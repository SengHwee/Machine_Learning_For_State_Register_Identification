module altor32_lite(clk_i, rst_i, intr_i, nmi_i, enable_i, \mem_dat_i[0] , \mem_dat_i[1] , \mem_dat_i[2] , \mem_dat_i[3] , \mem_dat_i[4] , \mem_dat_i[5] , \mem_dat_i[6] , \mem_dat_i[7] , \mem_dat_i[8] , \mem_dat_i[9] , \mem_dat_i[10] , \mem_dat_i[11] , \mem_dat_i[12] , \mem_dat_i[13] , \mem_dat_i[14] , \mem_dat_i[15] , \mem_dat_i[16] , \mem_dat_i[17] , \mem_dat_i[18] , \mem_dat_i[19] , \mem_dat_i[20] , \mem_dat_i[21] , \mem_dat_i[22] , \mem_dat_i[23] , \mem_dat_i[24] , \mem_dat_i[25] , \mem_dat_i[26] , \mem_dat_i[27] , \mem_dat_i[28] , \mem_dat_i[29] , \mem_dat_i[30] , \mem_dat_i[31] , mem_stall_i, mem_ack_i, fault_o, break_o, \mem_addr_o[0] , \mem_addr_o[1] , \mem_addr_o[2] , \mem_addr_o[3] , \mem_addr_o[4] , \mem_addr_o[5] , \mem_addr_o[6] , \mem_addr_o[7] , \mem_addr_o[8] , \mem_addr_o[9] , \mem_addr_o[10] , \mem_addr_o[11] , \mem_addr_o[12] , \mem_addr_o[13] , \mem_addr_o[14] , \mem_addr_o[15] , \mem_addr_o[16] , \mem_addr_o[17] , \mem_addr_o[18] , \mem_addr_o[19] , \mem_addr_o[20] , \mem_addr_o[21] , \mem_addr_o[22] , \mem_addr_o[23] , \mem_addr_o[24] , \mem_addr_o[25] , \mem_addr_o[26] , \mem_addr_o[27] , \mem_addr_o[28] , \mem_addr_o[29] , \mem_addr_o[30] , \mem_addr_o[31] , \mem_dat_o[0] , \mem_dat_o[1] , \mem_dat_o[2] , \mem_dat_o[3] , \mem_dat_o[4] , \mem_dat_o[5] , \mem_dat_o[6] , \mem_dat_o[7] , \mem_dat_o[8] , \mem_dat_o[9] , \mem_dat_o[10] , \mem_dat_o[11] , \mem_dat_o[12] , \mem_dat_o[13] , \mem_dat_o[14] , \mem_dat_o[15] , \mem_dat_o[16] , \mem_dat_o[17] , \mem_dat_o[18] , \mem_dat_o[19] , \mem_dat_o[20] , \mem_dat_o[21] , \mem_dat_o[22] , \mem_dat_o[23] , \mem_dat_o[24] , \mem_dat_o[25] , \mem_dat_o[26] , \mem_dat_o[27] , \mem_dat_o[28] , \mem_dat_o[29] , \mem_dat_o[30] , \mem_dat_o[31] , \mem_cti_o[0] , \mem_cti_o[1] , \mem_cti_o[2] , mem_cyc_o, mem_stb_o, mem_we_o, \mem_sel_o[0] , \mem_sel_o[1] , \mem_sel_o[2] , \mem_sel_o[3] );

wire REGFILE_SIM_reg_bank__0reg_r10_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r10_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r11_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r12_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r13_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r14_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r15_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r16_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r17_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r18_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r19_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r20_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r21_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r22_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r23_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r24_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r25_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r26_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r27_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r28_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r29_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r30_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r31_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r3_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r4_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r5_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r6_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r7_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r8_31_0__9_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__0_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__10_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__11_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__12_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__13_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__14_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__15_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__16_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__17_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__18_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__19_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__1_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__20_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__21_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__22_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__23_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__24_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__25_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__26_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__27_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__28_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__29_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__2_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__30_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__31_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__3_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__4_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__5_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__6_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__7_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__8_; 
wire REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__9_; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2099_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2111_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2115_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2120_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2121_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2124_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2132_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2136_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2144_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2147_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2150_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2156_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2162_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2174_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2180_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2182_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2186_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2192_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2204_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2206_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2210_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2216_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2222_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2234_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2246_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2249_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2252_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2255_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2261_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2264_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2267_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2270_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2273_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2276_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2279_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2282_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2285_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2288_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2291_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2294_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2297_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2300_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2303_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2306_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2309_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2312_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2315_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2318_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2321_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2324_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2327_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2330_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2333_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2336_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2344_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2347_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2350_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2353_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2356_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2359_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2362_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2365_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2368_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2371_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2374_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2377_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2380_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2383_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2386_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2389_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2392_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2395_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2398_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2401_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2404_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2407_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2410_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2413_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2416_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2419_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2422_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2425_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2428_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2431_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2434_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2436_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2439_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2445_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2448_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2451_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2454_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2457_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2460_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2463_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2466_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2469_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2475_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2478_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2481_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2487_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2490_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2493_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2499_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2502_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2505_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2511_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2514_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2521_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2523_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2527_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2535_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2539_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2551_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2557_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2559_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2563_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2566_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2569_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2571_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2574_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2575_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2577_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2578_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2581_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2582_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2583_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2586_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2587_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2589_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2590_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2593_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2595_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2598_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2599_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2601_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2602_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2605_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2608_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2611_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2614_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2620_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2623_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2626_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2629_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2632_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2633_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2635_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2638_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2641_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2644_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2647_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2650_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2653_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2656_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2657_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2659_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2662_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2665_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2666_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2668_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2671_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2674_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2677_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2678_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2680_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2683_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2686_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2689_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2690_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2692_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2695_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2698_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2701_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2702_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2704_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2706_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2710_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2713_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2714_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2718_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2722_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2725_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2726_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2728_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2730_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2734_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2737_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2738_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2740_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2742_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2746_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2749_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2750_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2752_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2754_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2758_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2761_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2762_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2764_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2765_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2766_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2770_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2773_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2774_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2776_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2778_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2782_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2785_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2786_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2788_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2789_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2790_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2794_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2797_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2798_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2800_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2801_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2804_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2806_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2809_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2810_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2812_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2813_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2816_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2817_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2820_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2822_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2825_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2826_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2828_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2831_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2832_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2834_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2835_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2838_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2840_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2843_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2844_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2846_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2847_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2850_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2852_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2855_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2856_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2858_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2859_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2862_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2864_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2867_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2868_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2870_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2871_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2874_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2876_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2879_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2880_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2882_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2883_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2886_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2887_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2888_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2892_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2895_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2896_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2898_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2899_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2902_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2904_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2907_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2908_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2910_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2911_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2914_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2920_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2923_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2926_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2932_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2935_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2938_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2944_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2947_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2948_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2950_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2956_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2959_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2961_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2969_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2972_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2973_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2981_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2985_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2991_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2993_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2997_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n2999_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3003_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3005_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3009_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3011_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3015_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3017_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3021_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3023_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3027_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3029_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3033_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3035_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3039_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3041_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3047_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3051_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3058_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3059_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3060_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3061_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3064_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3067_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3070_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3071_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3073_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3076_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3079_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3082_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3083_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3085_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3088_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3091_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3094_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3095_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3097_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3103_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3115_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3118_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3121_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3124_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3128_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3133_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3136_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3148_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3168_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3180_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3183_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3188_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3192_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3204_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3208_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3213_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3216_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3228_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3243_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3249_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3252_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3253_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3255_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3261_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3264_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3267_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3273_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3276_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3277_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3279_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3285_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3291_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3294_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3297_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3303_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3306_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3309_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3315_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3318_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3321_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3327_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3330_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3333_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3347_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3350_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3353_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3359_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3362_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3365_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3371_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3374_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3375_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3377_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3383_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3386_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3389_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3395_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3398_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3399_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3401_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3407_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3410_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3413_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3419_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3422_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3425_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3426_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3428_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3431_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3434_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3447_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3450_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3459_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3520_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3523_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3532_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3535_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3559_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3564_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3568_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3571_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3574_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3576_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3577_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3580_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3582_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3583_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3586_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3588_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3589_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3592_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3595_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3598_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3601_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3604_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3607_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3610_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3613_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3616_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3619_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3622_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3625_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3628_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3631_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3633_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3634_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3637_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3640_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3643_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3646_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3649_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3652_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3655_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3657_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3658_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3661_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3664_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3666_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3667_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3670_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3673_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3676_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3678_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3679_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3682_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3685_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3688_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3690_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3691_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3694_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3697_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3702_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3703_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3706_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3711_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3714_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3715_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3718_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3723_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3726_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3727_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3730_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3735_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3738_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3739_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3742_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3747_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3750_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3751_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3754_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3759_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3762_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3763_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3765_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3766_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3771_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3774_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3775_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3778_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3783_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3786_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3787_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3789_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3790_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3795_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3798_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3799_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3801_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3804_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3807_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3810_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3811_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3813_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3815_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3816_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3819_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3822_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3825_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3827_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3828_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3831_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3833_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3834_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3837_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3840_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3843_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3845_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3846_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3849_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3852_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3855_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3857_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3858_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3861_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3864_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3867_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3869_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3870_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3873_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3876_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3879_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3881_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3882_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3885_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3887_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3888_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3893_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3896_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3897_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3899_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3902_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3905_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3908_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3909_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3911_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3914_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3920_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3923_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3926_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3932_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3935_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3938_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3944_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3947_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3948_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3950_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3956_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3959_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3962_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3968_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3971_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3972_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3974_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3980_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3983_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3986_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3991_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3992_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3995_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3998_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n3999_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4003_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4004_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4007_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4010_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4011_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4015_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4016_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4019_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4022_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4023_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4027_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4028_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4031_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4034_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4035_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4039_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4040_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4043_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4047_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4051_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4059_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4060_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4063_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4066_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4069_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4071_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4072_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4075_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4078_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4081_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4083_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4084_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4087_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4090_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4093_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4095_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4096_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4099_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4108_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4111_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4120_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4123_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4128_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4132_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4138_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4148_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4178_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4182_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4188_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4206_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4208_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4218_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4238_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4253_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4274_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4277_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4286_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4292_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4304_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4316_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4328_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4340_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4352_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4364_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4372_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4375_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4384_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4396_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4399_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4408_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4426_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4436_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4445_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4448_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4450_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4454_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4457_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4460_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4466_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4469_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4472_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4478_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4481_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4484_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4490_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4493_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4496_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4502_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4505_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4508_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4514_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4520_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4521_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4524_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4532_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4536_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4548_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4557_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4560_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4564_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4566_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4569_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4572_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4575_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4576_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4578_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4581_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4582_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4584_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4587_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4588_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4590_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4593_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4596_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4599_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4602_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4605_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4608_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4611_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4614_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4620_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4623_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4626_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4629_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4632_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4633_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4635_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4638_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4641_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4644_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4647_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4650_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4653_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4656_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4657_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4659_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4664_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4665_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4667_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4668_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4671_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4673_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4676_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4677_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4679_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4680_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4683_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4685_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4688_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4689_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4691_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4692_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4695_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4697_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4701_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4703_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4704_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4707_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4711_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4713_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4715_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4719_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4723_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4725_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4727_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4728_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4731_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4735_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4737_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4739_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4740_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4743_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4747_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4749_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4751_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4752_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4755_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4759_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4761_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4763_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4764_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4765_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4767_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4771_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4773_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4775_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4776_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4779_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4783_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4785_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4787_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4788_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4789_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4791_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4794_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4797_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4799_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4800_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4803_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4806_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4809_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4811_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4812_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4815_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4817_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4820_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4823_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4826_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4827_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4829_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4832_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4833_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4835_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4838_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4841_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4844_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4845_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4847_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4850_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4853_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4856_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4857_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4859_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4862_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4865_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4868_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4869_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4871_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4874_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4877_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4880_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4881_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4883_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4886_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4887_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4889_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4892_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4895_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4897_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4898_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4901_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4904_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4907_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4909_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4910_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4913_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4921_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4925_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4933_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4937_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4945_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4948_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4949_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4957_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4961_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4969_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4972_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4973_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4981_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4985_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4989_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4992_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4993_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4997_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n4998_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5001_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5004_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5005_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5009_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5010_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5013_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5016_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5017_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5021_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5022_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5025_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5028_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5029_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5033_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5034_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5037_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5040_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5041_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5046_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5049_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5052_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5058_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5060_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5061_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5064_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5066_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5069_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5070_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5072_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5073_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5076_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5078_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5081_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5082_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5084_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5085_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5088_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5090_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5093_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5094_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5096_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5097_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5108_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5118_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5121_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5123_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5133_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5138_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5147_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5150_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5153_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5162_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5174_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5178_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5182_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5183_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5186_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5198_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5206_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5210_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5213_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5218_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5222_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5234_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5238_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5243_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5246_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5253_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5274_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5277_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5286_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5292_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5304_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5316_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5328_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5340_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5344_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5352_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5364_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5372_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5375_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5384_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5396_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5399_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5408_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5426_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5436_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5439_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5447_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5450_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5459_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5521_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5524_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5527_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5536_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5539_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5548_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5551_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5557_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5559_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5560_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5563_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5564_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5566_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5568_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5569_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5571_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5572_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5574_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5575_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5576_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5577_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5578_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5580_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5581_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5582_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5583_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5584_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5586_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5587_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5588_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5589_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5590_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5592_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5593_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5595_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5596_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5598_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5599_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5601_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5602_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5604_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5605_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5607_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5608_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5610_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5611_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5613_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5614_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5616_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5619_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5620_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5622_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5623_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5625_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5626_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5628_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5629_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5631_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5632_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5633_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5634_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5635_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5637_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5638_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5640_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5641_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5643_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5644_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5646_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5647_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5649_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5650_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5652_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5653_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5655_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5656_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5658_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5659_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5661_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5662_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5664_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5665_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5666_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5667_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5668_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5670_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5671_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5673_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5674_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5676_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5677_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5678_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5679_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5680_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5682_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5683_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5685_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5686_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5688_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5689_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5690_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5691_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5692_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5694_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5695_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5697_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5698_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5701_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5702_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5703_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5704_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5706_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5707_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5710_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5711_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5713_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5714_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5715_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5719_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5722_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5723_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5725_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5726_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5727_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5728_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5730_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5731_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5734_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5735_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5737_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5738_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5739_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5740_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5742_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5743_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5746_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5747_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5749_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5750_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5751_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5752_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5754_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5755_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5758_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5759_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5761_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5762_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5763_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5764_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5765_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5766_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5767_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5770_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5771_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5773_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5774_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5775_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5776_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5778_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5782_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5783_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5785_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5786_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5787_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5788_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5789_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5790_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5791_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5794_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5795_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5797_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5798_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5799_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5800_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5801_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5803_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5804_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5806_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5807_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5809_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5810_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5811_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5812_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5813_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5815_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5816_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5817_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5819_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5820_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5822_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5823_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5825_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5826_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5827_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5828_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5829_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5831_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5832_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5833_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5834_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5835_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5837_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5838_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5841_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5843_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5844_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5845_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5846_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5847_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5849_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5850_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5852_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5853_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5855_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5856_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5857_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5858_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5859_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5861_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5862_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5864_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5865_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5867_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5868_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5869_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5870_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5871_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5873_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5874_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5876_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5877_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5879_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5880_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5881_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5882_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5883_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5885_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5886_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5887_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5888_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5889_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5892_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5893_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5895_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5896_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5897_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5898_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5899_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5902_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5904_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5905_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5907_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5908_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5909_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5910_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5911_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5913_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5914_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5917_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5920_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5921_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5923_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5925_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5926_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5929_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5932_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5933_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5935_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5937_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5938_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5941_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5944_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5945_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5947_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5948_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5949_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5950_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5953_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5956_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5957_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5959_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5961_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5965_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5968_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5969_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5971_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5972_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5973_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5974_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5977_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5980_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5981_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5983_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5985_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5986_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5989_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5991_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5992_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5993_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5995_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5997_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5998_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n5999_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6001_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6003_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6004_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6005_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6007_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6009_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6010_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6011_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6013_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6015_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6016_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6017_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6019_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6021_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6022_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6025_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6027_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6028_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6029_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6031_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6033_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6034_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6035_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6037_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6039_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6040_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6041_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6043_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6046_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6047_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6049_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6051_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6052_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6055_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6058_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6059_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6060_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6061_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6063_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6064_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6066_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6067_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6069_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6070_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6071_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6072_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6073_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6075_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6076_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6078_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6079_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6081_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6082_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6083_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6085_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6087_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6088_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6090_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6091_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6093_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6094_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6095_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6096_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6097_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6099_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6103_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6108_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6111_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6115_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6118_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6120_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6121_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6123_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6124_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6128_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6132_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6133_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6136_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6138_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6144_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6147_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6148_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6150_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6153_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6156_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6162_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6168_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6174_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6178_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6180_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6182_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6183_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6186_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6188_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6192_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6198_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6204_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6208_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6210_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6213_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6216_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6218_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6222_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6228_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6234_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6238_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6243_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6246_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6249_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6252_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6253_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6255_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6258_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6261_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6264_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6270_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6273_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6274_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6276_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6277_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6279_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6282_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6285_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6286_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6288_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6291_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6292_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6294_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6297_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6300_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6303_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6304_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6306_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6309_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6312_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6315_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6316_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6318_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6321_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6324_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6327_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6330_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6333_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6336_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6340_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6344_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6347_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6350_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6352_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6353_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6356_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6359_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6362_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6364_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6365_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6368_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6371_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6372_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6374_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6375_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6377_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6380_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6383_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6384_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6386_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6392_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6395_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6396_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6398_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6399_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6401_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6404_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6407_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6408_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6410_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6413_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6416_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6419_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6422_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6425_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6426_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6428_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6431_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6434_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6436_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6439_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6445_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6447_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6448_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6451_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6454_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6457_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6459_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6460_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6463_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6466_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6469_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6472_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6475_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6478_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6481_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6484_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6487_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6490_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6493_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6496_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6499_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6502_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6505_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6508_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6514_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6520_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6521_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6523_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6524_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6527_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6532_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6535_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6536_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6539_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6548_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6551_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6557_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6559_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6560_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6563_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6564_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6566_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6568_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6569_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6571_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6574_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6575_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6576_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6577_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6578_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6580_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6581_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6582_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6583_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6584_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6586_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6587_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6588_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6589_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6590_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6592_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6593_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6595_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6596_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6598_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6599_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6601_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6602_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6604_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6605_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6607_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6608_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6610_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6611_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6613_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6614_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6616_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6619_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6620_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6622_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6623_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6625_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6626_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6628_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6629_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6631_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6632_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6634_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6635_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6637_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6638_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6640_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6641_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6643_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6644_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6646_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6647_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6649_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6650_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6652_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6653_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6655_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6656_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6657_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6658_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6659_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6661_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6662_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6664_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6665_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6666_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6667_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6668_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6670_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6671_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6673_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6674_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6676_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6677_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6678_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6679_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6680_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6682_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6683_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6685_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6686_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6688_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6689_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6690_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6691_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6692_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6695_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6697_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6698_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6701_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6702_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6703_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6704_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6706_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6707_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6710_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6711_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6713_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6714_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6715_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6718_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6719_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6722_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6723_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6725_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6726_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6727_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6728_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6730_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6731_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6734_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6735_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6737_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6738_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6739_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6740_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6742_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6743_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6746_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6747_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6749_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6750_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6751_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6752_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6754_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6758_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6759_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6761_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6762_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6763_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6764_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6765_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6766_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6767_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6770_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6771_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6773_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6774_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6775_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6776_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6778_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6779_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6782_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6783_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6785_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6786_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6787_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6788_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6789_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6790_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6791_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6794_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6795_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6797_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6798_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6799_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6800_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6801_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6803_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6804_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6806_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6807_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6809_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6810_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6811_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6812_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6813_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6815_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6817_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6819_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6820_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6822_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6823_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6825_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6826_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6827_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6828_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6829_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6831_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6832_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6833_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6834_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6835_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6837_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6838_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6840_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6841_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6843_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6844_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6845_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6846_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6847_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6849_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6850_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6852_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6853_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6855_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6856_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6857_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6858_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6859_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6861_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6862_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6864_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6865_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6867_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6868_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6869_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6870_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6871_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6873_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6874_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6876_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6879_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6880_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6881_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6882_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6883_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6885_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6886_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6887_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6888_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6889_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6892_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6893_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6895_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6896_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6897_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6898_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6899_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6901_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6902_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6904_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6905_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6907_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6908_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6909_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6910_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6911_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6913_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6914_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6917_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6920_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6921_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6923_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6925_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6926_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6929_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6932_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6933_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6935_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6937_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6941_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6944_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6945_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6947_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6948_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6949_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6950_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6953_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6956_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6957_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6959_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6961_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6962_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6965_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6968_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6969_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6971_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6972_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6973_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6974_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6977_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6980_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6981_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6983_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6985_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6986_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6989_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6991_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6992_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6993_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6995_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6997_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n6998_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7001_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7003_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7004_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7005_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7007_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7009_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7010_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7011_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7013_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7015_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7016_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7017_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7019_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7021_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7022_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7023_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7025_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7027_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7028_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7029_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7031_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7033_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7034_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7035_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7037_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7039_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7040_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7041_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7043_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7046_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7047_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7049_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7051_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7052_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7055_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7058_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7059_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7061_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7063_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7064_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7066_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7067_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7069_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7070_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7071_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7072_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7073_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7075_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7076_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7078_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7079_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7081_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7082_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7083_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7084_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7085_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7087_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7088_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7090_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7091_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7093_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7094_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7095_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7096_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7097_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7099_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7103_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7108_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7111_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7115_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7118_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7120_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7123_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7124_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7128_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7132_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7133_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7136_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7138_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7144_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7147_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7148_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7150_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7153_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7156_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7162_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7168_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7174_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7178_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7180_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7183_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7186_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7188_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7192_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7198_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7204_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7206_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7208_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7210_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7213_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7216_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7218_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7222_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7228_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7234_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7238_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7246_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7249_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7252_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7253_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7255_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7258_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7261_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7264_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7267_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7270_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7273_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7274_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7276_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7277_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7279_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7282_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7285_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7286_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7288_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7291_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7292_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7294_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7297_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7300_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7303_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7306_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7309_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7312_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7315_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7316_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7318_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7321_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7324_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7327_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7328_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7330_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7333_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7336_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7340_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7344_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7347_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7350_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7352_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7353_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7356_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7359_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7362_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7364_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7368_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7371_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7372_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7374_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7375_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7377_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7380_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7383_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7384_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7386_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7389_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7392_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7395_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7396_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7398_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7399_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7401_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7404_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7407_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7408_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7410_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7413_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7416_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7419_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7422_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7425_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7428_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7431_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7434_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7436_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7439_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7445_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7447_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7448_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7450_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7451_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7454_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7457_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7459_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7460_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7463_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7466_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7469_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7472_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7475_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7478_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7481_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7484_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7490_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7493_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7496_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7499_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7502_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7505_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7508_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7511_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7514_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7520_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7521_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7523_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7524_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7527_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7532_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7535_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7536_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7539_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7551_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7557_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7559_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7560_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7563_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7564_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7566_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7568_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7569_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7571_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7572_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7574_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7575_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7576_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7577_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7578_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7580_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7581_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7582_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7583_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7584_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7586_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7587_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7588_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7589_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7590_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7592_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7593_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7595_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7596_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7598_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7599_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7601_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7602_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7604_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7605_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7607_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7608_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7610_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7611_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7613_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7614_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7616_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7619_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7620_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7622_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7623_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7625_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7626_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7628_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7629_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7631_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7632_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7633_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7634_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7635_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7637_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7638_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7640_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7641_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7643_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7644_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7646_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7647_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7649_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7650_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7652_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7653_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7655_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7656_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7657_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7658_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7659_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7661_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7662_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7664_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7665_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7666_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7668_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7670_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7671_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7673_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7674_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7676_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7677_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7678_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7679_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7680_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7682_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7683_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7685_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7686_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7688_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7689_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7690_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7691_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7692_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7694_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7695_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7697_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7698_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7701_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7702_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7703_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7704_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7706_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7707_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7710_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7711_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7713_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7714_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7715_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7718_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7719_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7722_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7723_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7725_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7726_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7727_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7730_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7731_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7734_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7735_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7737_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7738_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7739_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7740_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7742_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7743_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7746_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7747_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7749_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7750_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7751_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7752_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7754_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7755_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7758_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7759_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7761_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7762_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7763_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7764_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7765_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7766_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7767_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7770_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7771_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7773_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7774_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7775_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7776_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7778_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7779_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7782_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7783_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7785_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7786_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7787_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7788_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7790_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7791_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7794_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7795_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7797_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7798_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7799_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7800_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7801_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7803_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7804_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7806_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7807_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7809_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7810_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7811_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7812_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7813_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7815_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7816_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7817_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7819_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7820_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7822_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7823_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7825_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7826_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7827_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7828_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7829_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7831_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7832_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7833_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7834_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7835_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7837_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7838_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7840_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7841_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7843_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7844_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7845_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7846_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7847_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7849_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7852_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7853_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7855_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7856_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7857_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7858_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7859_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7861_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7862_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7864_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7865_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7867_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7868_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7869_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7870_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7871_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7873_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7874_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7876_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7877_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7879_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7880_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7881_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7882_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7883_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7885_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7886_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7887_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7888_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7889_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7892_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7893_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7895_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7896_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7897_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7898_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7899_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7901_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7902_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7904_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7905_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7907_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7908_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7909_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7910_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7913_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7914_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7917_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7920_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7921_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7923_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7925_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7926_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7929_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7932_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7933_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7935_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7937_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7938_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7941_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7944_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7945_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7947_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7948_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7949_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7950_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7953_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7956_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7957_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7959_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7961_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7962_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7965_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7968_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7969_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7971_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7973_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7974_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7977_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7980_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7981_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7983_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7985_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7986_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7989_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7991_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7992_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7993_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7995_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7997_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7998_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n7999_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8001_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8003_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8004_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8005_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8007_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8009_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8010_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8011_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8013_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8015_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8016_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8017_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8019_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8021_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8022_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8023_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8025_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8027_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8028_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8029_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8031_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8034_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8035_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8037_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8039_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8040_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8041_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8043_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8046_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8047_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8049_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8051_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8052_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8055_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8058_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8059_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8060_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8061_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8063_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8064_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8066_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8067_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8069_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8070_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8071_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8072_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8073_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8075_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8076_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8078_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8079_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8081_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8082_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8083_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8084_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8085_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8087_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8088_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8090_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8091_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8093_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8095_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8096_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8097_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8099_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8103_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8108_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8111_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8115_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8118_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8120_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8121_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8123_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8124_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8128_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8131_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8132_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8133_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8136_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8138_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8144_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8147_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8148_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8150_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8153_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8156_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8162_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8168_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8174_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8178_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8180_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8182_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8183_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8186_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8188_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8192_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8198_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8204_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8206_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8208_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8210_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8213_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8218_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8222_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8228_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8234_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8238_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8243_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8246_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8249_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8252_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8253_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8255_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8258_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8261_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8264_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8267_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8270_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8273_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8274_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8276_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8279_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8282_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8285_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8286_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8288_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8291_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8292_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8294_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8297_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8300_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8303_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8304_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8306_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8309_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8312_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8314_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8315_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8316_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8318_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8321_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8324_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8327_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8328_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8330_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8333_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8336_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8340_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8344_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8347_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8350_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8352_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8353_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8356_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8359_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8362_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8364_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8365_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8368_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8371_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8372_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8374_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8375_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8377_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8380_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8383_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8384_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8386_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8389_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8392_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8395_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8396_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8398_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8401_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8404_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8407_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8408_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8410_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8413_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8416_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8419_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8422_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8425_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8426_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8428_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8431_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8434_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8436_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8439_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8445_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8447_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8448_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8450_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8451_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8454_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8457_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8459_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8463_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8466_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8469_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8472_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8475_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8478_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8481_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8484_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8487_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8490_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8493_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8496_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8497_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8499_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8502_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8505_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8508_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8511_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8514_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8520_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8523_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8524_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8527_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8532_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8535_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8536_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8539_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8548_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8551_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8557_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8558_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8559_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8560_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8561_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8562_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8563_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8564_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8565_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8566_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8567_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8568_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8569_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8570_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8571_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8572_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8573_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8574_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8575_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8576_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8577_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8578_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8579_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8580_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8581_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8583_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8584_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8585_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8586_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8587_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8588_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8589_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8590_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8591_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8592_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8593_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8594_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8595_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8596_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8597_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8598_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8599_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8600_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8601_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8602_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8603_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8604_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8605_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8606_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8607_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8608_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8609_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8610_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8611_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8612_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8613_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8614_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8615_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8616_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8617_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8618_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8619_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8620_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8621_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8622_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8623_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8624_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8625_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8626_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8627_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8628_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8629_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8630_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8631_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8632_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8633_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8634_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8635_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8636_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8637_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8638_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8639_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8640_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8641_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8642_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8644_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8645_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8646_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8647_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8648_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8649_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8650_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8651_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8652_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8653_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8654_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8655_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8656_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8657_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8658_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8659_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8660_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8661_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8662_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8663_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8664_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8665_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8666_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8667_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8668_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8669_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8670_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8671_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8672_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8673_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8674_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8675_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8676_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8677_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8678_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8679_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8680_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8681_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8682_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8683_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8684_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8685_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8686_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8687_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8688_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8689_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8690_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8691_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8692_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8693_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8694_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8695_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8696_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8697_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8698_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8699_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8700_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8701_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8702_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8703_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8705_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8706_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8707_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8708_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8709_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8710_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8711_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8712_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8713_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8714_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8715_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8716_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8717_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8718_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8719_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8720_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8721_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8722_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8723_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8724_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8725_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8726_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8727_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8728_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8729_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8730_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8731_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8732_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8733_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8734_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8735_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8736_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8737_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8738_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8739_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8740_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8741_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8742_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8743_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8744_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8745_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8746_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8747_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8748_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8749_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8750_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8751_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8752_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8753_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8754_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8755_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8756_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8757_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8758_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8759_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8760_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8761_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8762_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8763_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8764_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8766_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8767_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8768_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8769_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8770_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8771_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8772_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8773_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8774_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8775_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8776_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8777_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8778_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8779_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8780_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8781_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8782_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8783_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8784_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8785_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8786_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8787_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8788_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8789_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8790_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8791_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8792_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8793_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8794_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8795_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8796_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8797_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8798_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8799_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8800_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8801_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8802_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8803_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8804_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8805_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8806_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8807_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8808_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8809_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8810_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8811_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8812_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8813_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8814_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8815_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8816_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8817_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8818_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8819_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8820_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8821_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8822_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8823_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8824_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8825_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8827_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8828_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8829_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8830_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8831_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8832_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8833_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8834_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8835_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8836_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8837_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8838_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8839_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8840_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8841_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8842_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8843_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8844_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8845_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8846_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8847_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8848_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8849_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8850_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8851_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8852_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8853_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8854_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8855_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8856_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8857_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8858_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8859_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8860_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8861_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8862_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8863_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8864_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8865_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8866_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8867_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8868_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8869_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8870_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8871_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8872_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8873_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8874_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8875_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8876_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8877_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8878_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8879_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8880_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8881_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8882_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8883_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8884_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8885_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8886_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8888_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8889_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8890_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8891_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8892_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8893_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8894_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8895_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8896_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8897_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8898_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8899_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8900_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8901_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8902_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8903_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8904_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8905_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8906_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8907_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8908_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8909_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8910_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8911_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8912_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8913_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8914_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8915_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8916_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8917_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8918_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8919_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8920_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8921_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8922_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8923_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8924_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8925_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8926_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8927_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8928_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8929_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8930_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8931_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8932_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8933_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8934_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8935_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8936_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8937_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8938_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8939_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8940_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8941_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8942_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8943_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8944_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8945_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8946_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8947_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8949_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8950_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8951_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8952_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8953_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8954_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8955_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8956_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8957_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8958_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8959_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8960_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8961_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8962_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8963_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8964_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8965_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8966_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8967_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8968_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8969_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8970_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8971_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8972_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8973_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8974_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8975_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8976_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8977_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8978_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8979_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8980_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8981_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8982_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8983_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8984_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8985_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8986_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8987_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8988_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8989_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8990_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8991_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8992_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8993_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8994_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8995_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8996_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8997_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8998_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n8999_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9000_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9001_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9002_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9003_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9004_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9005_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9006_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9007_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9008_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9010_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9011_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9012_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9013_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9014_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9015_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9016_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9017_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9018_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9019_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9020_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9021_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9022_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9023_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9024_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9025_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9026_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9027_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9028_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9029_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9030_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9031_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9032_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9033_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9034_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9035_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9036_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9037_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9038_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9039_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9040_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9041_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9042_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9043_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9044_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9045_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9046_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9047_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9048_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9049_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9050_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9051_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9052_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9053_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9054_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9055_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9056_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9057_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9058_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9059_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9060_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9061_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9062_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9063_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9064_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9065_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9066_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9067_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9068_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9069_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9071_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9072_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9073_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9074_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9075_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9076_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9077_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9078_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9079_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9080_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9081_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9082_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9083_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9084_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9085_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9086_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9087_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9088_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9089_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9090_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9091_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9092_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9093_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9094_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9095_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9096_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9097_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9098_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9099_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9100_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9101_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9102_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9103_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9104_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9105_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9106_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9107_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9108_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9109_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9110_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9111_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9112_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9113_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9114_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9115_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9116_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9117_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9118_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9119_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9120_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9121_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9122_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9123_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9124_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9125_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9126_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9127_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9128_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9129_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9130_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9132_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9133_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9134_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9135_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9136_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9137_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9138_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9139_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9140_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9141_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9142_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9143_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9144_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9145_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9146_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9147_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9148_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9149_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9150_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9151_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9152_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9153_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9154_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9155_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9156_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9157_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9158_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9159_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9160_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9161_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9162_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9163_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9164_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9165_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9166_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9167_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9168_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9169_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9170_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9171_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9172_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9173_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9174_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9175_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9176_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9177_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9178_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9179_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9180_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9181_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9182_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9183_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9184_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9185_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9186_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9187_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9188_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9189_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9190_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9191_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9193_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9194_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9195_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9196_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9197_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9198_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9199_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9200_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9201_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9202_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9203_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9204_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9205_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9206_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9207_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9208_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9209_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9210_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9211_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9212_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9213_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9214_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9215_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9216_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9217_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9218_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9219_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9220_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9221_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9222_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9223_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9224_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9225_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9226_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9227_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9228_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9229_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9230_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9231_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9232_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9233_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9234_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9235_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9236_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9237_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9238_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9239_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9240_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9241_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9242_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9243_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9244_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9245_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9246_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9247_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9248_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9249_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9250_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9251_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9252_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9254_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9255_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9256_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9257_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9258_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9259_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9260_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9261_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9262_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9263_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9264_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9265_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9266_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9267_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9268_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9269_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9270_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9271_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9272_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9273_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9274_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9275_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9276_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9277_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9278_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9279_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9280_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9281_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9282_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9283_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9284_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9285_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9286_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9287_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9288_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9289_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9290_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9291_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9292_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9293_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9294_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9295_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9296_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9297_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9298_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9299_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9300_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9301_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9302_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9303_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9304_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9305_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9306_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9307_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9308_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9309_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9310_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9311_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9312_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9313_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9315_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9316_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9317_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9318_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9319_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9320_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9321_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9322_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9323_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9324_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9325_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9326_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9327_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9328_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9329_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9330_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9331_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9332_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9333_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9334_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9335_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9336_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9337_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9338_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9339_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9340_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9341_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9342_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9343_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9344_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9345_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9346_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9347_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9348_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9349_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9350_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9351_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9352_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9353_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9354_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9355_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9356_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9357_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9358_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9359_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9360_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9361_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9362_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9363_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9364_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9365_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9366_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9367_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9368_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9369_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9370_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9371_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9372_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9373_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9374_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9376_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9377_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9378_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9379_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9380_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9381_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9382_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9383_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9384_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9385_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9386_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9387_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9388_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9389_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9390_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9391_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9392_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9393_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9394_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9395_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9396_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9397_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9398_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9399_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9400_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9401_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9402_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9403_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9404_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9405_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9406_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9407_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9408_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9409_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9410_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9411_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9412_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9413_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9414_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9415_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9416_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9417_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9418_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9419_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9420_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9421_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9422_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9423_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9424_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9425_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9426_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9427_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9428_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9429_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9430_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9431_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9432_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9433_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9434_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9435_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9437_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9438_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9439_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9440_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9441_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9442_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9443_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9444_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9445_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9446_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9447_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9448_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9449_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9450_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9451_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9452_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9453_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9454_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9455_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9456_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9457_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9458_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9459_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9460_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9461_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9462_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9463_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9464_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9465_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9466_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9467_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9468_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9469_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9470_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9471_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9472_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9473_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9474_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9475_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9476_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9477_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9478_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9479_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9480_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9481_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9482_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9483_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9484_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9485_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9486_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9487_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9488_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9489_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9490_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9491_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9492_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9493_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9494_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9495_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9496_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9498_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9499_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9500_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9501_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9502_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9503_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9504_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9505_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9506_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9507_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9508_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9509_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9510_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9511_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9512_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9513_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9514_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9515_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9516_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9517_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9518_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9519_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9520_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9521_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9522_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9523_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9524_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9525_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9526_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9527_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9528_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9529_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9530_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9531_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9532_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9533_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9534_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9535_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9536_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9537_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9538_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9539_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9540_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9541_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9542_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9543_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9544_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9545_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9546_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9547_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9548_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9549_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9550_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9551_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9552_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9553_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9554_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9555_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9556_; 
wire REGFILE_SIM_reg_bank__abc_34819_new_n9557_; 
wire REGFILE_SIM_reg_bank_ra_i_0_; 
wire REGFILE_SIM_reg_bank_ra_i_1_; 
wire REGFILE_SIM_reg_bank_ra_i_2_; 
wire REGFILE_SIM_reg_bank_ra_i_3_; 
wire REGFILE_SIM_reg_bank_ra_i_4_; 
wire REGFILE_SIM_reg_bank_ra_i_4_bF_buf0_; 
wire REGFILE_SIM_reg_bank_ra_i_4_bF_buf1_; 
wire REGFILE_SIM_reg_bank_ra_i_4_bF_buf2_; 
wire REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_; 
wire REGFILE_SIM_reg_bank_rb_i_0_; 
wire REGFILE_SIM_reg_bank_rb_i_1_; 
wire REGFILE_SIM_reg_bank_rb_i_2_; 
wire REGFILE_SIM_reg_bank_rb_i_3_; 
wire REGFILE_SIM_reg_bank_rb_i_4_; 
wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf0_; 
wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf1_; 
wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf2_; 
wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf3_; 
wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf4_; 
wire REGFILE_SIM_reg_bank_rb_i_4_bF_buf5_; 
wire REGFILE_SIM_reg_bank_rd_i_0_; 
wire REGFILE_SIM_reg_bank_rd_i_1_; 
wire REGFILE_SIM_reg_bank_rd_i_2_; 
wire REGFILE_SIM_reg_bank_rd_i_3_; 
wire REGFILE_SIM_reg_bank_rd_i_4_; 
wire REGFILE_SIM_reg_bank_reg_r10_0_; 
wire REGFILE_SIM_reg_bank_reg_r10_10_; 
wire REGFILE_SIM_reg_bank_reg_r10_11_; 
wire REGFILE_SIM_reg_bank_reg_r10_12_; 
wire REGFILE_SIM_reg_bank_reg_r10_13_; 
wire REGFILE_SIM_reg_bank_reg_r10_14_; 
wire REGFILE_SIM_reg_bank_reg_r10_15_; 
wire REGFILE_SIM_reg_bank_reg_r10_16_; 
wire REGFILE_SIM_reg_bank_reg_r10_17_; 
wire REGFILE_SIM_reg_bank_reg_r10_18_; 
wire REGFILE_SIM_reg_bank_reg_r10_19_; 
wire REGFILE_SIM_reg_bank_reg_r10_1_; 
wire REGFILE_SIM_reg_bank_reg_r10_20_; 
wire REGFILE_SIM_reg_bank_reg_r10_21_; 
wire REGFILE_SIM_reg_bank_reg_r10_22_; 
wire REGFILE_SIM_reg_bank_reg_r10_23_; 
wire REGFILE_SIM_reg_bank_reg_r10_24_; 
wire REGFILE_SIM_reg_bank_reg_r10_25_; 
wire REGFILE_SIM_reg_bank_reg_r10_26_; 
wire REGFILE_SIM_reg_bank_reg_r10_27_; 
wire REGFILE_SIM_reg_bank_reg_r10_28_; 
wire REGFILE_SIM_reg_bank_reg_r10_29_; 
wire REGFILE_SIM_reg_bank_reg_r10_2_; 
wire REGFILE_SIM_reg_bank_reg_r10_30_; 
wire REGFILE_SIM_reg_bank_reg_r10_31_; 
wire REGFILE_SIM_reg_bank_reg_r10_3_; 
wire REGFILE_SIM_reg_bank_reg_r10_4_; 
wire REGFILE_SIM_reg_bank_reg_r10_5_; 
wire REGFILE_SIM_reg_bank_reg_r10_6_; 
wire REGFILE_SIM_reg_bank_reg_r10_7_; 
wire REGFILE_SIM_reg_bank_reg_r10_8_; 
wire REGFILE_SIM_reg_bank_reg_r10_9_; 
wire REGFILE_SIM_reg_bank_reg_r11_0_; 
wire REGFILE_SIM_reg_bank_reg_r11_10_; 
wire REGFILE_SIM_reg_bank_reg_r11_11_; 
wire REGFILE_SIM_reg_bank_reg_r11_12_; 
wire REGFILE_SIM_reg_bank_reg_r11_13_; 
wire REGFILE_SIM_reg_bank_reg_r11_14_; 
wire REGFILE_SIM_reg_bank_reg_r11_15_; 
wire REGFILE_SIM_reg_bank_reg_r11_16_; 
wire REGFILE_SIM_reg_bank_reg_r11_17_; 
wire REGFILE_SIM_reg_bank_reg_r11_18_; 
wire REGFILE_SIM_reg_bank_reg_r11_19_; 
wire REGFILE_SIM_reg_bank_reg_r11_1_; 
wire REGFILE_SIM_reg_bank_reg_r11_20_; 
wire REGFILE_SIM_reg_bank_reg_r11_21_; 
wire REGFILE_SIM_reg_bank_reg_r11_22_; 
wire REGFILE_SIM_reg_bank_reg_r11_23_; 
wire REGFILE_SIM_reg_bank_reg_r11_24_; 
wire REGFILE_SIM_reg_bank_reg_r11_25_; 
wire REGFILE_SIM_reg_bank_reg_r11_26_; 
wire REGFILE_SIM_reg_bank_reg_r11_27_; 
wire REGFILE_SIM_reg_bank_reg_r11_28_; 
wire REGFILE_SIM_reg_bank_reg_r11_29_; 
wire REGFILE_SIM_reg_bank_reg_r11_2_; 
wire REGFILE_SIM_reg_bank_reg_r11_30_; 
wire REGFILE_SIM_reg_bank_reg_r11_31_; 
wire REGFILE_SIM_reg_bank_reg_r11_3_; 
wire REGFILE_SIM_reg_bank_reg_r11_4_; 
wire REGFILE_SIM_reg_bank_reg_r11_5_; 
wire REGFILE_SIM_reg_bank_reg_r11_6_; 
wire REGFILE_SIM_reg_bank_reg_r11_7_; 
wire REGFILE_SIM_reg_bank_reg_r11_8_; 
wire REGFILE_SIM_reg_bank_reg_r11_9_; 
wire REGFILE_SIM_reg_bank_reg_r12_0_; 
wire REGFILE_SIM_reg_bank_reg_r12_10_; 
wire REGFILE_SIM_reg_bank_reg_r12_11_; 
wire REGFILE_SIM_reg_bank_reg_r12_12_; 
wire REGFILE_SIM_reg_bank_reg_r12_13_; 
wire REGFILE_SIM_reg_bank_reg_r12_14_; 
wire REGFILE_SIM_reg_bank_reg_r12_15_; 
wire REGFILE_SIM_reg_bank_reg_r12_16_; 
wire REGFILE_SIM_reg_bank_reg_r12_17_; 
wire REGFILE_SIM_reg_bank_reg_r12_18_; 
wire REGFILE_SIM_reg_bank_reg_r12_19_; 
wire REGFILE_SIM_reg_bank_reg_r12_1_; 
wire REGFILE_SIM_reg_bank_reg_r12_20_; 
wire REGFILE_SIM_reg_bank_reg_r12_21_; 
wire REGFILE_SIM_reg_bank_reg_r12_22_; 
wire REGFILE_SIM_reg_bank_reg_r12_23_; 
wire REGFILE_SIM_reg_bank_reg_r12_24_; 
wire REGFILE_SIM_reg_bank_reg_r12_25_; 
wire REGFILE_SIM_reg_bank_reg_r12_26_; 
wire REGFILE_SIM_reg_bank_reg_r12_27_; 
wire REGFILE_SIM_reg_bank_reg_r12_28_; 
wire REGFILE_SIM_reg_bank_reg_r12_29_; 
wire REGFILE_SIM_reg_bank_reg_r12_2_; 
wire REGFILE_SIM_reg_bank_reg_r12_30_; 
wire REGFILE_SIM_reg_bank_reg_r12_31_; 
wire REGFILE_SIM_reg_bank_reg_r12_3_; 
wire REGFILE_SIM_reg_bank_reg_r12_4_; 
wire REGFILE_SIM_reg_bank_reg_r12_5_; 
wire REGFILE_SIM_reg_bank_reg_r12_6_; 
wire REGFILE_SIM_reg_bank_reg_r12_7_; 
wire REGFILE_SIM_reg_bank_reg_r12_8_; 
wire REGFILE_SIM_reg_bank_reg_r12_9_; 
wire REGFILE_SIM_reg_bank_reg_r13_0_; 
wire REGFILE_SIM_reg_bank_reg_r13_10_; 
wire REGFILE_SIM_reg_bank_reg_r13_11_; 
wire REGFILE_SIM_reg_bank_reg_r13_12_; 
wire REGFILE_SIM_reg_bank_reg_r13_13_; 
wire REGFILE_SIM_reg_bank_reg_r13_14_; 
wire REGFILE_SIM_reg_bank_reg_r13_15_; 
wire REGFILE_SIM_reg_bank_reg_r13_16_; 
wire REGFILE_SIM_reg_bank_reg_r13_17_; 
wire REGFILE_SIM_reg_bank_reg_r13_18_; 
wire REGFILE_SIM_reg_bank_reg_r13_19_; 
wire REGFILE_SIM_reg_bank_reg_r13_1_; 
wire REGFILE_SIM_reg_bank_reg_r13_20_; 
wire REGFILE_SIM_reg_bank_reg_r13_21_; 
wire REGFILE_SIM_reg_bank_reg_r13_22_; 
wire REGFILE_SIM_reg_bank_reg_r13_23_; 
wire REGFILE_SIM_reg_bank_reg_r13_24_; 
wire REGFILE_SIM_reg_bank_reg_r13_25_; 
wire REGFILE_SIM_reg_bank_reg_r13_26_; 
wire REGFILE_SIM_reg_bank_reg_r13_27_; 
wire REGFILE_SIM_reg_bank_reg_r13_28_; 
wire REGFILE_SIM_reg_bank_reg_r13_29_; 
wire REGFILE_SIM_reg_bank_reg_r13_2_; 
wire REGFILE_SIM_reg_bank_reg_r13_30_; 
wire REGFILE_SIM_reg_bank_reg_r13_31_; 
wire REGFILE_SIM_reg_bank_reg_r13_3_; 
wire REGFILE_SIM_reg_bank_reg_r13_4_; 
wire REGFILE_SIM_reg_bank_reg_r13_5_; 
wire REGFILE_SIM_reg_bank_reg_r13_6_; 
wire REGFILE_SIM_reg_bank_reg_r13_7_; 
wire REGFILE_SIM_reg_bank_reg_r13_8_; 
wire REGFILE_SIM_reg_bank_reg_r13_9_; 
wire REGFILE_SIM_reg_bank_reg_r14_0_; 
wire REGFILE_SIM_reg_bank_reg_r14_10_; 
wire REGFILE_SIM_reg_bank_reg_r14_11_; 
wire REGFILE_SIM_reg_bank_reg_r14_12_; 
wire REGFILE_SIM_reg_bank_reg_r14_13_; 
wire REGFILE_SIM_reg_bank_reg_r14_14_; 
wire REGFILE_SIM_reg_bank_reg_r14_15_; 
wire REGFILE_SIM_reg_bank_reg_r14_16_; 
wire REGFILE_SIM_reg_bank_reg_r14_17_; 
wire REGFILE_SIM_reg_bank_reg_r14_18_; 
wire REGFILE_SIM_reg_bank_reg_r14_19_; 
wire REGFILE_SIM_reg_bank_reg_r14_1_; 
wire REGFILE_SIM_reg_bank_reg_r14_20_; 
wire REGFILE_SIM_reg_bank_reg_r14_21_; 
wire REGFILE_SIM_reg_bank_reg_r14_22_; 
wire REGFILE_SIM_reg_bank_reg_r14_23_; 
wire REGFILE_SIM_reg_bank_reg_r14_24_; 
wire REGFILE_SIM_reg_bank_reg_r14_25_; 
wire REGFILE_SIM_reg_bank_reg_r14_26_; 
wire REGFILE_SIM_reg_bank_reg_r14_27_; 
wire REGFILE_SIM_reg_bank_reg_r14_28_; 
wire REGFILE_SIM_reg_bank_reg_r14_29_; 
wire REGFILE_SIM_reg_bank_reg_r14_2_; 
wire REGFILE_SIM_reg_bank_reg_r14_30_; 
wire REGFILE_SIM_reg_bank_reg_r14_31_; 
wire REGFILE_SIM_reg_bank_reg_r14_3_; 
wire REGFILE_SIM_reg_bank_reg_r14_4_; 
wire REGFILE_SIM_reg_bank_reg_r14_5_; 
wire REGFILE_SIM_reg_bank_reg_r14_6_; 
wire REGFILE_SIM_reg_bank_reg_r14_7_; 
wire REGFILE_SIM_reg_bank_reg_r14_8_; 
wire REGFILE_SIM_reg_bank_reg_r14_9_; 
wire REGFILE_SIM_reg_bank_reg_r15_0_; 
wire REGFILE_SIM_reg_bank_reg_r15_10_; 
wire REGFILE_SIM_reg_bank_reg_r15_11_; 
wire REGFILE_SIM_reg_bank_reg_r15_12_; 
wire REGFILE_SIM_reg_bank_reg_r15_13_; 
wire REGFILE_SIM_reg_bank_reg_r15_14_; 
wire REGFILE_SIM_reg_bank_reg_r15_15_; 
wire REGFILE_SIM_reg_bank_reg_r15_16_; 
wire REGFILE_SIM_reg_bank_reg_r15_17_; 
wire REGFILE_SIM_reg_bank_reg_r15_18_; 
wire REGFILE_SIM_reg_bank_reg_r15_19_; 
wire REGFILE_SIM_reg_bank_reg_r15_1_; 
wire REGFILE_SIM_reg_bank_reg_r15_20_; 
wire REGFILE_SIM_reg_bank_reg_r15_21_; 
wire REGFILE_SIM_reg_bank_reg_r15_22_; 
wire REGFILE_SIM_reg_bank_reg_r15_23_; 
wire REGFILE_SIM_reg_bank_reg_r15_24_; 
wire REGFILE_SIM_reg_bank_reg_r15_25_; 
wire REGFILE_SIM_reg_bank_reg_r15_26_; 
wire REGFILE_SIM_reg_bank_reg_r15_27_; 
wire REGFILE_SIM_reg_bank_reg_r15_28_; 
wire REGFILE_SIM_reg_bank_reg_r15_29_; 
wire REGFILE_SIM_reg_bank_reg_r15_2_; 
wire REGFILE_SIM_reg_bank_reg_r15_30_; 
wire REGFILE_SIM_reg_bank_reg_r15_31_; 
wire REGFILE_SIM_reg_bank_reg_r15_3_; 
wire REGFILE_SIM_reg_bank_reg_r15_4_; 
wire REGFILE_SIM_reg_bank_reg_r15_5_; 
wire REGFILE_SIM_reg_bank_reg_r15_6_; 
wire REGFILE_SIM_reg_bank_reg_r15_7_; 
wire REGFILE_SIM_reg_bank_reg_r15_8_; 
wire REGFILE_SIM_reg_bank_reg_r15_9_; 
wire REGFILE_SIM_reg_bank_reg_r16_0_; 
wire REGFILE_SIM_reg_bank_reg_r16_10_; 
wire REGFILE_SIM_reg_bank_reg_r16_11_; 
wire REGFILE_SIM_reg_bank_reg_r16_12_; 
wire REGFILE_SIM_reg_bank_reg_r16_13_; 
wire REGFILE_SIM_reg_bank_reg_r16_14_; 
wire REGFILE_SIM_reg_bank_reg_r16_15_; 
wire REGFILE_SIM_reg_bank_reg_r16_16_; 
wire REGFILE_SIM_reg_bank_reg_r16_17_; 
wire REGFILE_SIM_reg_bank_reg_r16_18_; 
wire REGFILE_SIM_reg_bank_reg_r16_19_; 
wire REGFILE_SIM_reg_bank_reg_r16_1_; 
wire REGFILE_SIM_reg_bank_reg_r16_20_; 
wire REGFILE_SIM_reg_bank_reg_r16_21_; 
wire REGFILE_SIM_reg_bank_reg_r16_22_; 
wire REGFILE_SIM_reg_bank_reg_r16_23_; 
wire REGFILE_SIM_reg_bank_reg_r16_24_; 
wire REGFILE_SIM_reg_bank_reg_r16_25_; 
wire REGFILE_SIM_reg_bank_reg_r16_26_; 
wire REGFILE_SIM_reg_bank_reg_r16_27_; 
wire REGFILE_SIM_reg_bank_reg_r16_28_; 
wire REGFILE_SIM_reg_bank_reg_r16_29_; 
wire REGFILE_SIM_reg_bank_reg_r16_2_; 
wire REGFILE_SIM_reg_bank_reg_r16_30_; 
wire REGFILE_SIM_reg_bank_reg_r16_31_; 
wire REGFILE_SIM_reg_bank_reg_r16_3_; 
wire REGFILE_SIM_reg_bank_reg_r16_4_; 
wire REGFILE_SIM_reg_bank_reg_r16_5_; 
wire REGFILE_SIM_reg_bank_reg_r16_6_; 
wire REGFILE_SIM_reg_bank_reg_r16_7_; 
wire REGFILE_SIM_reg_bank_reg_r16_8_; 
wire REGFILE_SIM_reg_bank_reg_r16_9_; 
wire REGFILE_SIM_reg_bank_reg_r17_0_; 
wire REGFILE_SIM_reg_bank_reg_r17_10_; 
wire REGFILE_SIM_reg_bank_reg_r17_11_; 
wire REGFILE_SIM_reg_bank_reg_r17_12_; 
wire REGFILE_SIM_reg_bank_reg_r17_13_; 
wire REGFILE_SIM_reg_bank_reg_r17_14_; 
wire REGFILE_SIM_reg_bank_reg_r17_15_; 
wire REGFILE_SIM_reg_bank_reg_r17_16_; 
wire REGFILE_SIM_reg_bank_reg_r17_17_; 
wire REGFILE_SIM_reg_bank_reg_r17_18_; 
wire REGFILE_SIM_reg_bank_reg_r17_19_; 
wire REGFILE_SIM_reg_bank_reg_r17_1_; 
wire REGFILE_SIM_reg_bank_reg_r17_20_; 
wire REGFILE_SIM_reg_bank_reg_r17_21_; 
wire REGFILE_SIM_reg_bank_reg_r17_22_; 
wire REGFILE_SIM_reg_bank_reg_r17_23_; 
wire REGFILE_SIM_reg_bank_reg_r17_24_; 
wire REGFILE_SIM_reg_bank_reg_r17_25_; 
wire REGFILE_SIM_reg_bank_reg_r17_26_; 
wire REGFILE_SIM_reg_bank_reg_r17_27_; 
wire REGFILE_SIM_reg_bank_reg_r17_28_; 
wire REGFILE_SIM_reg_bank_reg_r17_29_; 
wire REGFILE_SIM_reg_bank_reg_r17_2_; 
wire REGFILE_SIM_reg_bank_reg_r17_30_; 
wire REGFILE_SIM_reg_bank_reg_r17_31_; 
wire REGFILE_SIM_reg_bank_reg_r17_3_; 
wire REGFILE_SIM_reg_bank_reg_r17_4_; 
wire REGFILE_SIM_reg_bank_reg_r17_5_; 
wire REGFILE_SIM_reg_bank_reg_r17_6_; 
wire REGFILE_SIM_reg_bank_reg_r17_7_; 
wire REGFILE_SIM_reg_bank_reg_r17_8_; 
wire REGFILE_SIM_reg_bank_reg_r17_9_; 
wire REGFILE_SIM_reg_bank_reg_r18_0_; 
wire REGFILE_SIM_reg_bank_reg_r18_10_; 
wire REGFILE_SIM_reg_bank_reg_r18_11_; 
wire REGFILE_SIM_reg_bank_reg_r18_12_; 
wire REGFILE_SIM_reg_bank_reg_r18_13_; 
wire REGFILE_SIM_reg_bank_reg_r18_14_; 
wire REGFILE_SIM_reg_bank_reg_r18_15_; 
wire REGFILE_SIM_reg_bank_reg_r18_16_; 
wire REGFILE_SIM_reg_bank_reg_r18_17_; 
wire REGFILE_SIM_reg_bank_reg_r18_18_; 
wire REGFILE_SIM_reg_bank_reg_r18_19_; 
wire REGFILE_SIM_reg_bank_reg_r18_1_; 
wire REGFILE_SIM_reg_bank_reg_r18_20_; 
wire REGFILE_SIM_reg_bank_reg_r18_21_; 
wire REGFILE_SIM_reg_bank_reg_r18_22_; 
wire REGFILE_SIM_reg_bank_reg_r18_23_; 
wire REGFILE_SIM_reg_bank_reg_r18_24_; 
wire REGFILE_SIM_reg_bank_reg_r18_25_; 
wire REGFILE_SIM_reg_bank_reg_r18_26_; 
wire REGFILE_SIM_reg_bank_reg_r18_27_; 
wire REGFILE_SIM_reg_bank_reg_r18_28_; 
wire REGFILE_SIM_reg_bank_reg_r18_29_; 
wire REGFILE_SIM_reg_bank_reg_r18_2_; 
wire REGFILE_SIM_reg_bank_reg_r18_30_; 
wire REGFILE_SIM_reg_bank_reg_r18_31_; 
wire REGFILE_SIM_reg_bank_reg_r18_3_; 
wire REGFILE_SIM_reg_bank_reg_r18_4_; 
wire REGFILE_SIM_reg_bank_reg_r18_5_; 
wire REGFILE_SIM_reg_bank_reg_r18_6_; 
wire REGFILE_SIM_reg_bank_reg_r18_7_; 
wire REGFILE_SIM_reg_bank_reg_r18_8_; 
wire REGFILE_SIM_reg_bank_reg_r18_9_; 
wire REGFILE_SIM_reg_bank_reg_r19_0_; 
wire REGFILE_SIM_reg_bank_reg_r19_10_; 
wire REGFILE_SIM_reg_bank_reg_r19_11_; 
wire REGFILE_SIM_reg_bank_reg_r19_12_; 
wire REGFILE_SIM_reg_bank_reg_r19_13_; 
wire REGFILE_SIM_reg_bank_reg_r19_14_; 
wire REGFILE_SIM_reg_bank_reg_r19_15_; 
wire REGFILE_SIM_reg_bank_reg_r19_16_; 
wire REGFILE_SIM_reg_bank_reg_r19_17_; 
wire REGFILE_SIM_reg_bank_reg_r19_18_; 
wire REGFILE_SIM_reg_bank_reg_r19_19_; 
wire REGFILE_SIM_reg_bank_reg_r19_1_; 
wire REGFILE_SIM_reg_bank_reg_r19_20_; 
wire REGFILE_SIM_reg_bank_reg_r19_21_; 
wire REGFILE_SIM_reg_bank_reg_r19_22_; 
wire REGFILE_SIM_reg_bank_reg_r19_23_; 
wire REGFILE_SIM_reg_bank_reg_r19_24_; 
wire REGFILE_SIM_reg_bank_reg_r19_25_; 
wire REGFILE_SIM_reg_bank_reg_r19_26_; 
wire REGFILE_SIM_reg_bank_reg_r19_27_; 
wire REGFILE_SIM_reg_bank_reg_r19_28_; 
wire REGFILE_SIM_reg_bank_reg_r19_29_; 
wire REGFILE_SIM_reg_bank_reg_r19_2_; 
wire REGFILE_SIM_reg_bank_reg_r19_30_; 
wire REGFILE_SIM_reg_bank_reg_r19_31_; 
wire REGFILE_SIM_reg_bank_reg_r19_3_; 
wire REGFILE_SIM_reg_bank_reg_r19_4_; 
wire REGFILE_SIM_reg_bank_reg_r19_5_; 
wire REGFILE_SIM_reg_bank_reg_r19_6_; 
wire REGFILE_SIM_reg_bank_reg_r19_7_; 
wire REGFILE_SIM_reg_bank_reg_r19_8_; 
wire REGFILE_SIM_reg_bank_reg_r19_9_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_0_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_10_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_11_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_12_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_13_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_14_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_15_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_16_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_17_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_18_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_19_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_1_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_20_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_21_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_22_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_23_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_24_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_25_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_26_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_27_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_28_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_29_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_2_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_30_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_31_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_3_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_4_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_5_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_6_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_7_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_8_; 
wire REGFILE_SIM_reg_bank_reg_r1_sp_9_; 
wire REGFILE_SIM_reg_bank_reg_r20_0_; 
wire REGFILE_SIM_reg_bank_reg_r20_10_; 
wire REGFILE_SIM_reg_bank_reg_r20_11_; 
wire REGFILE_SIM_reg_bank_reg_r20_12_; 
wire REGFILE_SIM_reg_bank_reg_r20_13_; 
wire REGFILE_SIM_reg_bank_reg_r20_14_; 
wire REGFILE_SIM_reg_bank_reg_r20_15_; 
wire REGFILE_SIM_reg_bank_reg_r20_16_; 
wire REGFILE_SIM_reg_bank_reg_r20_17_; 
wire REGFILE_SIM_reg_bank_reg_r20_18_; 
wire REGFILE_SIM_reg_bank_reg_r20_19_; 
wire REGFILE_SIM_reg_bank_reg_r20_1_; 
wire REGFILE_SIM_reg_bank_reg_r20_20_; 
wire REGFILE_SIM_reg_bank_reg_r20_21_; 
wire REGFILE_SIM_reg_bank_reg_r20_22_; 
wire REGFILE_SIM_reg_bank_reg_r20_23_; 
wire REGFILE_SIM_reg_bank_reg_r20_24_; 
wire REGFILE_SIM_reg_bank_reg_r20_25_; 
wire REGFILE_SIM_reg_bank_reg_r20_26_; 
wire REGFILE_SIM_reg_bank_reg_r20_27_; 
wire REGFILE_SIM_reg_bank_reg_r20_28_; 
wire REGFILE_SIM_reg_bank_reg_r20_29_; 
wire REGFILE_SIM_reg_bank_reg_r20_2_; 
wire REGFILE_SIM_reg_bank_reg_r20_30_; 
wire REGFILE_SIM_reg_bank_reg_r20_31_; 
wire REGFILE_SIM_reg_bank_reg_r20_3_; 
wire REGFILE_SIM_reg_bank_reg_r20_4_; 
wire REGFILE_SIM_reg_bank_reg_r20_5_; 
wire REGFILE_SIM_reg_bank_reg_r20_6_; 
wire REGFILE_SIM_reg_bank_reg_r20_7_; 
wire REGFILE_SIM_reg_bank_reg_r20_8_; 
wire REGFILE_SIM_reg_bank_reg_r20_9_; 
wire REGFILE_SIM_reg_bank_reg_r21_0_; 
wire REGFILE_SIM_reg_bank_reg_r21_10_; 
wire REGFILE_SIM_reg_bank_reg_r21_11_; 
wire REGFILE_SIM_reg_bank_reg_r21_12_; 
wire REGFILE_SIM_reg_bank_reg_r21_13_; 
wire REGFILE_SIM_reg_bank_reg_r21_14_; 
wire REGFILE_SIM_reg_bank_reg_r21_15_; 
wire REGFILE_SIM_reg_bank_reg_r21_16_; 
wire REGFILE_SIM_reg_bank_reg_r21_17_; 
wire REGFILE_SIM_reg_bank_reg_r21_18_; 
wire REGFILE_SIM_reg_bank_reg_r21_19_; 
wire REGFILE_SIM_reg_bank_reg_r21_1_; 
wire REGFILE_SIM_reg_bank_reg_r21_20_; 
wire REGFILE_SIM_reg_bank_reg_r21_21_; 
wire REGFILE_SIM_reg_bank_reg_r21_22_; 
wire REGFILE_SIM_reg_bank_reg_r21_23_; 
wire REGFILE_SIM_reg_bank_reg_r21_24_; 
wire REGFILE_SIM_reg_bank_reg_r21_25_; 
wire REGFILE_SIM_reg_bank_reg_r21_26_; 
wire REGFILE_SIM_reg_bank_reg_r21_27_; 
wire REGFILE_SIM_reg_bank_reg_r21_28_; 
wire REGFILE_SIM_reg_bank_reg_r21_29_; 
wire REGFILE_SIM_reg_bank_reg_r21_2_; 
wire REGFILE_SIM_reg_bank_reg_r21_30_; 
wire REGFILE_SIM_reg_bank_reg_r21_31_; 
wire REGFILE_SIM_reg_bank_reg_r21_3_; 
wire REGFILE_SIM_reg_bank_reg_r21_4_; 
wire REGFILE_SIM_reg_bank_reg_r21_5_; 
wire REGFILE_SIM_reg_bank_reg_r21_6_; 
wire REGFILE_SIM_reg_bank_reg_r21_7_; 
wire REGFILE_SIM_reg_bank_reg_r21_8_; 
wire REGFILE_SIM_reg_bank_reg_r21_9_; 
wire REGFILE_SIM_reg_bank_reg_r22_0_; 
wire REGFILE_SIM_reg_bank_reg_r22_10_; 
wire REGFILE_SIM_reg_bank_reg_r22_11_; 
wire REGFILE_SIM_reg_bank_reg_r22_12_; 
wire REGFILE_SIM_reg_bank_reg_r22_13_; 
wire REGFILE_SIM_reg_bank_reg_r22_14_; 
wire REGFILE_SIM_reg_bank_reg_r22_15_; 
wire REGFILE_SIM_reg_bank_reg_r22_16_; 
wire REGFILE_SIM_reg_bank_reg_r22_17_; 
wire REGFILE_SIM_reg_bank_reg_r22_18_; 
wire REGFILE_SIM_reg_bank_reg_r22_19_; 
wire REGFILE_SIM_reg_bank_reg_r22_1_; 
wire REGFILE_SIM_reg_bank_reg_r22_20_; 
wire REGFILE_SIM_reg_bank_reg_r22_21_; 
wire REGFILE_SIM_reg_bank_reg_r22_22_; 
wire REGFILE_SIM_reg_bank_reg_r22_23_; 
wire REGFILE_SIM_reg_bank_reg_r22_24_; 
wire REGFILE_SIM_reg_bank_reg_r22_25_; 
wire REGFILE_SIM_reg_bank_reg_r22_26_; 
wire REGFILE_SIM_reg_bank_reg_r22_27_; 
wire REGFILE_SIM_reg_bank_reg_r22_28_; 
wire REGFILE_SIM_reg_bank_reg_r22_29_; 
wire REGFILE_SIM_reg_bank_reg_r22_2_; 
wire REGFILE_SIM_reg_bank_reg_r22_30_; 
wire REGFILE_SIM_reg_bank_reg_r22_31_; 
wire REGFILE_SIM_reg_bank_reg_r22_3_; 
wire REGFILE_SIM_reg_bank_reg_r22_4_; 
wire REGFILE_SIM_reg_bank_reg_r22_5_; 
wire REGFILE_SIM_reg_bank_reg_r22_6_; 
wire REGFILE_SIM_reg_bank_reg_r22_7_; 
wire REGFILE_SIM_reg_bank_reg_r22_8_; 
wire REGFILE_SIM_reg_bank_reg_r22_9_; 
wire REGFILE_SIM_reg_bank_reg_r23_0_; 
wire REGFILE_SIM_reg_bank_reg_r23_10_; 
wire REGFILE_SIM_reg_bank_reg_r23_11_; 
wire REGFILE_SIM_reg_bank_reg_r23_12_; 
wire REGFILE_SIM_reg_bank_reg_r23_13_; 
wire REGFILE_SIM_reg_bank_reg_r23_14_; 
wire REGFILE_SIM_reg_bank_reg_r23_15_; 
wire REGFILE_SIM_reg_bank_reg_r23_16_; 
wire REGFILE_SIM_reg_bank_reg_r23_17_; 
wire REGFILE_SIM_reg_bank_reg_r23_18_; 
wire REGFILE_SIM_reg_bank_reg_r23_19_; 
wire REGFILE_SIM_reg_bank_reg_r23_1_; 
wire REGFILE_SIM_reg_bank_reg_r23_20_; 
wire REGFILE_SIM_reg_bank_reg_r23_21_; 
wire REGFILE_SIM_reg_bank_reg_r23_22_; 
wire REGFILE_SIM_reg_bank_reg_r23_23_; 
wire REGFILE_SIM_reg_bank_reg_r23_24_; 
wire REGFILE_SIM_reg_bank_reg_r23_25_; 
wire REGFILE_SIM_reg_bank_reg_r23_26_; 
wire REGFILE_SIM_reg_bank_reg_r23_27_; 
wire REGFILE_SIM_reg_bank_reg_r23_28_; 
wire REGFILE_SIM_reg_bank_reg_r23_29_; 
wire REGFILE_SIM_reg_bank_reg_r23_2_; 
wire REGFILE_SIM_reg_bank_reg_r23_30_; 
wire REGFILE_SIM_reg_bank_reg_r23_31_; 
wire REGFILE_SIM_reg_bank_reg_r23_3_; 
wire REGFILE_SIM_reg_bank_reg_r23_4_; 
wire REGFILE_SIM_reg_bank_reg_r23_5_; 
wire REGFILE_SIM_reg_bank_reg_r23_6_; 
wire REGFILE_SIM_reg_bank_reg_r23_7_; 
wire REGFILE_SIM_reg_bank_reg_r23_8_; 
wire REGFILE_SIM_reg_bank_reg_r23_9_; 
wire REGFILE_SIM_reg_bank_reg_r24_0_; 
wire REGFILE_SIM_reg_bank_reg_r24_10_; 
wire REGFILE_SIM_reg_bank_reg_r24_11_; 
wire REGFILE_SIM_reg_bank_reg_r24_12_; 
wire REGFILE_SIM_reg_bank_reg_r24_13_; 
wire REGFILE_SIM_reg_bank_reg_r24_14_; 
wire REGFILE_SIM_reg_bank_reg_r24_15_; 
wire REGFILE_SIM_reg_bank_reg_r24_16_; 
wire REGFILE_SIM_reg_bank_reg_r24_17_; 
wire REGFILE_SIM_reg_bank_reg_r24_18_; 
wire REGFILE_SIM_reg_bank_reg_r24_19_; 
wire REGFILE_SIM_reg_bank_reg_r24_1_; 
wire REGFILE_SIM_reg_bank_reg_r24_20_; 
wire REGFILE_SIM_reg_bank_reg_r24_21_; 
wire REGFILE_SIM_reg_bank_reg_r24_22_; 
wire REGFILE_SIM_reg_bank_reg_r24_23_; 
wire REGFILE_SIM_reg_bank_reg_r24_24_; 
wire REGFILE_SIM_reg_bank_reg_r24_25_; 
wire REGFILE_SIM_reg_bank_reg_r24_26_; 
wire REGFILE_SIM_reg_bank_reg_r24_27_; 
wire REGFILE_SIM_reg_bank_reg_r24_28_; 
wire REGFILE_SIM_reg_bank_reg_r24_29_; 
wire REGFILE_SIM_reg_bank_reg_r24_2_; 
wire REGFILE_SIM_reg_bank_reg_r24_30_; 
wire REGFILE_SIM_reg_bank_reg_r24_31_; 
wire REGFILE_SIM_reg_bank_reg_r24_3_; 
wire REGFILE_SIM_reg_bank_reg_r24_4_; 
wire REGFILE_SIM_reg_bank_reg_r24_5_; 
wire REGFILE_SIM_reg_bank_reg_r24_6_; 
wire REGFILE_SIM_reg_bank_reg_r24_7_; 
wire REGFILE_SIM_reg_bank_reg_r24_8_; 
wire REGFILE_SIM_reg_bank_reg_r24_9_; 
wire REGFILE_SIM_reg_bank_reg_r25_0_; 
wire REGFILE_SIM_reg_bank_reg_r25_10_; 
wire REGFILE_SIM_reg_bank_reg_r25_11_; 
wire REGFILE_SIM_reg_bank_reg_r25_12_; 
wire REGFILE_SIM_reg_bank_reg_r25_13_; 
wire REGFILE_SIM_reg_bank_reg_r25_14_; 
wire REGFILE_SIM_reg_bank_reg_r25_15_; 
wire REGFILE_SIM_reg_bank_reg_r25_16_; 
wire REGFILE_SIM_reg_bank_reg_r25_17_; 
wire REGFILE_SIM_reg_bank_reg_r25_18_; 
wire REGFILE_SIM_reg_bank_reg_r25_19_; 
wire REGFILE_SIM_reg_bank_reg_r25_1_; 
wire REGFILE_SIM_reg_bank_reg_r25_20_; 
wire REGFILE_SIM_reg_bank_reg_r25_21_; 
wire REGFILE_SIM_reg_bank_reg_r25_22_; 
wire REGFILE_SIM_reg_bank_reg_r25_23_; 
wire REGFILE_SIM_reg_bank_reg_r25_24_; 
wire REGFILE_SIM_reg_bank_reg_r25_25_; 
wire REGFILE_SIM_reg_bank_reg_r25_26_; 
wire REGFILE_SIM_reg_bank_reg_r25_27_; 
wire REGFILE_SIM_reg_bank_reg_r25_28_; 
wire REGFILE_SIM_reg_bank_reg_r25_29_; 
wire REGFILE_SIM_reg_bank_reg_r25_2_; 
wire REGFILE_SIM_reg_bank_reg_r25_30_; 
wire REGFILE_SIM_reg_bank_reg_r25_31_; 
wire REGFILE_SIM_reg_bank_reg_r25_3_; 
wire REGFILE_SIM_reg_bank_reg_r25_4_; 
wire REGFILE_SIM_reg_bank_reg_r25_5_; 
wire REGFILE_SIM_reg_bank_reg_r25_6_; 
wire REGFILE_SIM_reg_bank_reg_r25_7_; 
wire REGFILE_SIM_reg_bank_reg_r25_8_; 
wire REGFILE_SIM_reg_bank_reg_r25_9_; 
wire REGFILE_SIM_reg_bank_reg_r26_0_; 
wire REGFILE_SIM_reg_bank_reg_r26_10_; 
wire REGFILE_SIM_reg_bank_reg_r26_11_; 
wire REGFILE_SIM_reg_bank_reg_r26_12_; 
wire REGFILE_SIM_reg_bank_reg_r26_13_; 
wire REGFILE_SIM_reg_bank_reg_r26_14_; 
wire REGFILE_SIM_reg_bank_reg_r26_15_; 
wire REGFILE_SIM_reg_bank_reg_r26_16_; 
wire REGFILE_SIM_reg_bank_reg_r26_17_; 
wire REGFILE_SIM_reg_bank_reg_r26_18_; 
wire REGFILE_SIM_reg_bank_reg_r26_19_; 
wire REGFILE_SIM_reg_bank_reg_r26_1_; 
wire REGFILE_SIM_reg_bank_reg_r26_20_; 
wire REGFILE_SIM_reg_bank_reg_r26_21_; 
wire REGFILE_SIM_reg_bank_reg_r26_22_; 
wire REGFILE_SIM_reg_bank_reg_r26_23_; 
wire REGFILE_SIM_reg_bank_reg_r26_24_; 
wire REGFILE_SIM_reg_bank_reg_r26_25_; 
wire REGFILE_SIM_reg_bank_reg_r26_26_; 
wire REGFILE_SIM_reg_bank_reg_r26_27_; 
wire REGFILE_SIM_reg_bank_reg_r26_28_; 
wire REGFILE_SIM_reg_bank_reg_r26_29_; 
wire REGFILE_SIM_reg_bank_reg_r26_2_; 
wire REGFILE_SIM_reg_bank_reg_r26_30_; 
wire REGFILE_SIM_reg_bank_reg_r26_31_; 
wire REGFILE_SIM_reg_bank_reg_r26_3_; 
wire REGFILE_SIM_reg_bank_reg_r26_4_; 
wire REGFILE_SIM_reg_bank_reg_r26_5_; 
wire REGFILE_SIM_reg_bank_reg_r26_6_; 
wire REGFILE_SIM_reg_bank_reg_r26_7_; 
wire REGFILE_SIM_reg_bank_reg_r26_8_; 
wire REGFILE_SIM_reg_bank_reg_r26_9_; 
wire REGFILE_SIM_reg_bank_reg_r27_0_; 
wire REGFILE_SIM_reg_bank_reg_r27_10_; 
wire REGFILE_SIM_reg_bank_reg_r27_11_; 
wire REGFILE_SIM_reg_bank_reg_r27_12_; 
wire REGFILE_SIM_reg_bank_reg_r27_13_; 
wire REGFILE_SIM_reg_bank_reg_r27_14_; 
wire REGFILE_SIM_reg_bank_reg_r27_15_; 
wire REGFILE_SIM_reg_bank_reg_r27_16_; 
wire REGFILE_SIM_reg_bank_reg_r27_17_; 
wire REGFILE_SIM_reg_bank_reg_r27_18_; 
wire REGFILE_SIM_reg_bank_reg_r27_19_; 
wire REGFILE_SIM_reg_bank_reg_r27_1_; 
wire REGFILE_SIM_reg_bank_reg_r27_20_; 
wire REGFILE_SIM_reg_bank_reg_r27_21_; 
wire REGFILE_SIM_reg_bank_reg_r27_22_; 
wire REGFILE_SIM_reg_bank_reg_r27_23_; 
wire REGFILE_SIM_reg_bank_reg_r27_24_; 
wire REGFILE_SIM_reg_bank_reg_r27_25_; 
wire REGFILE_SIM_reg_bank_reg_r27_26_; 
wire REGFILE_SIM_reg_bank_reg_r27_27_; 
wire REGFILE_SIM_reg_bank_reg_r27_28_; 
wire REGFILE_SIM_reg_bank_reg_r27_29_; 
wire REGFILE_SIM_reg_bank_reg_r27_2_; 
wire REGFILE_SIM_reg_bank_reg_r27_30_; 
wire REGFILE_SIM_reg_bank_reg_r27_31_; 
wire REGFILE_SIM_reg_bank_reg_r27_3_; 
wire REGFILE_SIM_reg_bank_reg_r27_4_; 
wire REGFILE_SIM_reg_bank_reg_r27_5_; 
wire REGFILE_SIM_reg_bank_reg_r27_6_; 
wire REGFILE_SIM_reg_bank_reg_r27_7_; 
wire REGFILE_SIM_reg_bank_reg_r27_8_; 
wire REGFILE_SIM_reg_bank_reg_r27_9_; 
wire REGFILE_SIM_reg_bank_reg_r28_0_; 
wire REGFILE_SIM_reg_bank_reg_r28_10_; 
wire REGFILE_SIM_reg_bank_reg_r28_11_; 
wire REGFILE_SIM_reg_bank_reg_r28_12_; 
wire REGFILE_SIM_reg_bank_reg_r28_13_; 
wire REGFILE_SIM_reg_bank_reg_r28_14_; 
wire REGFILE_SIM_reg_bank_reg_r28_15_; 
wire REGFILE_SIM_reg_bank_reg_r28_16_; 
wire REGFILE_SIM_reg_bank_reg_r28_17_; 
wire REGFILE_SIM_reg_bank_reg_r28_18_; 
wire REGFILE_SIM_reg_bank_reg_r28_19_; 
wire REGFILE_SIM_reg_bank_reg_r28_1_; 
wire REGFILE_SIM_reg_bank_reg_r28_20_; 
wire REGFILE_SIM_reg_bank_reg_r28_21_; 
wire REGFILE_SIM_reg_bank_reg_r28_22_; 
wire REGFILE_SIM_reg_bank_reg_r28_23_; 
wire REGFILE_SIM_reg_bank_reg_r28_24_; 
wire REGFILE_SIM_reg_bank_reg_r28_25_; 
wire REGFILE_SIM_reg_bank_reg_r28_26_; 
wire REGFILE_SIM_reg_bank_reg_r28_27_; 
wire REGFILE_SIM_reg_bank_reg_r28_28_; 
wire REGFILE_SIM_reg_bank_reg_r28_29_; 
wire REGFILE_SIM_reg_bank_reg_r28_2_; 
wire REGFILE_SIM_reg_bank_reg_r28_30_; 
wire REGFILE_SIM_reg_bank_reg_r28_31_; 
wire REGFILE_SIM_reg_bank_reg_r28_3_; 
wire REGFILE_SIM_reg_bank_reg_r28_4_; 
wire REGFILE_SIM_reg_bank_reg_r28_5_; 
wire REGFILE_SIM_reg_bank_reg_r28_6_; 
wire REGFILE_SIM_reg_bank_reg_r28_7_; 
wire REGFILE_SIM_reg_bank_reg_r28_8_; 
wire REGFILE_SIM_reg_bank_reg_r28_9_; 
wire REGFILE_SIM_reg_bank_reg_r29_0_; 
wire REGFILE_SIM_reg_bank_reg_r29_10_; 
wire REGFILE_SIM_reg_bank_reg_r29_11_; 
wire REGFILE_SIM_reg_bank_reg_r29_12_; 
wire REGFILE_SIM_reg_bank_reg_r29_13_; 
wire REGFILE_SIM_reg_bank_reg_r29_14_; 
wire REGFILE_SIM_reg_bank_reg_r29_15_; 
wire REGFILE_SIM_reg_bank_reg_r29_16_; 
wire REGFILE_SIM_reg_bank_reg_r29_17_; 
wire REGFILE_SIM_reg_bank_reg_r29_18_; 
wire REGFILE_SIM_reg_bank_reg_r29_19_; 
wire REGFILE_SIM_reg_bank_reg_r29_1_; 
wire REGFILE_SIM_reg_bank_reg_r29_20_; 
wire REGFILE_SIM_reg_bank_reg_r29_21_; 
wire REGFILE_SIM_reg_bank_reg_r29_22_; 
wire REGFILE_SIM_reg_bank_reg_r29_23_; 
wire REGFILE_SIM_reg_bank_reg_r29_24_; 
wire REGFILE_SIM_reg_bank_reg_r29_25_; 
wire REGFILE_SIM_reg_bank_reg_r29_26_; 
wire REGFILE_SIM_reg_bank_reg_r29_27_; 
wire REGFILE_SIM_reg_bank_reg_r29_28_; 
wire REGFILE_SIM_reg_bank_reg_r29_29_; 
wire REGFILE_SIM_reg_bank_reg_r29_2_; 
wire REGFILE_SIM_reg_bank_reg_r29_30_; 
wire REGFILE_SIM_reg_bank_reg_r29_31_; 
wire REGFILE_SIM_reg_bank_reg_r29_3_; 
wire REGFILE_SIM_reg_bank_reg_r29_4_; 
wire REGFILE_SIM_reg_bank_reg_r29_5_; 
wire REGFILE_SIM_reg_bank_reg_r29_6_; 
wire REGFILE_SIM_reg_bank_reg_r29_7_; 
wire REGFILE_SIM_reg_bank_reg_r29_8_; 
wire REGFILE_SIM_reg_bank_reg_r29_9_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_0_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_10_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_11_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_12_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_13_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_14_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_15_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_16_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_17_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_18_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_19_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_1_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_20_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_21_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_22_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_23_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_24_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_25_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_26_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_27_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_28_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_29_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_2_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_30_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_31_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_3_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_4_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_5_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_6_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_7_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_8_; 
wire REGFILE_SIM_reg_bank_reg_r2_fp_9_; 
wire REGFILE_SIM_reg_bank_reg_r30_0_; 
wire REGFILE_SIM_reg_bank_reg_r30_10_; 
wire REGFILE_SIM_reg_bank_reg_r30_11_; 
wire REGFILE_SIM_reg_bank_reg_r30_12_; 
wire REGFILE_SIM_reg_bank_reg_r30_13_; 
wire REGFILE_SIM_reg_bank_reg_r30_14_; 
wire REGFILE_SIM_reg_bank_reg_r30_15_; 
wire REGFILE_SIM_reg_bank_reg_r30_16_; 
wire REGFILE_SIM_reg_bank_reg_r30_17_; 
wire REGFILE_SIM_reg_bank_reg_r30_18_; 
wire REGFILE_SIM_reg_bank_reg_r30_19_; 
wire REGFILE_SIM_reg_bank_reg_r30_1_; 
wire REGFILE_SIM_reg_bank_reg_r30_20_; 
wire REGFILE_SIM_reg_bank_reg_r30_21_; 
wire REGFILE_SIM_reg_bank_reg_r30_22_; 
wire REGFILE_SIM_reg_bank_reg_r30_23_; 
wire REGFILE_SIM_reg_bank_reg_r30_24_; 
wire REGFILE_SIM_reg_bank_reg_r30_25_; 
wire REGFILE_SIM_reg_bank_reg_r30_26_; 
wire REGFILE_SIM_reg_bank_reg_r30_27_; 
wire REGFILE_SIM_reg_bank_reg_r30_28_; 
wire REGFILE_SIM_reg_bank_reg_r30_29_; 
wire REGFILE_SIM_reg_bank_reg_r30_2_; 
wire REGFILE_SIM_reg_bank_reg_r30_30_; 
wire REGFILE_SIM_reg_bank_reg_r30_31_; 
wire REGFILE_SIM_reg_bank_reg_r30_3_; 
wire REGFILE_SIM_reg_bank_reg_r30_4_; 
wire REGFILE_SIM_reg_bank_reg_r30_5_; 
wire REGFILE_SIM_reg_bank_reg_r30_6_; 
wire REGFILE_SIM_reg_bank_reg_r30_7_; 
wire REGFILE_SIM_reg_bank_reg_r30_8_; 
wire REGFILE_SIM_reg_bank_reg_r30_9_; 
wire REGFILE_SIM_reg_bank_reg_r31_0_; 
wire REGFILE_SIM_reg_bank_reg_r31_10_; 
wire REGFILE_SIM_reg_bank_reg_r31_11_; 
wire REGFILE_SIM_reg_bank_reg_r31_12_; 
wire REGFILE_SIM_reg_bank_reg_r31_13_; 
wire REGFILE_SIM_reg_bank_reg_r31_14_; 
wire REGFILE_SIM_reg_bank_reg_r31_15_; 
wire REGFILE_SIM_reg_bank_reg_r31_16_; 
wire REGFILE_SIM_reg_bank_reg_r31_17_; 
wire REGFILE_SIM_reg_bank_reg_r31_18_; 
wire REGFILE_SIM_reg_bank_reg_r31_19_; 
wire REGFILE_SIM_reg_bank_reg_r31_1_; 
wire REGFILE_SIM_reg_bank_reg_r31_20_; 
wire REGFILE_SIM_reg_bank_reg_r31_21_; 
wire REGFILE_SIM_reg_bank_reg_r31_22_; 
wire REGFILE_SIM_reg_bank_reg_r31_23_; 
wire REGFILE_SIM_reg_bank_reg_r31_24_; 
wire REGFILE_SIM_reg_bank_reg_r31_25_; 
wire REGFILE_SIM_reg_bank_reg_r31_26_; 
wire REGFILE_SIM_reg_bank_reg_r31_27_; 
wire REGFILE_SIM_reg_bank_reg_r31_28_; 
wire REGFILE_SIM_reg_bank_reg_r31_29_; 
wire REGFILE_SIM_reg_bank_reg_r31_2_; 
wire REGFILE_SIM_reg_bank_reg_r31_30_; 
wire REGFILE_SIM_reg_bank_reg_r31_31_; 
wire REGFILE_SIM_reg_bank_reg_r31_3_; 
wire REGFILE_SIM_reg_bank_reg_r31_4_; 
wire REGFILE_SIM_reg_bank_reg_r31_5_; 
wire REGFILE_SIM_reg_bank_reg_r31_6_; 
wire REGFILE_SIM_reg_bank_reg_r31_7_; 
wire REGFILE_SIM_reg_bank_reg_r31_8_; 
wire REGFILE_SIM_reg_bank_reg_r31_9_; 
wire REGFILE_SIM_reg_bank_reg_r3_0_; 
wire REGFILE_SIM_reg_bank_reg_r3_10_; 
wire REGFILE_SIM_reg_bank_reg_r3_11_; 
wire REGFILE_SIM_reg_bank_reg_r3_12_; 
wire REGFILE_SIM_reg_bank_reg_r3_13_; 
wire REGFILE_SIM_reg_bank_reg_r3_14_; 
wire REGFILE_SIM_reg_bank_reg_r3_15_; 
wire REGFILE_SIM_reg_bank_reg_r3_16_; 
wire REGFILE_SIM_reg_bank_reg_r3_17_; 
wire REGFILE_SIM_reg_bank_reg_r3_18_; 
wire REGFILE_SIM_reg_bank_reg_r3_19_; 
wire REGFILE_SIM_reg_bank_reg_r3_1_; 
wire REGFILE_SIM_reg_bank_reg_r3_20_; 
wire REGFILE_SIM_reg_bank_reg_r3_21_; 
wire REGFILE_SIM_reg_bank_reg_r3_22_; 
wire REGFILE_SIM_reg_bank_reg_r3_23_; 
wire REGFILE_SIM_reg_bank_reg_r3_24_; 
wire REGFILE_SIM_reg_bank_reg_r3_25_; 
wire REGFILE_SIM_reg_bank_reg_r3_26_; 
wire REGFILE_SIM_reg_bank_reg_r3_27_; 
wire REGFILE_SIM_reg_bank_reg_r3_28_; 
wire REGFILE_SIM_reg_bank_reg_r3_29_; 
wire REGFILE_SIM_reg_bank_reg_r3_2_; 
wire REGFILE_SIM_reg_bank_reg_r3_30_; 
wire REGFILE_SIM_reg_bank_reg_r3_31_; 
wire REGFILE_SIM_reg_bank_reg_r3_3_; 
wire REGFILE_SIM_reg_bank_reg_r3_4_; 
wire REGFILE_SIM_reg_bank_reg_r3_5_; 
wire REGFILE_SIM_reg_bank_reg_r3_6_; 
wire REGFILE_SIM_reg_bank_reg_r3_7_; 
wire REGFILE_SIM_reg_bank_reg_r3_8_; 
wire REGFILE_SIM_reg_bank_reg_r3_9_; 
wire REGFILE_SIM_reg_bank_reg_r4_0_; 
wire REGFILE_SIM_reg_bank_reg_r4_10_; 
wire REGFILE_SIM_reg_bank_reg_r4_11_; 
wire REGFILE_SIM_reg_bank_reg_r4_12_; 
wire REGFILE_SIM_reg_bank_reg_r4_13_; 
wire REGFILE_SIM_reg_bank_reg_r4_14_; 
wire REGFILE_SIM_reg_bank_reg_r4_15_; 
wire REGFILE_SIM_reg_bank_reg_r4_16_; 
wire REGFILE_SIM_reg_bank_reg_r4_17_; 
wire REGFILE_SIM_reg_bank_reg_r4_18_; 
wire REGFILE_SIM_reg_bank_reg_r4_19_; 
wire REGFILE_SIM_reg_bank_reg_r4_1_; 
wire REGFILE_SIM_reg_bank_reg_r4_20_; 
wire REGFILE_SIM_reg_bank_reg_r4_21_; 
wire REGFILE_SIM_reg_bank_reg_r4_22_; 
wire REGFILE_SIM_reg_bank_reg_r4_23_; 
wire REGFILE_SIM_reg_bank_reg_r4_24_; 
wire REGFILE_SIM_reg_bank_reg_r4_25_; 
wire REGFILE_SIM_reg_bank_reg_r4_26_; 
wire REGFILE_SIM_reg_bank_reg_r4_27_; 
wire REGFILE_SIM_reg_bank_reg_r4_28_; 
wire REGFILE_SIM_reg_bank_reg_r4_29_; 
wire REGFILE_SIM_reg_bank_reg_r4_2_; 
wire REGFILE_SIM_reg_bank_reg_r4_30_; 
wire REGFILE_SIM_reg_bank_reg_r4_31_; 
wire REGFILE_SIM_reg_bank_reg_r4_3_; 
wire REGFILE_SIM_reg_bank_reg_r4_4_; 
wire REGFILE_SIM_reg_bank_reg_r4_5_; 
wire REGFILE_SIM_reg_bank_reg_r4_6_; 
wire REGFILE_SIM_reg_bank_reg_r4_7_; 
wire REGFILE_SIM_reg_bank_reg_r4_8_; 
wire REGFILE_SIM_reg_bank_reg_r4_9_; 
wire REGFILE_SIM_reg_bank_reg_r5_0_; 
wire REGFILE_SIM_reg_bank_reg_r5_10_; 
wire REGFILE_SIM_reg_bank_reg_r5_11_; 
wire REGFILE_SIM_reg_bank_reg_r5_12_; 
wire REGFILE_SIM_reg_bank_reg_r5_13_; 
wire REGFILE_SIM_reg_bank_reg_r5_14_; 
wire REGFILE_SIM_reg_bank_reg_r5_15_; 
wire REGFILE_SIM_reg_bank_reg_r5_16_; 
wire REGFILE_SIM_reg_bank_reg_r5_17_; 
wire REGFILE_SIM_reg_bank_reg_r5_18_; 
wire REGFILE_SIM_reg_bank_reg_r5_19_; 
wire REGFILE_SIM_reg_bank_reg_r5_1_; 
wire REGFILE_SIM_reg_bank_reg_r5_20_; 
wire REGFILE_SIM_reg_bank_reg_r5_21_; 
wire REGFILE_SIM_reg_bank_reg_r5_22_; 
wire REGFILE_SIM_reg_bank_reg_r5_23_; 
wire REGFILE_SIM_reg_bank_reg_r5_24_; 
wire REGFILE_SIM_reg_bank_reg_r5_25_; 
wire REGFILE_SIM_reg_bank_reg_r5_26_; 
wire REGFILE_SIM_reg_bank_reg_r5_27_; 
wire REGFILE_SIM_reg_bank_reg_r5_28_; 
wire REGFILE_SIM_reg_bank_reg_r5_29_; 
wire REGFILE_SIM_reg_bank_reg_r5_2_; 
wire REGFILE_SIM_reg_bank_reg_r5_30_; 
wire REGFILE_SIM_reg_bank_reg_r5_31_; 
wire REGFILE_SIM_reg_bank_reg_r5_3_; 
wire REGFILE_SIM_reg_bank_reg_r5_4_; 
wire REGFILE_SIM_reg_bank_reg_r5_5_; 
wire REGFILE_SIM_reg_bank_reg_r5_6_; 
wire REGFILE_SIM_reg_bank_reg_r5_7_; 
wire REGFILE_SIM_reg_bank_reg_r5_8_; 
wire REGFILE_SIM_reg_bank_reg_r5_9_; 
wire REGFILE_SIM_reg_bank_reg_r6_0_; 
wire REGFILE_SIM_reg_bank_reg_r6_10_; 
wire REGFILE_SIM_reg_bank_reg_r6_11_; 
wire REGFILE_SIM_reg_bank_reg_r6_12_; 
wire REGFILE_SIM_reg_bank_reg_r6_13_; 
wire REGFILE_SIM_reg_bank_reg_r6_14_; 
wire REGFILE_SIM_reg_bank_reg_r6_15_; 
wire REGFILE_SIM_reg_bank_reg_r6_16_; 
wire REGFILE_SIM_reg_bank_reg_r6_17_; 
wire REGFILE_SIM_reg_bank_reg_r6_18_; 
wire REGFILE_SIM_reg_bank_reg_r6_19_; 
wire REGFILE_SIM_reg_bank_reg_r6_1_; 
wire REGFILE_SIM_reg_bank_reg_r6_20_; 
wire REGFILE_SIM_reg_bank_reg_r6_21_; 
wire REGFILE_SIM_reg_bank_reg_r6_22_; 
wire REGFILE_SIM_reg_bank_reg_r6_23_; 
wire REGFILE_SIM_reg_bank_reg_r6_24_; 
wire REGFILE_SIM_reg_bank_reg_r6_25_; 
wire REGFILE_SIM_reg_bank_reg_r6_26_; 
wire REGFILE_SIM_reg_bank_reg_r6_27_; 
wire REGFILE_SIM_reg_bank_reg_r6_28_; 
wire REGFILE_SIM_reg_bank_reg_r6_29_; 
wire REGFILE_SIM_reg_bank_reg_r6_2_; 
wire REGFILE_SIM_reg_bank_reg_r6_30_; 
wire REGFILE_SIM_reg_bank_reg_r6_31_; 
wire REGFILE_SIM_reg_bank_reg_r6_3_; 
wire REGFILE_SIM_reg_bank_reg_r6_4_; 
wire REGFILE_SIM_reg_bank_reg_r6_5_; 
wire REGFILE_SIM_reg_bank_reg_r6_6_; 
wire REGFILE_SIM_reg_bank_reg_r6_7_; 
wire REGFILE_SIM_reg_bank_reg_r6_8_; 
wire REGFILE_SIM_reg_bank_reg_r6_9_; 
wire REGFILE_SIM_reg_bank_reg_r7_0_; 
wire REGFILE_SIM_reg_bank_reg_r7_10_; 
wire REGFILE_SIM_reg_bank_reg_r7_11_; 
wire REGFILE_SIM_reg_bank_reg_r7_12_; 
wire REGFILE_SIM_reg_bank_reg_r7_13_; 
wire REGFILE_SIM_reg_bank_reg_r7_14_; 
wire REGFILE_SIM_reg_bank_reg_r7_15_; 
wire REGFILE_SIM_reg_bank_reg_r7_16_; 
wire REGFILE_SIM_reg_bank_reg_r7_17_; 
wire REGFILE_SIM_reg_bank_reg_r7_18_; 
wire REGFILE_SIM_reg_bank_reg_r7_19_; 
wire REGFILE_SIM_reg_bank_reg_r7_1_; 
wire REGFILE_SIM_reg_bank_reg_r7_20_; 
wire REGFILE_SIM_reg_bank_reg_r7_21_; 
wire REGFILE_SIM_reg_bank_reg_r7_22_; 
wire REGFILE_SIM_reg_bank_reg_r7_23_; 
wire REGFILE_SIM_reg_bank_reg_r7_24_; 
wire REGFILE_SIM_reg_bank_reg_r7_25_; 
wire REGFILE_SIM_reg_bank_reg_r7_26_; 
wire REGFILE_SIM_reg_bank_reg_r7_27_; 
wire REGFILE_SIM_reg_bank_reg_r7_28_; 
wire REGFILE_SIM_reg_bank_reg_r7_29_; 
wire REGFILE_SIM_reg_bank_reg_r7_2_; 
wire REGFILE_SIM_reg_bank_reg_r7_30_; 
wire REGFILE_SIM_reg_bank_reg_r7_31_; 
wire REGFILE_SIM_reg_bank_reg_r7_3_; 
wire REGFILE_SIM_reg_bank_reg_r7_4_; 
wire REGFILE_SIM_reg_bank_reg_r7_5_; 
wire REGFILE_SIM_reg_bank_reg_r7_6_; 
wire REGFILE_SIM_reg_bank_reg_r7_7_; 
wire REGFILE_SIM_reg_bank_reg_r7_8_; 
wire REGFILE_SIM_reg_bank_reg_r7_9_; 
wire REGFILE_SIM_reg_bank_reg_r8_0_; 
wire REGFILE_SIM_reg_bank_reg_r8_10_; 
wire REGFILE_SIM_reg_bank_reg_r8_11_; 
wire REGFILE_SIM_reg_bank_reg_r8_12_; 
wire REGFILE_SIM_reg_bank_reg_r8_13_; 
wire REGFILE_SIM_reg_bank_reg_r8_14_; 
wire REGFILE_SIM_reg_bank_reg_r8_15_; 
wire REGFILE_SIM_reg_bank_reg_r8_16_; 
wire REGFILE_SIM_reg_bank_reg_r8_17_; 
wire REGFILE_SIM_reg_bank_reg_r8_18_; 
wire REGFILE_SIM_reg_bank_reg_r8_19_; 
wire REGFILE_SIM_reg_bank_reg_r8_1_; 
wire REGFILE_SIM_reg_bank_reg_r8_20_; 
wire REGFILE_SIM_reg_bank_reg_r8_21_; 
wire REGFILE_SIM_reg_bank_reg_r8_22_; 
wire REGFILE_SIM_reg_bank_reg_r8_23_; 
wire REGFILE_SIM_reg_bank_reg_r8_24_; 
wire REGFILE_SIM_reg_bank_reg_r8_25_; 
wire REGFILE_SIM_reg_bank_reg_r8_26_; 
wire REGFILE_SIM_reg_bank_reg_r8_27_; 
wire REGFILE_SIM_reg_bank_reg_r8_28_; 
wire REGFILE_SIM_reg_bank_reg_r8_29_; 
wire REGFILE_SIM_reg_bank_reg_r8_2_; 
wire REGFILE_SIM_reg_bank_reg_r8_30_; 
wire REGFILE_SIM_reg_bank_reg_r8_31_; 
wire REGFILE_SIM_reg_bank_reg_r8_3_; 
wire REGFILE_SIM_reg_bank_reg_r8_4_; 
wire REGFILE_SIM_reg_bank_reg_r8_5_; 
wire REGFILE_SIM_reg_bank_reg_r8_6_; 
wire REGFILE_SIM_reg_bank_reg_r8_7_; 
wire REGFILE_SIM_reg_bank_reg_r8_8_; 
wire REGFILE_SIM_reg_bank_reg_r8_9_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_0_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_10_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_11_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_12_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_13_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_14_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_15_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_16_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_17_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_18_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_19_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_1_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_20_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_21_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_22_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_23_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_24_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_25_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_26_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_27_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_28_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_29_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_2_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_30_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_31_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_3_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_4_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_5_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_6_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_7_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_8_; 
wire REGFILE_SIM_reg_bank_reg_r9_lr_9_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_0_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_10_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_11_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_12_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_13_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_14_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_15_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_16_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_17_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_18_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_19_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_1_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_20_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_21_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_22_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_23_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_24_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_25_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_26_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_27_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_28_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_29_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_2_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_30_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_31_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_3_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_4_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_5_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_6_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_7_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_8_; 
wire REGFILE_SIM_reg_bank_reg_ra_o_9_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_0_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_10_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_11_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_12_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_13_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_14_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_15_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_16_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_17_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_18_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_19_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_1_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_20_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_21_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_22_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_23_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_24_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_25_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_26_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_27_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_28_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_29_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_2_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_30_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_31_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_3_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_4_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_5_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_6_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_7_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_8_; 
wire REGFILE_SIM_reg_bank_reg_rb_o_9_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_10_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_11_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_12_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_13_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_14_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_15_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_16_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_17_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_18_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_19_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_20_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_21_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_22_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_23_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_24_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_25_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_26_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_27_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_28_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_29_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_30_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_31_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_4_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_5_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_6_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_7_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_8_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_9_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_; 
wire REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_; 
wire REGFILE_SIM_reg_bank_wr_i; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf0; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf1; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf2; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf3; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf4; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf5; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf6; 
wire REGFILE_SIM_reg_bank_wr_i_bF_buf7; 
wire _0epc_q_31_0__0_; 
wire _0epc_q_31_0__10_; 
wire _0epc_q_31_0__11_; 
wire _0epc_q_31_0__12_; 
wire _0epc_q_31_0__13_; 
wire _0epc_q_31_0__14_; 
wire _0epc_q_31_0__15_; 
wire _0epc_q_31_0__16_; 
wire _0epc_q_31_0__17_; 
wire _0epc_q_31_0__18_; 
wire _0epc_q_31_0__19_; 
wire _0epc_q_31_0__1_; 
wire _0epc_q_31_0__20_; 
wire _0epc_q_31_0__21_; 
wire _0epc_q_31_0__22_; 
wire _0epc_q_31_0__23_; 
wire _0epc_q_31_0__24_; 
wire _0epc_q_31_0__25_; 
wire _0epc_q_31_0__26_; 
wire _0epc_q_31_0__27_; 
wire _0epc_q_31_0__28_; 
wire _0epc_q_31_0__29_; 
wire _0epc_q_31_0__2_; 
wire _0epc_q_31_0__30_; 
wire _0epc_q_31_0__31_; 
wire _0epc_q_31_0__3_; 
wire _0epc_q_31_0__4_; 
wire _0epc_q_31_0__5_; 
wire _0epc_q_31_0__6_; 
wire _0epc_q_31_0__7_; 
wire _0epc_q_31_0__8_; 
wire _0epc_q_31_0__9_; 
wire _0esr_q_31_0__10_; 
wire _0esr_q_31_0__2_; 
wire _0esr_q_31_0__9_; 
wire _0ex_rd_q_4_0__0_; 
wire _0ex_rd_q_4_0__1_; 
wire _0ex_rd_q_4_0__2_; 
wire _0ex_rd_q_4_0__3_; 
wire _0ex_rd_q_4_0__4_; 
wire _0fault_o_0_0_; 
wire _0mem_addr_o_31_0__0_; 
wire _0mem_addr_o_31_0__10_; 
wire _0mem_addr_o_31_0__11_; 
wire _0mem_addr_o_31_0__12_; 
wire _0mem_addr_o_31_0__13_; 
wire _0mem_addr_o_31_0__14_; 
wire _0mem_addr_o_31_0__15_; 
wire _0mem_addr_o_31_0__16_; 
wire _0mem_addr_o_31_0__17_; 
wire _0mem_addr_o_31_0__18_; 
wire _0mem_addr_o_31_0__19_; 
wire _0mem_addr_o_31_0__1_; 
wire _0mem_addr_o_31_0__20_; 
wire _0mem_addr_o_31_0__21_; 
wire _0mem_addr_o_31_0__22_; 
wire _0mem_addr_o_31_0__23_; 
wire _0mem_addr_o_31_0__24_; 
wire _0mem_addr_o_31_0__25_; 
wire _0mem_addr_o_31_0__26_; 
wire _0mem_addr_o_31_0__27_; 
wire _0mem_addr_o_31_0__28_; 
wire _0mem_addr_o_31_0__29_; 
wire _0mem_addr_o_31_0__2_; 
wire _0mem_addr_o_31_0__30_; 
wire _0mem_addr_o_31_0__31_; 
wire _0mem_addr_o_31_0__3_; 
wire _0mem_addr_o_31_0__4_; 
wire _0mem_addr_o_31_0__5_; 
wire _0mem_addr_o_31_0__6_; 
wire _0mem_addr_o_31_0__7_; 
wire _0mem_addr_o_31_0__8_; 
wire _0mem_addr_o_31_0__9_; 
wire _0mem_cyc_o_0_0_; 
wire _0mem_dat_o_31_0__0_; 
wire _0mem_dat_o_31_0__10_; 
wire _0mem_dat_o_31_0__11_; 
wire _0mem_dat_o_31_0__12_; 
wire _0mem_dat_o_31_0__13_; 
wire _0mem_dat_o_31_0__14_; 
wire _0mem_dat_o_31_0__15_; 
wire _0mem_dat_o_31_0__16_; 
wire _0mem_dat_o_31_0__17_; 
wire _0mem_dat_o_31_0__18_; 
wire _0mem_dat_o_31_0__19_; 
wire _0mem_dat_o_31_0__1_; 
wire _0mem_dat_o_31_0__20_; 
wire _0mem_dat_o_31_0__21_; 
wire _0mem_dat_o_31_0__22_; 
wire _0mem_dat_o_31_0__23_; 
wire _0mem_dat_o_31_0__24_; 
wire _0mem_dat_o_31_0__25_; 
wire _0mem_dat_o_31_0__26_; 
wire _0mem_dat_o_31_0__27_; 
wire _0mem_dat_o_31_0__28_; 
wire _0mem_dat_o_31_0__29_; 
wire _0mem_dat_o_31_0__2_; 
wire _0mem_dat_o_31_0__30_; 
wire _0mem_dat_o_31_0__31_; 
wire _0mem_dat_o_31_0__3_; 
wire _0mem_dat_o_31_0__4_; 
wire _0mem_dat_o_31_0__5_; 
wire _0mem_dat_o_31_0__6_; 
wire _0mem_dat_o_31_0__7_; 
wire _0mem_dat_o_31_0__8_; 
wire _0mem_dat_o_31_0__9_; 
wire _0mem_offset_q_1_0__0_; 
wire _0mem_offset_q_1_0__1_; 
wire _0mem_sel_o_3_0__0_; 
wire _0mem_sel_o_3_0__1_; 
wire _0mem_sel_o_3_0__2_; 
wire _0mem_sel_o_3_0__3_; 
wire _0mem_stb_o_0_0_; 
wire _0mem_we_o_0_0_; 
wire _0nmi_q_0_0_; 
wire _0opcode_q_31_0__0_; 
wire _0opcode_q_31_0__10_; 
wire _0opcode_q_31_0__11_; 
wire _0opcode_q_31_0__12_; 
wire _0opcode_q_31_0__13_; 
wire _0opcode_q_31_0__14_; 
wire _0opcode_q_31_0__15_; 
wire _0opcode_q_31_0__16_; 
wire _0opcode_q_31_0__17_; 
wire _0opcode_q_31_0__18_; 
wire _0opcode_q_31_0__19_; 
wire _0opcode_q_31_0__1_; 
wire _0opcode_q_31_0__20_; 
wire _0opcode_q_31_0__21_; 
wire _0opcode_q_31_0__22_; 
wire _0opcode_q_31_0__23_; 
wire _0opcode_q_31_0__24_; 
wire _0opcode_q_31_0__25_; 
wire _0opcode_q_31_0__26_; 
wire _0opcode_q_31_0__27_; 
wire _0opcode_q_31_0__28_; 
wire _0opcode_q_31_0__29_; 
wire _0opcode_q_31_0__2_; 
wire _0opcode_q_31_0__30_; 
wire _0opcode_q_31_0__31_; 
wire _0opcode_q_31_0__3_; 
wire _0opcode_q_31_0__4_; 
wire _0opcode_q_31_0__5_; 
wire _0opcode_q_31_0__6_; 
wire _0opcode_q_31_0__7_; 
wire _0opcode_q_31_0__8_; 
wire _0opcode_q_31_0__9_; 
wire _0pc_q_31_0__0_; 
wire _0pc_q_31_0__10_; 
wire _0pc_q_31_0__11_; 
wire _0pc_q_31_0__12_; 
wire _0pc_q_31_0__13_; 
wire _0pc_q_31_0__14_; 
wire _0pc_q_31_0__15_; 
wire _0pc_q_31_0__16_; 
wire _0pc_q_31_0__17_; 
wire _0pc_q_31_0__18_; 
wire _0pc_q_31_0__19_; 
wire _0pc_q_31_0__1_; 
wire _0pc_q_31_0__20_; 
wire _0pc_q_31_0__21_; 
wire _0pc_q_31_0__22_; 
wire _0pc_q_31_0__23_; 
wire _0pc_q_31_0__24_; 
wire _0pc_q_31_0__25_; 
wire _0pc_q_31_0__26_; 
wire _0pc_q_31_0__27_; 
wire _0pc_q_31_0__28_; 
wire _0pc_q_31_0__29_; 
wire _0pc_q_31_0__2_; 
wire _0pc_q_31_0__30_; 
wire _0pc_q_31_0__31_; 
wire _0pc_q_31_0__3_; 
wire _0pc_q_31_0__4_; 
wire _0pc_q_31_0__5_; 
wire _0pc_q_31_0__6_; 
wire _0pc_q_31_0__7_; 
wire _0pc_q_31_0__8_; 
wire _0pc_q_31_0__9_; 
wire _0sr_q_31_0__10_; 
wire _0sr_q_31_0__2_; 
wire _0sr_q_31_0__9_; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2386; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6; 
wire _abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7; 
wire _abc_28031_auto_fsm_map_cc_170_map_fsm_2380_1_; 
wire _abc_28031_auto_fsm_map_cc_170_map_fsm_2380_2_; 
wire _abc_28031_auto_fsm_map_cc_170_map_fsm_2380_3_; 
wire _abc_28031_auto_fsm_map_cc_170_map_fsm_2380_4_; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf0; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf1; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf2; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8; 
wire _abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9; 
wire _abc_44694_new_n1000_; 
wire _abc_44694_new_n1001_; 
wire _abc_44694_new_n1002_; 
wire _abc_44694_new_n1003_; 
wire _abc_44694_new_n1004_; 
wire _abc_44694_new_n1005_; 
wire _abc_44694_new_n1006_; 
wire _abc_44694_new_n1007_; 
wire _abc_44694_new_n1008_; 
wire _abc_44694_new_n1009_; 
wire _abc_44694_new_n1010_; 
wire _abc_44694_new_n1011_; 
wire _abc_44694_new_n1012_; 
wire _abc_44694_new_n1013_; 
wire _abc_44694_new_n1014_; 
wire _abc_44694_new_n1015_; 
wire _abc_44694_new_n1016_; 
wire _abc_44694_new_n1017_; 
wire _abc_44694_new_n1018_; 
wire _abc_44694_new_n1019_; 
wire _abc_44694_new_n1019__bF_buf0; 
wire _abc_44694_new_n1019__bF_buf1; 
wire _abc_44694_new_n1019__bF_buf2; 
wire _abc_44694_new_n1019__bF_buf3; 
wire _abc_44694_new_n1019__bF_buf4; 
wire _abc_44694_new_n1020_; 
wire _abc_44694_new_n1021_; 
wire _abc_44694_new_n1022_; 
wire _abc_44694_new_n1023_; 
wire _abc_44694_new_n1024_; 
wire _abc_44694_new_n1025_; 
wire _abc_44694_new_n1026_; 
wire _abc_44694_new_n1027_; 
wire _abc_44694_new_n1028_; 
wire _abc_44694_new_n1029_; 
wire _abc_44694_new_n1030_; 
wire _abc_44694_new_n1031_; 
wire _abc_44694_new_n1032_; 
wire _abc_44694_new_n1033_; 
wire _abc_44694_new_n1034_; 
wire _abc_44694_new_n1035_; 
wire _abc_44694_new_n1036_; 
wire _abc_44694_new_n1037_; 
wire _abc_44694_new_n1038_; 
wire _abc_44694_new_n1039_; 
wire _abc_44694_new_n1040_; 
wire _abc_44694_new_n1041_; 
wire _abc_44694_new_n1042_; 
wire _abc_44694_new_n1043_; 
wire _abc_44694_new_n1044_; 
wire _abc_44694_new_n1045_; 
wire _abc_44694_new_n1046_; 
wire _abc_44694_new_n1047_; 
wire _abc_44694_new_n1048_; 
wire _abc_44694_new_n1049_; 
wire _abc_44694_new_n1050_; 
wire _abc_44694_new_n1051_; 
wire _abc_44694_new_n1052_; 
wire _abc_44694_new_n1053_; 
wire _abc_44694_new_n1054_; 
wire _abc_44694_new_n1055_; 
wire _abc_44694_new_n1056_; 
wire _abc_44694_new_n1057_; 
wire _abc_44694_new_n1058_; 
wire _abc_44694_new_n1059_; 
wire _abc_44694_new_n1060_; 
wire _abc_44694_new_n1061_; 
wire _abc_44694_new_n1062_; 
wire _abc_44694_new_n1063_; 
wire _abc_44694_new_n1064_; 
wire _abc_44694_new_n1065_; 
wire _abc_44694_new_n1066_; 
wire _abc_44694_new_n1067_; 
wire _abc_44694_new_n1068_; 
wire _abc_44694_new_n1069_; 
wire _abc_44694_new_n1070_; 
wire _abc_44694_new_n1071_; 
wire _abc_44694_new_n1072_; 
wire _abc_44694_new_n1073_; 
wire _abc_44694_new_n1074_; 
wire _abc_44694_new_n1075_; 
wire _abc_44694_new_n1076_; 
wire _abc_44694_new_n1077_; 
wire _abc_44694_new_n1078_; 
wire _abc_44694_new_n1079_; 
wire _abc_44694_new_n1080_; 
wire _abc_44694_new_n1081_; 
wire _abc_44694_new_n1082_; 
wire _abc_44694_new_n1083_; 
wire _abc_44694_new_n1084_; 
wire _abc_44694_new_n1084__bF_buf0; 
wire _abc_44694_new_n1084__bF_buf1; 
wire _abc_44694_new_n1084__bF_buf2; 
wire _abc_44694_new_n1084__bF_buf3; 
wire _abc_44694_new_n1085_; 
wire _abc_44694_new_n1086_; 
wire _abc_44694_new_n1087_; 
wire _abc_44694_new_n1087__bF_buf0; 
wire _abc_44694_new_n1087__bF_buf1; 
wire _abc_44694_new_n1087__bF_buf2; 
wire _abc_44694_new_n1087__bF_buf3; 
wire _abc_44694_new_n1088_; 
wire _abc_44694_new_n1089_; 
wire _abc_44694_new_n1090_; 
wire _abc_44694_new_n1091_; 
wire _abc_44694_new_n1092_; 
wire _abc_44694_new_n1093_; 
wire _abc_44694_new_n1094_; 
wire _abc_44694_new_n1095_; 
wire _abc_44694_new_n1096_; 
wire _abc_44694_new_n1097_; 
wire _abc_44694_new_n1098_; 
wire _abc_44694_new_n1099_; 
wire _abc_44694_new_n1100_; 
wire _abc_44694_new_n1101_; 
wire _abc_44694_new_n1102_; 
wire _abc_44694_new_n1103_; 
wire _abc_44694_new_n1104_; 
wire _abc_44694_new_n1105_; 
wire _abc_44694_new_n1106_; 
wire _abc_44694_new_n1107_; 
wire _abc_44694_new_n1108_; 
wire _abc_44694_new_n1109_; 
wire _abc_44694_new_n1110_; 
wire _abc_44694_new_n1111_; 
wire _abc_44694_new_n1112_; 
wire _abc_44694_new_n1113_; 
wire _abc_44694_new_n1114_; 
wire _abc_44694_new_n1114__bF_buf0; 
wire _abc_44694_new_n1114__bF_buf1; 
wire _abc_44694_new_n1114__bF_buf2; 
wire _abc_44694_new_n1114__bF_buf3; 
wire _abc_44694_new_n1114__bF_buf4; 
wire _abc_44694_new_n1115_; 
wire _abc_44694_new_n1116_; 
wire _abc_44694_new_n1117_; 
wire _abc_44694_new_n1118_; 
wire _abc_44694_new_n1119_; 
wire _abc_44694_new_n1120_; 
wire _abc_44694_new_n1121_; 
wire _abc_44694_new_n1122_; 
wire _abc_44694_new_n1123_; 
wire _abc_44694_new_n1124_; 
wire _abc_44694_new_n1125_; 
wire _abc_44694_new_n1126_; 
wire _abc_44694_new_n1127_; 
wire _abc_44694_new_n1128_; 
wire _abc_44694_new_n1129_; 
wire _abc_44694_new_n1130_; 
wire _abc_44694_new_n1131_; 
wire _abc_44694_new_n1132_; 
wire _abc_44694_new_n1133_; 
wire _abc_44694_new_n1134_; 
wire _abc_44694_new_n1135_; 
wire _abc_44694_new_n1136_; 
wire _abc_44694_new_n1137_; 
wire _abc_44694_new_n1138_; 
wire _abc_44694_new_n1139_; 
wire _abc_44694_new_n1140_; 
wire _abc_44694_new_n1141_; 
wire _abc_44694_new_n1142_; 
wire _abc_44694_new_n1143_; 
wire _abc_44694_new_n1144_; 
wire _abc_44694_new_n1145_; 
wire _abc_44694_new_n1146_; 
wire _abc_44694_new_n1147_; 
wire _abc_44694_new_n1148_; 
wire _abc_44694_new_n1149_; 
wire _abc_44694_new_n1150_; 
wire _abc_44694_new_n1151_; 
wire _abc_44694_new_n1152_; 
wire _abc_44694_new_n1153_; 
wire _abc_44694_new_n1154_; 
wire _abc_44694_new_n1155_; 
wire _abc_44694_new_n1156_; 
wire _abc_44694_new_n1157_; 
wire _abc_44694_new_n1158_; 
wire _abc_44694_new_n1159_; 
wire _abc_44694_new_n1160_; 
wire _abc_44694_new_n1161_; 
wire _abc_44694_new_n1162_; 
wire _abc_44694_new_n1163_; 
wire _abc_44694_new_n1164_; 
wire _abc_44694_new_n1165_; 
wire _abc_44694_new_n1166_; 
wire _abc_44694_new_n1167_; 
wire _abc_44694_new_n1168_; 
wire _abc_44694_new_n1169_; 
wire _abc_44694_new_n1170_; 
wire _abc_44694_new_n1171_; 
wire _abc_44694_new_n1172_; 
wire _abc_44694_new_n1173_; 
wire _abc_44694_new_n1174_; 
wire _abc_44694_new_n1175_; 
wire _abc_44694_new_n1176_; 
wire _abc_44694_new_n1177_; 
wire _abc_44694_new_n1178_; 
wire _abc_44694_new_n1178__bF_buf0; 
wire _abc_44694_new_n1178__bF_buf1; 
wire _abc_44694_new_n1178__bF_buf2; 
wire _abc_44694_new_n1178__bF_buf3; 
wire _abc_44694_new_n1178__bF_buf4; 
wire _abc_44694_new_n1179_; 
wire _abc_44694_new_n1179__bF_buf0; 
wire _abc_44694_new_n1179__bF_buf1; 
wire _abc_44694_new_n1179__bF_buf2; 
wire _abc_44694_new_n1179__bF_buf3; 
wire _abc_44694_new_n1180_; 
wire _abc_44694_new_n1181_; 
wire _abc_44694_new_n1181__bF_buf0; 
wire _abc_44694_new_n1181__bF_buf1; 
wire _abc_44694_new_n1181__bF_buf2; 
wire _abc_44694_new_n1181__bF_buf3; 
wire _abc_44694_new_n1182_; 
wire _abc_44694_new_n1183_; 
wire _abc_44694_new_n1184_; 
wire _abc_44694_new_n1185_; 
wire _abc_44694_new_n1185__bF_buf0; 
wire _abc_44694_new_n1185__bF_buf1; 
wire _abc_44694_new_n1185__bF_buf2; 
wire _abc_44694_new_n1185__bF_buf3; 
wire _abc_44694_new_n1186_; 
wire _abc_44694_new_n1186__bF_buf0; 
wire _abc_44694_new_n1186__bF_buf1; 
wire _abc_44694_new_n1186__bF_buf2; 
wire _abc_44694_new_n1186__bF_buf3; 
wire _abc_44694_new_n1187_; 
wire _abc_44694_new_n1188_; 
wire _abc_44694_new_n1189_; 
wire _abc_44694_new_n1190_; 
wire _abc_44694_new_n1191_; 
wire _abc_44694_new_n1192_; 
wire _abc_44694_new_n1193_; 
wire _abc_44694_new_n1194_; 
wire _abc_44694_new_n1194__bF_buf0; 
wire _abc_44694_new_n1194__bF_buf1; 
wire _abc_44694_new_n1194__bF_buf2; 
wire _abc_44694_new_n1194__bF_buf3; 
wire _abc_44694_new_n1194__bF_buf4; 
wire _abc_44694_new_n1195_; 
wire _abc_44694_new_n1196_; 
wire _abc_44694_new_n1197_; 
wire _abc_44694_new_n1198_; 
wire _abc_44694_new_n1199_; 
wire _abc_44694_new_n1200_; 
wire _abc_44694_new_n1201_; 
wire _abc_44694_new_n1202_; 
wire _abc_44694_new_n1203_; 
wire _abc_44694_new_n1204_; 
wire _abc_44694_new_n1205_; 
wire _abc_44694_new_n1206_; 
wire _abc_44694_new_n1207_; 
wire _abc_44694_new_n1207__bF_buf0; 
wire _abc_44694_new_n1207__bF_buf1; 
wire _abc_44694_new_n1207__bF_buf2; 
wire _abc_44694_new_n1207__bF_buf3; 
wire _abc_44694_new_n1207__bF_buf4; 
wire _abc_44694_new_n1207__bF_buf5; 
wire _abc_44694_new_n1208_; 
wire _abc_44694_new_n1209_; 
wire _abc_44694_new_n1210_; 
wire _abc_44694_new_n1210__bF_buf0; 
wire _abc_44694_new_n1210__bF_buf1; 
wire _abc_44694_new_n1210__bF_buf2; 
wire _abc_44694_new_n1210__bF_buf3; 
wire _abc_44694_new_n1210__bF_buf4; 
wire _abc_44694_new_n1210__bF_buf5; 
wire _abc_44694_new_n1210__bF_buf6; 
wire _abc_44694_new_n1210__bF_buf7; 
wire _abc_44694_new_n1211_; 
wire _abc_44694_new_n1212_; 
wire _abc_44694_new_n1213_; 
wire _abc_44694_new_n1214_; 
wire _abc_44694_new_n1215_; 
wire _abc_44694_new_n1216_; 
wire _abc_44694_new_n1218_; 
wire _abc_44694_new_n1219_; 
wire _abc_44694_new_n1220_; 
wire _abc_44694_new_n1221_; 
wire _abc_44694_new_n1222_; 
wire _abc_44694_new_n1223_; 
wire _abc_44694_new_n1224_; 
wire _abc_44694_new_n1225_; 
wire _abc_44694_new_n1226_; 
wire _abc_44694_new_n1227_; 
wire _abc_44694_new_n1228_; 
wire _abc_44694_new_n1229_; 
wire _abc_44694_new_n1230_; 
wire _abc_44694_new_n1231_; 
wire _abc_44694_new_n1232_; 
wire _abc_44694_new_n1233_; 
wire _abc_44694_new_n1234_; 
wire _abc_44694_new_n1235_; 
wire _abc_44694_new_n1236_; 
wire _abc_44694_new_n1237_; 
wire _abc_44694_new_n1238_; 
wire _abc_44694_new_n1239_; 
wire _abc_44694_new_n1240_; 
wire _abc_44694_new_n1241_; 
wire _abc_44694_new_n1242_; 
wire _abc_44694_new_n1243_; 
wire _abc_44694_new_n1244_; 
wire _abc_44694_new_n1245_; 
wire _abc_44694_new_n1246_; 
wire _abc_44694_new_n1247_; 
wire _abc_44694_new_n1248_; 
wire _abc_44694_new_n1249_; 
wire _abc_44694_new_n1250_; 
wire _abc_44694_new_n1251_; 
wire _abc_44694_new_n1252_; 
wire _abc_44694_new_n1253_; 
wire _abc_44694_new_n1254_; 
wire _abc_44694_new_n1255_; 
wire _abc_44694_new_n1256_; 
wire _abc_44694_new_n1257_; 
wire _abc_44694_new_n1258_; 
wire _abc_44694_new_n1259_; 
wire _abc_44694_new_n1260_; 
wire _abc_44694_new_n1261_; 
wire _abc_44694_new_n1262_; 
wire _abc_44694_new_n1263_; 
wire _abc_44694_new_n1264_; 
wire _abc_44694_new_n1265_; 
wire _abc_44694_new_n1266_; 
wire _abc_44694_new_n1267_; 
wire _abc_44694_new_n1268_; 
wire _abc_44694_new_n1269_; 
wire _abc_44694_new_n1270_; 
wire _abc_44694_new_n1271_; 
wire _abc_44694_new_n1272_; 
wire _abc_44694_new_n1273_; 
wire _abc_44694_new_n1274_; 
wire _abc_44694_new_n1275_; 
wire _abc_44694_new_n1276_; 
wire _abc_44694_new_n1277_; 
wire _abc_44694_new_n1278_; 
wire _abc_44694_new_n1278__bF_buf0; 
wire _abc_44694_new_n1278__bF_buf1; 
wire _abc_44694_new_n1278__bF_buf2; 
wire _abc_44694_new_n1278__bF_buf3; 
wire _abc_44694_new_n1278__bF_buf4; 
wire _abc_44694_new_n1278__bF_buf5; 
wire _abc_44694_new_n1279_; 
wire _abc_44694_new_n1280_; 
wire _abc_44694_new_n1281_; 
wire _abc_44694_new_n1282_; 
wire _abc_44694_new_n1283_; 
wire _abc_44694_new_n1284_; 
wire _abc_44694_new_n1285_; 
wire _abc_44694_new_n1286_; 
wire _abc_44694_new_n1287_; 
wire _abc_44694_new_n1288_; 
wire _abc_44694_new_n1289_; 
wire _abc_44694_new_n1291_; 
wire _abc_44694_new_n1292_; 
wire _abc_44694_new_n1293_; 
wire _abc_44694_new_n1294_; 
wire _abc_44694_new_n1295_; 
wire _abc_44694_new_n1296_; 
wire _abc_44694_new_n1297_; 
wire _abc_44694_new_n1298_; 
wire _abc_44694_new_n1299_; 
wire _abc_44694_new_n1300_; 
wire _abc_44694_new_n1301_; 
wire _abc_44694_new_n1302_; 
wire _abc_44694_new_n1303_; 
wire _abc_44694_new_n1304_; 
wire _abc_44694_new_n1305_; 
wire _abc_44694_new_n1306_; 
wire _abc_44694_new_n1307_; 
wire _abc_44694_new_n1308_; 
wire _abc_44694_new_n1309_; 
wire _abc_44694_new_n1310_; 
wire _abc_44694_new_n1311_; 
wire _abc_44694_new_n1312_; 
wire _abc_44694_new_n1313_; 
wire _abc_44694_new_n1314_; 
wire _abc_44694_new_n1316_; 
wire _abc_44694_new_n1317_; 
wire _abc_44694_new_n1318_; 
wire _abc_44694_new_n1319_; 
wire _abc_44694_new_n1320_; 
wire _abc_44694_new_n1321_; 
wire _abc_44694_new_n1323_; 
wire _abc_44694_new_n1324_; 
wire _abc_44694_new_n1325_; 
wire _abc_44694_new_n1326_; 
wire _abc_44694_new_n1328_; 
wire _abc_44694_new_n1329_; 
wire _abc_44694_new_n1330_; 
wire _abc_44694_new_n1331_; 
wire _abc_44694_new_n1332_; 
wire _abc_44694_new_n1334_; 
wire _abc_44694_new_n1334__bF_buf0; 
wire _abc_44694_new_n1334__bF_buf1; 
wire _abc_44694_new_n1334__bF_buf2; 
wire _abc_44694_new_n1334__bF_buf3; 
wire _abc_44694_new_n1334__bF_buf4; 
wire _abc_44694_new_n1335_; 
wire _abc_44694_new_n1336_; 
wire _abc_44694_new_n1337_; 
wire _abc_44694_new_n1337__bF_buf0; 
wire _abc_44694_new_n1337__bF_buf1; 
wire _abc_44694_new_n1337__bF_buf2; 
wire _abc_44694_new_n1337__bF_buf3; 
wire _abc_44694_new_n1337__bF_buf4; 
wire _abc_44694_new_n1338_; 
wire _abc_44694_new_n1339_; 
wire _abc_44694_new_n1340_; 
wire _abc_44694_new_n1340__bF_buf0; 
wire _abc_44694_new_n1340__bF_buf1; 
wire _abc_44694_new_n1340__bF_buf2; 
wire _abc_44694_new_n1340__bF_buf3; 
wire _abc_44694_new_n1340__bF_buf4; 
wire _abc_44694_new_n1341_; 
wire _abc_44694_new_n1342_; 
wire _abc_44694_new_n1343_; 
wire _abc_44694_new_n1344_; 
wire _abc_44694_new_n1345_; 
wire _abc_44694_new_n1346_; 
wire _abc_44694_new_n1347_; 
wire _abc_44694_new_n1347__bF_buf0; 
wire _abc_44694_new_n1347__bF_buf1; 
wire _abc_44694_new_n1347__bF_buf2; 
wire _abc_44694_new_n1347__bF_buf3; 
wire _abc_44694_new_n1347__bF_buf4; 
wire _abc_44694_new_n1348_; 
wire _abc_44694_new_n1348__bF_buf0; 
wire _abc_44694_new_n1348__bF_buf1; 
wire _abc_44694_new_n1348__bF_buf2; 
wire _abc_44694_new_n1348__bF_buf3; 
wire _abc_44694_new_n1348__bF_buf4; 
wire _abc_44694_new_n1348__bF_buf5; 
wire _abc_44694_new_n1349_; 
wire _abc_44694_new_n1350_; 
wire _abc_44694_new_n1351_; 
wire _abc_44694_new_n1352_; 
wire _abc_44694_new_n1353_; 
wire _abc_44694_new_n1354_; 
wire _abc_44694_new_n1355_; 
wire _abc_44694_new_n1356_; 
wire _abc_44694_new_n1357_; 
wire _abc_44694_new_n1358_; 
wire _abc_44694_new_n1359_; 
wire _abc_44694_new_n1360_; 
wire _abc_44694_new_n1362_; 
wire _abc_44694_new_n1363_; 
wire _abc_44694_new_n1364_; 
wire _abc_44694_new_n1365_; 
wire _abc_44694_new_n1366_; 
wire _abc_44694_new_n1367_; 
wire _abc_44694_new_n1368_; 
wire _abc_44694_new_n1369_; 
wire _abc_44694_new_n1370_; 
wire _abc_44694_new_n1371_; 
wire _abc_44694_new_n1372_; 
wire _abc_44694_new_n1373_; 
wire _abc_44694_new_n1374_; 
wire _abc_44694_new_n1375_; 
wire _abc_44694_new_n1376_; 
wire _abc_44694_new_n1377_; 
wire _abc_44694_new_n1378_; 
wire _abc_44694_new_n1379_; 
wire _abc_44694_new_n1380_; 
wire _abc_44694_new_n1382_; 
wire _abc_44694_new_n1382__bF_buf0; 
wire _abc_44694_new_n1382__bF_buf1; 
wire _abc_44694_new_n1382__bF_buf2; 
wire _abc_44694_new_n1382__bF_buf3; 
wire _abc_44694_new_n1383_; 
wire _abc_44694_new_n1384_; 
wire _abc_44694_new_n1385_; 
wire _abc_44694_new_n1386_; 
wire _abc_44694_new_n1387_; 
wire _abc_44694_new_n1388_; 
wire _abc_44694_new_n1389_; 
wire _abc_44694_new_n1390_; 
wire _abc_44694_new_n1391_; 
wire _abc_44694_new_n1392_; 
wire _abc_44694_new_n1393_; 
wire _abc_44694_new_n1394_; 
wire _abc_44694_new_n1395_; 
wire _abc_44694_new_n1396_; 
wire _abc_44694_new_n1397_; 
wire _abc_44694_new_n1398_; 
wire _abc_44694_new_n1399_; 
wire _abc_44694_new_n1399__bF_buf0; 
wire _abc_44694_new_n1399__bF_buf1; 
wire _abc_44694_new_n1399__bF_buf2; 
wire _abc_44694_new_n1399__bF_buf3; 
wire _abc_44694_new_n1399__bF_buf4; 
wire _abc_44694_new_n1400_; 
wire _abc_44694_new_n1400__bF_buf0; 
wire _abc_44694_new_n1400__bF_buf1; 
wire _abc_44694_new_n1400__bF_buf2; 
wire _abc_44694_new_n1400__bF_buf3; 
wire _abc_44694_new_n1400__bF_buf4; 
wire _abc_44694_new_n1401_; 
wire _abc_44694_new_n1402_; 
wire _abc_44694_new_n1403_; 
wire _abc_44694_new_n1404_; 
wire _abc_44694_new_n1405_; 
wire _abc_44694_new_n1406_; 
wire _abc_44694_new_n1407_; 
wire _abc_44694_new_n1408_; 
wire _abc_44694_new_n1409_; 
wire _abc_44694_new_n1410_; 
wire _abc_44694_new_n1411_; 
wire _abc_44694_new_n1412_; 
wire _abc_44694_new_n1413_; 
wire _abc_44694_new_n1414_; 
wire _abc_44694_new_n1415_; 
wire _abc_44694_new_n1416_; 
wire _abc_44694_new_n1417_; 
wire _abc_44694_new_n1418_; 
wire _abc_44694_new_n1419_; 
wire _abc_44694_new_n1420_; 
wire _abc_44694_new_n1421_; 
wire _abc_44694_new_n1422_; 
wire _abc_44694_new_n1424_; 
wire _abc_44694_new_n1425_; 
wire _abc_44694_new_n1426_; 
wire _abc_44694_new_n1427_; 
wire _abc_44694_new_n1428_; 
wire _abc_44694_new_n1429_; 
wire _abc_44694_new_n1430_; 
wire _abc_44694_new_n1431_; 
wire _abc_44694_new_n1432_; 
wire _abc_44694_new_n1433_; 
wire _abc_44694_new_n1434_; 
wire _abc_44694_new_n1435_; 
wire _abc_44694_new_n1436_; 
wire _abc_44694_new_n1437_; 
wire _abc_44694_new_n1438_; 
wire _abc_44694_new_n1439_; 
wire _abc_44694_new_n1440_; 
wire _abc_44694_new_n1441_; 
wire _abc_44694_new_n1442_; 
wire _abc_44694_new_n1443_; 
wire _abc_44694_new_n1444_; 
wire _abc_44694_new_n1445_; 
wire _abc_44694_new_n1446_; 
wire _abc_44694_new_n1447_; 
wire _abc_44694_new_n1448_; 
wire _abc_44694_new_n1449_; 
wire _abc_44694_new_n1450_; 
wire _abc_44694_new_n1451_; 
wire _abc_44694_new_n1452_; 
wire _abc_44694_new_n1453_; 
wire _abc_44694_new_n1454_; 
wire _abc_44694_new_n1455_; 
wire _abc_44694_new_n1456_; 
wire _abc_44694_new_n1457_; 
wire _abc_44694_new_n1458_; 
wire _abc_44694_new_n1460_; 
wire _abc_44694_new_n1461_; 
wire _abc_44694_new_n1462_; 
wire _abc_44694_new_n1463_; 
wire _abc_44694_new_n1464_; 
wire _abc_44694_new_n1465_; 
wire _abc_44694_new_n1466_; 
wire _abc_44694_new_n1467_; 
wire _abc_44694_new_n1468_; 
wire _abc_44694_new_n1469_; 
wire _abc_44694_new_n1470_; 
wire _abc_44694_new_n1471_; 
wire _abc_44694_new_n1472_; 
wire _abc_44694_new_n1473_; 
wire _abc_44694_new_n1474_; 
wire _abc_44694_new_n1475_; 
wire _abc_44694_new_n1476_; 
wire _abc_44694_new_n1477_; 
wire _abc_44694_new_n1478_; 
wire _abc_44694_new_n1479_; 
wire _abc_44694_new_n1480_; 
wire _abc_44694_new_n1481_; 
wire _abc_44694_new_n1482_; 
wire _abc_44694_new_n1483_; 
wire _abc_44694_new_n1484_; 
wire _abc_44694_new_n1485_; 
wire _abc_44694_new_n1486_; 
wire _abc_44694_new_n1487_; 
wire _abc_44694_new_n1488_; 
wire _abc_44694_new_n1489_; 
wire _abc_44694_new_n1490_; 
wire _abc_44694_new_n1491_; 
wire _abc_44694_new_n1492_; 
wire _abc_44694_new_n1493_; 
wire _abc_44694_new_n1494_; 
wire _abc_44694_new_n1495_; 
wire _abc_44694_new_n1496_; 
wire _abc_44694_new_n1498_; 
wire _abc_44694_new_n1499_; 
wire _abc_44694_new_n1500_; 
wire _abc_44694_new_n1501_; 
wire _abc_44694_new_n1502_; 
wire _abc_44694_new_n1503_; 
wire _abc_44694_new_n1504_; 
wire _abc_44694_new_n1505_; 
wire _abc_44694_new_n1506_; 
wire _abc_44694_new_n1507_; 
wire _abc_44694_new_n1508_; 
wire _abc_44694_new_n1509_; 
wire _abc_44694_new_n1510_; 
wire _abc_44694_new_n1511_; 
wire _abc_44694_new_n1512_; 
wire _abc_44694_new_n1513_; 
wire _abc_44694_new_n1514_; 
wire _abc_44694_new_n1515_; 
wire _abc_44694_new_n1516_; 
wire _abc_44694_new_n1517_; 
wire _abc_44694_new_n1518_; 
wire _abc_44694_new_n1519_; 
wire _abc_44694_new_n1520_; 
wire _abc_44694_new_n1521_; 
wire _abc_44694_new_n1522_; 
wire _abc_44694_new_n1522__bF_buf0; 
wire _abc_44694_new_n1522__bF_buf1; 
wire _abc_44694_new_n1522__bF_buf2; 
wire _abc_44694_new_n1522__bF_buf3; 
wire _abc_44694_new_n1522__bF_buf4; 
wire _abc_44694_new_n1523_; 
wire _abc_44694_new_n1524_; 
wire _abc_44694_new_n1525_; 
wire _abc_44694_new_n1526_; 
wire _abc_44694_new_n1527_; 
wire _abc_44694_new_n1528_; 
wire _abc_44694_new_n1529_; 
wire _abc_44694_new_n1530_; 
wire _abc_44694_new_n1531_; 
wire _abc_44694_new_n1532_; 
wire _abc_44694_new_n1533_; 
wire _abc_44694_new_n1535_; 
wire _abc_44694_new_n1536_; 
wire _abc_44694_new_n1537_; 
wire _abc_44694_new_n1538_; 
wire _abc_44694_new_n1539_; 
wire _abc_44694_new_n1540_; 
wire _abc_44694_new_n1541_; 
wire _abc_44694_new_n1542_; 
wire _abc_44694_new_n1543_; 
wire _abc_44694_new_n1544_; 
wire _abc_44694_new_n1545_; 
wire _abc_44694_new_n1546_; 
wire _abc_44694_new_n1547_; 
wire _abc_44694_new_n1548_; 
wire _abc_44694_new_n1549_; 
wire _abc_44694_new_n1550_; 
wire _abc_44694_new_n1551_; 
wire _abc_44694_new_n1552_; 
wire _abc_44694_new_n1553_; 
wire _abc_44694_new_n1554_; 
wire _abc_44694_new_n1555_; 
wire _abc_44694_new_n1556_; 
wire _abc_44694_new_n1557_; 
wire _abc_44694_new_n1558_; 
wire _abc_44694_new_n1559_; 
wire _abc_44694_new_n1560_; 
wire _abc_44694_new_n1561_; 
wire _abc_44694_new_n1562_; 
wire _abc_44694_new_n1563_; 
wire _abc_44694_new_n1564_; 
wire _abc_44694_new_n1565_; 
wire _abc_44694_new_n1566_; 
wire _abc_44694_new_n1567_; 
wire _abc_44694_new_n1568_; 
wire _abc_44694_new_n1569_; 
wire _abc_44694_new_n1570_; 
wire _abc_44694_new_n1571_; 
wire _abc_44694_new_n1572_; 
wire _abc_44694_new_n1573_; 
wire _abc_44694_new_n1575_; 
wire _abc_44694_new_n1576_; 
wire _abc_44694_new_n1577_; 
wire _abc_44694_new_n1578_; 
wire _abc_44694_new_n1579_; 
wire _abc_44694_new_n1580_; 
wire _abc_44694_new_n1581_; 
wire _abc_44694_new_n1582_; 
wire _abc_44694_new_n1583_; 
wire _abc_44694_new_n1584_; 
wire _abc_44694_new_n1585_; 
wire _abc_44694_new_n1586_; 
wire _abc_44694_new_n1587_; 
wire _abc_44694_new_n1588_; 
wire _abc_44694_new_n1589_; 
wire _abc_44694_new_n1590_; 
wire _abc_44694_new_n1591_; 
wire _abc_44694_new_n1592_; 
wire _abc_44694_new_n1593_; 
wire _abc_44694_new_n1594_; 
wire _abc_44694_new_n1595_; 
wire _abc_44694_new_n1596_; 
wire _abc_44694_new_n1597_; 
wire _abc_44694_new_n1598_; 
wire _abc_44694_new_n1599_; 
wire _abc_44694_new_n1600_; 
wire _abc_44694_new_n1601_; 
wire _abc_44694_new_n1602_; 
wire _abc_44694_new_n1603_; 
wire _abc_44694_new_n1604_; 
wire _abc_44694_new_n1605_; 
wire _abc_44694_new_n1606_; 
wire _abc_44694_new_n1607_; 
wire _abc_44694_new_n1608_; 
wire _abc_44694_new_n1609_; 
wire _abc_44694_new_n1610_; 
wire _abc_44694_new_n1611_; 
wire _abc_44694_new_n1612_; 
wire _abc_44694_new_n1614_; 
wire _abc_44694_new_n1615_; 
wire _abc_44694_new_n1616_; 
wire _abc_44694_new_n1617_; 
wire _abc_44694_new_n1618_; 
wire _abc_44694_new_n1619_; 
wire _abc_44694_new_n1620_; 
wire _abc_44694_new_n1621_; 
wire _abc_44694_new_n1622_; 
wire _abc_44694_new_n1623_; 
wire _abc_44694_new_n1624_; 
wire _abc_44694_new_n1625_; 
wire _abc_44694_new_n1626_; 
wire _abc_44694_new_n1627_; 
wire _abc_44694_new_n1628_; 
wire _abc_44694_new_n1629_; 
wire _abc_44694_new_n1630_; 
wire _abc_44694_new_n1631_; 
wire _abc_44694_new_n1632_; 
wire _abc_44694_new_n1633_; 
wire _abc_44694_new_n1634_; 
wire _abc_44694_new_n1635_; 
wire _abc_44694_new_n1636_; 
wire _abc_44694_new_n1637_; 
wire _abc_44694_new_n1638_; 
wire _abc_44694_new_n1639_; 
wire _abc_44694_new_n1640_; 
wire _abc_44694_new_n1641_; 
wire _abc_44694_new_n1642_; 
wire _abc_44694_new_n1643_; 
wire _abc_44694_new_n1644_; 
wire _abc_44694_new_n1645_; 
wire _abc_44694_new_n1646_; 
wire _abc_44694_new_n1647_; 
wire _abc_44694_new_n1648_; 
wire _abc_44694_new_n1649_; 
wire _abc_44694_new_n1651_; 
wire _abc_44694_new_n1652_; 
wire _abc_44694_new_n1653_; 
wire _abc_44694_new_n1654_; 
wire _abc_44694_new_n1655_; 
wire _abc_44694_new_n1656_; 
wire _abc_44694_new_n1657_; 
wire _abc_44694_new_n1658_; 
wire _abc_44694_new_n1659_; 
wire _abc_44694_new_n1660_; 
wire _abc_44694_new_n1661_; 
wire _abc_44694_new_n1662_; 
wire _abc_44694_new_n1663_; 
wire _abc_44694_new_n1664_; 
wire _abc_44694_new_n1665_; 
wire _abc_44694_new_n1666_; 
wire _abc_44694_new_n1667_; 
wire _abc_44694_new_n1668_; 
wire _abc_44694_new_n1669_; 
wire _abc_44694_new_n1670_; 
wire _abc_44694_new_n1671_; 
wire _abc_44694_new_n1672_; 
wire _abc_44694_new_n1673_; 
wire _abc_44694_new_n1674_; 
wire _abc_44694_new_n1675_; 
wire _abc_44694_new_n1676_; 
wire _abc_44694_new_n1677_; 
wire _abc_44694_new_n1678_; 
wire _abc_44694_new_n1679_; 
wire _abc_44694_new_n1680_; 
wire _abc_44694_new_n1681_; 
wire _abc_44694_new_n1682_; 
wire _abc_44694_new_n1683_; 
wire _abc_44694_new_n1684_; 
wire _abc_44694_new_n1685_; 
wire _abc_44694_new_n1686_; 
wire _abc_44694_new_n1687_; 
wire _abc_44694_new_n1688_; 
wire _abc_44694_new_n1689_; 
wire _abc_44694_new_n1690_; 
wire _abc_44694_new_n1691_; 
wire _abc_44694_new_n1693_; 
wire _abc_44694_new_n1694_; 
wire _abc_44694_new_n1695_; 
wire _abc_44694_new_n1696_; 
wire _abc_44694_new_n1697_; 
wire _abc_44694_new_n1698_; 
wire _abc_44694_new_n1699_; 
wire _abc_44694_new_n1700_; 
wire _abc_44694_new_n1701_; 
wire _abc_44694_new_n1702_; 
wire _abc_44694_new_n1703_; 
wire _abc_44694_new_n1704_; 
wire _abc_44694_new_n1705_; 
wire _abc_44694_new_n1706_; 
wire _abc_44694_new_n1707_; 
wire _abc_44694_new_n1708_; 
wire _abc_44694_new_n1709_; 
wire _abc_44694_new_n1710_; 
wire _abc_44694_new_n1711_; 
wire _abc_44694_new_n1712_; 
wire _abc_44694_new_n1713_; 
wire _abc_44694_new_n1714_; 
wire _abc_44694_new_n1715_; 
wire _abc_44694_new_n1716_; 
wire _abc_44694_new_n1717_; 
wire _abc_44694_new_n1718_; 
wire _abc_44694_new_n1719_; 
wire _abc_44694_new_n1720_; 
wire _abc_44694_new_n1721_; 
wire _abc_44694_new_n1722_; 
wire _abc_44694_new_n1723_; 
wire _abc_44694_new_n1724_; 
wire _abc_44694_new_n1725_; 
wire _abc_44694_new_n1726_; 
wire _abc_44694_new_n1727_; 
wire _abc_44694_new_n1728_; 
wire _abc_44694_new_n1729_; 
wire _abc_44694_new_n1731_; 
wire _abc_44694_new_n1732_; 
wire _abc_44694_new_n1733_; 
wire _abc_44694_new_n1734_; 
wire _abc_44694_new_n1735_; 
wire _abc_44694_new_n1736_; 
wire _abc_44694_new_n1737_; 
wire _abc_44694_new_n1738_; 
wire _abc_44694_new_n1739_; 
wire _abc_44694_new_n1740_; 
wire _abc_44694_new_n1741_; 
wire _abc_44694_new_n1742_; 
wire _abc_44694_new_n1743_; 
wire _abc_44694_new_n1744_; 
wire _abc_44694_new_n1745_; 
wire _abc_44694_new_n1746_; 
wire _abc_44694_new_n1747_; 
wire _abc_44694_new_n1748_; 
wire _abc_44694_new_n1749_; 
wire _abc_44694_new_n1750_; 
wire _abc_44694_new_n1751_; 
wire _abc_44694_new_n1752_; 
wire _abc_44694_new_n1753_; 
wire _abc_44694_new_n1754_; 
wire _abc_44694_new_n1755_; 
wire _abc_44694_new_n1756_; 
wire _abc_44694_new_n1757_; 
wire _abc_44694_new_n1758_; 
wire _abc_44694_new_n1759_; 
wire _abc_44694_new_n1760_; 
wire _abc_44694_new_n1761_; 
wire _abc_44694_new_n1762_; 
wire _abc_44694_new_n1763_; 
wire _abc_44694_new_n1764_; 
wire _abc_44694_new_n1765_; 
wire _abc_44694_new_n1767_; 
wire _abc_44694_new_n1768_; 
wire _abc_44694_new_n1769_; 
wire _abc_44694_new_n1770_; 
wire _abc_44694_new_n1771_; 
wire _abc_44694_new_n1772_; 
wire _abc_44694_new_n1773_; 
wire _abc_44694_new_n1774_; 
wire _abc_44694_new_n1775_; 
wire _abc_44694_new_n1776_; 
wire _abc_44694_new_n1777_; 
wire _abc_44694_new_n1778_; 
wire _abc_44694_new_n1779_; 
wire _abc_44694_new_n1780_; 
wire _abc_44694_new_n1781_; 
wire _abc_44694_new_n1782_; 
wire _abc_44694_new_n1783_; 
wire _abc_44694_new_n1784_; 
wire _abc_44694_new_n1785_; 
wire _abc_44694_new_n1786_; 
wire _abc_44694_new_n1787_; 
wire _abc_44694_new_n1788_; 
wire _abc_44694_new_n1789_; 
wire _abc_44694_new_n1790_; 
wire _abc_44694_new_n1791_; 
wire _abc_44694_new_n1792_; 
wire _abc_44694_new_n1793_; 
wire _abc_44694_new_n1794_; 
wire _abc_44694_new_n1795_; 
wire _abc_44694_new_n1796_; 
wire _abc_44694_new_n1797_; 
wire _abc_44694_new_n1798_; 
wire _abc_44694_new_n1799_; 
wire _abc_44694_new_n1800_; 
wire _abc_44694_new_n1801_; 
wire _abc_44694_new_n1802_; 
wire _abc_44694_new_n1803_; 
wire _abc_44694_new_n1804_; 
wire _abc_44694_new_n1805_; 
wire _abc_44694_new_n1806_; 
wire _abc_44694_new_n1807_; 
wire _abc_44694_new_n1809_; 
wire _abc_44694_new_n1810_; 
wire _abc_44694_new_n1811_; 
wire _abc_44694_new_n1812_; 
wire _abc_44694_new_n1813_; 
wire _abc_44694_new_n1814_; 
wire _abc_44694_new_n1815_; 
wire _abc_44694_new_n1816_; 
wire _abc_44694_new_n1817_; 
wire _abc_44694_new_n1818_; 
wire _abc_44694_new_n1819_; 
wire _abc_44694_new_n1820_; 
wire _abc_44694_new_n1821_; 
wire _abc_44694_new_n1822_; 
wire _abc_44694_new_n1823_; 
wire _abc_44694_new_n1824_; 
wire _abc_44694_new_n1825_; 
wire _abc_44694_new_n1826_; 
wire _abc_44694_new_n1827_; 
wire _abc_44694_new_n1828_; 
wire _abc_44694_new_n1829_; 
wire _abc_44694_new_n1830_; 
wire _abc_44694_new_n1831_; 
wire _abc_44694_new_n1832_; 
wire _abc_44694_new_n1833_; 
wire _abc_44694_new_n1834_; 
wire _abc_44694_new_n1835_; 
wire _abc_44694_new_n1836_; 
wire _abc_44694_new_n1837_; 
wire _abc_44694_new_n1838_; 
wire _abc_44694_new_n1839_; 
wire _abc_44694_new_n1840_; 
wire _abc_44694_new_n1841_; 
wire _abc_44694_new_n1842_; 
wire _abc_44694_new_n1843_; 
wire _abc_44694_new_n1844_; 
wire _abc_44694_new_n1845_; 
wire _abc_44694_new_n1846_; 
wire _abc_44694_new_n1848_; 
wire _abc_44694_new_n1849_; 
wire _abc_44694_new_n1850_; 
wire _abc_44694_new_n1851_; 
wire _abc_44694_new_n1852_; 
wire _abc_44694_new_n1853_; 
wire _abc_44694_new_n1854_; 
wire _abc_44694_new_n1855_; 
wire _abc_44694_new_n1856_; 
wire _abc_44694_new_n1857_; 
wire _abc_44694_new_n1858_; 
wire _abc_44694_new_n1859_; 
wire _abc_44694_new_n1860_; 
wire _abc_44694_new_n1861_; 
wire _abc_44694_new_n1862_; 
wire _abc_44694_new_n1863_; 
wire _abc_44694_new_n1864_; 
wire _abc_44694_new_n1865_; 
wire _abc_44694_new_n1866_; 
wire _abc_44694_new_n1867_; 
wire _abc_44694_new_n1868_; 
wire _abc_44694_new_n1869_; 
wire _abc_44694_new_n1870_; 
wire _abc_44694_new_n1871_; 
wire _abc_44694_new_n1872_; 
wire _abc_44694_new_n1873_; 
wire _abc_44694_new_n1874_; 
wire _abc_44694_new_n1875_; 
wire _abc_44694_new_n1876_; 
wire _abc_44694_new_n1877_; 
wire _abc_44694_new_n1878_; 
wire _abc_44694_new_n1879_; 
wire _abc_44694_new_n1880_; 
wire _abc_44694_new_n1881_; 
wire _abc_44694_new_n1882_; 
wire _abc_44694_new_n1883_; 
wire _abc_44694_new_n1885_; 
wire _abc_44694_new_n1886_; 
wire _abc_44694_new_n1887_; 
wire _abc_44694_new_n1888_; 
wire _abc_44694_new_n1889_; 
wire _abc_44694_new_n1890_; 
wire _abc_44694_new_n1891_; 
wire _abc_44694_new_n1892_; 
wire _abc_44694_new_n1893_; 
wire _abc_44694_new_n1894_; 
wire _abc_44694_new_n1895_; 
wire _abc_44694_new_n1896_; 
wire _abc_44694_new_n1897_; 
wire _abc_44694_new_n1898_; 
wire _abc_44694_new_n1899_; 
wire _abc_44694_new_n1900_; 
wire _abc_44694_new_n1901_; 
wire _abc_44694_new_n1902_; 
wire _abc_44694_new_n1903_; 
wire _abc_44694_new_n1904_; 
wire _abc_44694_new_n1905_; 
wire _abc_44694_new_n1906_; 
wire _abc_44694_new_n1907_; 
wire _abc_44694_new_n1908_; 
wire _abc_44694_new_n1909_; 
wire _abc_44694_new_n1910_; 
wire _abc_44694_new_n1911_; 
wire _abc_44694_new_n1912_; 
wire _abc_44694_new_n1913_; 
wire _abc_44694_new_n1914_; 
wire _abc_44694_new_n1915_; 
wire _abc_44694_new_n1916_; 
wire _abc_44694_new_n1917_; 
wire _abc_44694_new_n1918_; 
wire _abc_44694_new_n1919_; 
wire _abc_44694_new_n1921_; 
wire _abc_44694_new_n1922_; 
wire _abc_44694_new_n1923_; 
wire _abc_44694_new_n1924_; 
wire _abc_44694_new_n1925_; 
wire _abc_44694_new_n1926_; 
wire _abc_44694_new_n1927_; 
wire _abc_44694_new_n1928_; 
wire _abc_44694_new_n1929_; 
wire _abc_44694_new_n1930_; 
wire _abc_44694_new_n1931_; 
wire _abc_44694_new_n1932_; 
wire _abc_44694_new_n1933_; 
wire _abc_44694_new_n1934_; 
wire _abc_44694_new_n1935_; 
wire _abc_44694_new_n1936_; 
wire _abc_44694_new_n1937_; 
wire _abc_44694_new_n1938_; 
wire _abc_44694_new_n1939_; 
wire _abc_44694_new_n1940_; 
wire _abc_44694_new_n1941_; 
wire _abc_44694_new_n1942_; 
wire _abc_44694_new_n1943_; 
wire _abc_44694_new_n1944_; 
wire _abc_44694_new_n1945_; 
wire _abc_44694_new_n1946_; 
wire _abc_44694_new_n1947_; 
wire _abc_44694_new_n1948_; 
wire _abc_44694_new_n1949_; 
wire _abc_44694_new_n1950_; 
wire _abc_44694_new_n1951_; 
wire _abc_44694_new_n1952_; 
wire _abc_44694_new_n1953_; 
wire _abc_44694_new_n1954_; 
wire _abc_44694_new_n1955_; 
wire _abc_44694_new_n1956_; 
wire _abc_44694_new_n1957_; 
wire _abc_44694_new_n1958_; 
wire _abc_44694_new_n1959_; 
wire _abc_44694_new_n1960_; 
wire _abc_44694_new_n1961_; 
wire _abc_44694_new_n1962_; 
wire _abc_44694_new_n1963_; 
wire _abc_44694_new_n1964_; 
wire _abc_44694_new_n1965_; 
wire _abc_44694_new_n1967_; 
wire _abc_44694_new_n1968_; 
wire _abc_44694_new_n1969_; 
wire _abc_44694_new_n1970_; 
wire _abc_44694_new_n1971_; 
wire _abc_44694_new_n1972_; 
wire _abc_44694_new_n1973_; 
wire _abc_44694_new_n1974_; 
wire _abc_44694_new_n1975_; 
wire _abc_44694_new_n1976_; 
wire _abc_44694_new_n1977_; 
wire _abc_44694_new_n1978_; 
wire _abc_44694_new_n1979_; 
wire _abc_44694_new_n1980_; 
wire _abc_44694_new_n1981_; 
wire _abc_44694_new_n1982_; 
wire _abc_44694_new_n1983_; 
wire _abc_44694_new_n1984_; 
wire _abc_44694_new_n1985_; 
wire _abc_44694_new_n1986_; 
wire _abc_44694_new_n1987_; 
wire _abc_44694_new_n1988_; 
wire _abc_44694_new_n1989_; 
wire _abc_44694_new_n1990_; 
wire _abc_44694_new_n1991_; 
wire _abc_44694_new_n1992_; 
wire _abc_44694_new_n1993_; 
wire _abc_44694_new_n1994_; 
wire _abc_44694_new_n1995_; 
wire _abc_44694_new_n1996_; 
wire _abc_44694_new_n1997_; 
wire _abc_44694_new_n1998_; 
wire _abc_44694_new_n1999_; 
wire _abc_44694_new_n2000_; 
wire _abc_44694_new_n2001_; 
wire _abc_44694_new_n2003_; 
wire _abc_44694_new_n2004_; 
wire _abc_44694_new_n2005_; 
wire _abc_44694_new_n2006_; 
wire _abc_44694_new_n2007_; 
wire _abc_44694_new_n2008_; 
wire _abc_44694_new_n2009_; 
wire _abc_44694_new_n2010_; 
wire _abc_44694_new_n2011_; 
wire _abc_44694_new_n2012_; 
wire _abc_44694_new_n2013_; 
wire _abc_44694_new_n2014_; 
wire _abc_44694_new_n2015_; 
wire _abc_44694_new_n2016_; 
wire _abc_44694_new_n2017_; 
wire _abc_44694_new_n2018_; 
wire _abc_44694_new_n2019_; 
wire _abc_44694_new_n2020_; 
wire _abc_44694_new_n2021_; 
wire _abc_44694_new_n2022_; 
wire _abc_44694_new_n2023_; 
wire _abc_44694_new_n2024_; 
wire _abc_44694_new_n2025_; 
wire _abc_44694_new_n2026_; 
wire _abc_44694_new_n2027_; 
wire _abc_44694_new_n2028_; 
wire _abc_44694_new_n2029_; 
wire _abc_44694_new_n2030_; 
wire _abc_44694_new_n2031_; 
wire _abc_44694_new_n2032_; 
wire _abc_44694_new_n2033_; 
wire _abc_44694_new_n2034_; 
wire _abc_44694_new_n2035_; 
wire _abc_44694_new_n2036_; 
wire _abc_44694_new_n2037_; 
wire _abc_44694_new_n2039_; 
wire _abc_44694_new_n2040_; 
wire _abc_44694_new_n2041_; 
wire _abc_44694_new_n2042_; 
wire _abc_44694_new_n2043_; 
wire _abc_44694_new_n2044_; 
wire _abc_44694_new_n2045_; 
wire _abc_44694_new_n2046_; 
wire _abc_44694_new_n2047_; 
wire _abc_44694_new_n2048_; 
wire _abc_44694_new_n2049_; 
wire _abc_44694_new_n2050_; 
wire _abc_44694_new_n2051_; 
wire _abc_44694_new_n2052_; 
wire _abc_44694_new_n2053_; 
wire _abc_44694_new_n2054_; 
wire _abc_44694_new_n2055_; 
wire _abc_44694_new_n2056_; 
wire _abc_44694_new_n2057_; 
wire _abc_44694_new_n2058_; 
wire _abc_44694_new_n2059_; 
wire _abc_44694_new_n2060_; 
wire _abc_44694_new_n2061_; 
wire _abc_44694_new_n2062_; 
wire _abc_44694_new_n2063_; 
wire _abc_44694_new_n2064_; 
wire _abc_44694_new_n2065_; 
wire _abc_44694_new_n2066_; 
wire _abc_44694_new_n2067_; 
wire _abc_44694_new_n2068_; 
wire _abc_44694_new_n2069_; 
wire _abc_44694_new_n2070_; 
wire _abc_44694_new_n2071_; 
wire _abc_44694_new_n2072_; 
wire _abc_44694_new_n2073_; 
wire _abc_44694_new_n2075_; 
wire _abc_44694_new_n2076_; 
wire _abc_44694_new_n2077_; 
wire _abc_44694_new_n2078_; 
wire _abc_44694_new_n2079_; 
wire _abc_44694_new_n2080_; 
wire _abc_44694_new_n2081_; 
wire _abc_44694_new_n2082_; 
wire _abc_44694_new_n2083_; 
wire _abc_44694_new_n2084_; 
wire _abc_44694_new_n2085_; 
wire _abc_44694_new_n2086_; 
wire _abc_44694_new_n2087_; 
wire _abc_44694_new_n2088_; 
wire _abc_44694_new_n2089_; 
wire _abc_44694_new_n2090_; 
wire _abc_44694_new_n2091_; 
wire _abc_44694_new_n2092_; 
wire _abc_44694_new_n2093_; 
wire _abc_44694_new_n2094_; 
wire _abc_44694_new_n2095_; 
wire _abc_44694_new_n2096_; 
wire _abc_44694_new_n2097_; 
wire _abc_44694_new_n2098_; 
wire _abc_44694_new_n2099_; 
wire _abc_44694_new_n2100_; 
wire _abc_44694_new_n2101_; 
wire _abc_44694_new_n2102_; 
wire _abc_44694_new_n2103_; 
wire _abc_44694_new_n2104_; 
wire _abc_44694_new_n2105_; 
wire _abc_44694_new_n2106_; 
wire _abc_44694_new_n2107_; 
wire _abc_44694_new_n2108_; 
wire _abc_44694_new_n2109_; 
wire _abc_44694_new_n2110_; 
wire _abc_44694_new_n2111_; 
wire _abc_44694_new_n2112_; 
wire _abc_44694_new_n2113_; 
wire _abc_44694_new_n2114_; 
wire _abc_44694_new_n2115_; 
wire _abc_44694_new_n2116_; 
wire _abc_44694_new_n2117_; 
wire _abc_44694_new_n2118_; 
wire _abc_44694_new_n2119_; 
wire _abc_44694_new_n2120_; 
wire _abc_44694_new_n2121_; 
wire _abc_44694_new_n2122_; 
wire _abc_44694_new_n2124_; 
wire _abc_44694_new_n2125_; 
wire _abc_44694_new_n2126_; 
wire _abc_44694_new_n2127_; 
wire _abc_44694_new_n2128_; 
wire _abc_44694_new_n2129_; 
wire _abc_44694_new_n2130_; 
wire _abc_44694_new_n2131_; 
wire _abc_44694_new_n2132_; 
wire _abc_44694_new_n2133_; 
wire _abc_44694_new_n2134_; 
wire _abc_44694_new_n2135_; 
wire _abc_44694_new_n2136_; 
wire _abc_44694_new_n2137_; 
wire _abc_44694_new_n2138_; 
wire _abc_44694_new_n2139_; 
wire _abc_44694_new_n2140_; 
wire _abc_44694_new_n2141_; 
wire _abc_44694_new_n2142_; 
wire _abc_44694_new_n2143_; 
wire _abc_44694_new_n2144_; 
wire _abc_44694_new_n2145_; 
wire _abc_44694_new_n2146_; 
wire _abc_44694_new_n2147_; 
wire _abc_44694_new_n2148_; 
wire _abc_44694_new_n2149_; 
wire _abc_44694_new_n2150_; 
wire _abc_44694_new_n2151_; 
wire _abc_44694_new_n2152_; 
wire _abc_44694_new_n2153_; 
wire _abc_44694_new_n2154_; 
wire _abc_44694_new_n2155_; 
wire _abc_44694_new_n2156_; 
wire _abc_44694_new_n2157_; 
wire _abc_44694_new_n2158_; 
wire _abc_44694_new_n2159_; 
wire _abc_44694_new_n2160_; 
wire _abc_44694_new_n2161_; 
wire _abc_44694_new_n2163_; 
wire _abc_44694_new_n2164_; 
wire _abc_44694_new_n2165_; 
wire _abc_44694_new_n2166_; 
wire _abc_44694_new_n2167_; 
wire _abc_44694_new_n2168_; 
wire _abc_44694_new_n2169_; 
wire _abc_44694_new_n2170_; 
wire _abc_44694_new_n2171_; 
wire _abc_44694_new_n2172_; 
wire _abc_44694_new_n2173_; 
wire _abc_44694_new_n2174_; 
wire _abc_44694_new_n2175_; 
wire _abc_44694_new_n2176_; 
wire _abc_44694_new_n2177_; 
wire _abc_44694_new_n2178_; 
wire _abc_44694_new_n2179_; 
wire _abc_44694_new_n2180_; 
wire _abc_44694_new_n2181_; 
wire _abc_44694_new_n2182_; 
wire _abc_44694_new_n2183_; 
wire _abc_44694_new_n2184_; 
wire _abc_44694_new_n2185_; 
wire _abc_44694_new_n2186_; 
wire _abc_44694_new_n2187_; 
wire _abc_44694_new_n2188_; 
wire _abc_44694_new_n2189_; 
wire _abc_44694_new_n2190_; 
wire _abc_44694_new_n2191_; 
wire _abc_44694_new_n2192_; 
wire _abc_44694_new_n2193_; 
wire _abc_44694_new_n2194_; 
wire _abc_44694_new_n2195_; 
wire _abc_44694_new_n2196_; 
wire _abc_44694_new_n2197_; 
wire _abc_44694_new_n2198_; 
wire _abc_44694_new_n2200_; 
wire _abc_44694_new_n2201_; 
wire _abc_44694_new_n2202_; 
wire _abc_44694_new_n2203_; 
wire _abc_44694_new_n2204_; 
wire _abc_44694_new_n2205_; 
wire _abc_44694_new_n2206_; 
wire _abc_44694_new_n2207_; 
wire _abc_44694_new_n2208_; 
wire _abc_44694_new_n2209_; 
wire _abc_44694_new_n2210_; 
wire _abc_44694_new_n2211_; 
wire _abc_44694_new_n2212_; 
wire _abc_44694_new_n2213_; 
wire _abc_44694_new_n2214_; 
wire _abc_44694_new_n2215_; 
wire _abc_44694_new_n2216_; 
wire _abc_44694_new_n2217_; 
wire _abc_44694_new_n2218_; 
wire _abc_44694_new_n2219_; 
wire _abc_44694_new_n2220_; 
wire _abc_44694_new_n2221_; 
wire _abc_44694_new_n2222_; 
wire _abc_44694_new_n2223_; 
wire _abc_44694_new_n2224_; 
wire _abc_44694_new_n2225_; 
wire _abc_44694_new_n2226_; 
wire _abc_44694_new_n2227_; 
wire _abc_44694_new_n2228_; 
wire _abc_44694_new_n2229_; 
wire _abc_44694_new_n2230_; 
wire _abc_44694_new_n2231_; 
wire _abc_44694_new_n2232_; 
wire _abc_44694_new_n2233_; 
wire _abc_44694_new_n2234_; 
wire _abc_44694_new_n2236_; 
wire _abc_44694_new_n2237_; 
wire _abc_44694_new_n2238_; 
wire _abc_44694_new_n2239_; 
wire _abc_44694_new_n2240_; 
wire _abc_44694_new_n2241_; 
wire _abc_44694_new_n2242_; 
wire _abc_44694_new_n2243_; 
wire _abc_44694_new_n2244_; 
wire _abc_44694_new_n2245_; 
wire _abc_44694_new_n2246_; 
wire _abc_44694_new_n2247_; 
wire _abc_44694_new_n2248_; 
wire _abc_44694_new_n2249_; 
wire _abc_44694_new_n2250_; 
wire _abc_44694_new_n2251_; 
wire _abc_44694_new_n2252_; 
wire _abc_44694_new_n2253_; 
wire _abc_44694_new_n2254_; 
wire _abc_44694_new_n2255_; 
wire _abc_44694_new_n2256_; 
wire _abc_44694_new_n2257_; 
wire _abc_44694_new_n2258_; 
wire _abc_44694_new_n2259_; 
wire _abc_44694_new_n2260_; 
wire _abc_44694_new_n2261_; 
wire _abc_44694_new_n2262_; 
wire _abc_44694_new_n2263_; 
wire _abc_44694_new_n2264_; 
wire _abc_44694_new_n2265_; 
wire _abc_44694_new_n2266_; 
wire _abc_44694_new_n2267_; 
wire _abc_44694_new_n2268_; 
wire _abc_44694_new_n2269_; 
wire _abc_44694_new_n2270_; 
wire _abc_44694_new_n2271_; 
wire _abc_44694_new_n2272_; 
wire _abc_44694_new_n2273_; 
wire _abc_44694_new_n2274_; 
wire _abc_44694_new_n2275_; 
wire _abc_44694_new_n2276_; 
wire _abc_44694_new_n2277_; 
wire _abc_44694_new_n2278_; 
wire _abc_44694_new_n2279_; 
wire _abc_44694_new_n2280_; 
wire _abc_44694_new_n2282_; 
wire _abc_44694_new_n2283_; 
wire _abc_44694_new_n2284_; 
wire _abc_44694_new_n2285_; 
wire _abc_44694_new_n2286_; 
wire _abc_44694_new_n2287_; 
wire _abc_44694_new_n2288_; 
wire _abc_44694_new_n2289_; 
wire _abc_44694_new_n2290_; 
wire _abc_44694_new_n2291_; 
wire _abc_44694_new_n2292_; 
wire _abc_44694_new_n2293_; 
wire _abc_44694_new_n2294_; 
wire _abc_44694_new_n2295_; 
wire _abc_44694_new_n2296_; 
wire _abc_44694_new_n2297_; 
wire _abc_44694_new_n2298_; 
wire _abc_44694_new_n2299_; 
wire _abc_44694_new_n2300_; 
wire _abc_44694_new_n2301_; 
wire _abc_44694_new_n2302_; 
wire _abc_44694_new_n2303_; 
wire _abc_44694_new_n2304_; 
wire _abc_44694_new_n2305_; 
wire _abc_44694_new_n2306_; 
wire _abc_44694_new_n2307_; 
wire _abc_44694_new_n2308_; 
wire _abc_44694_new_n2309_; 
wire _abc_44694_new_n2310_; 
wire _abc_44694_new_n2311_; 
wire _abc_44694_new_n2312_; 
wire _abc_44694_new_n2313_; 
wire _abc_44694_new_n2314_; 
wire _abc_44694_new_n2315_; 
wire _abc_44694_new_n2316_; 
wire _abc_44694_new_n2317_; 
wire _abc_44694_new_n2318_; 
wire _abc_44694_new_n2319_; 
wire _abc_44694_new_n2321_; 
wire _abc_44694_new_n2322_; 
wire _abc_44694_new_n2323_; 
wire _abc_44694_new_n2324_; 
wire _abc_44694_new_n2325_; 
wire _abc_44694_new_n2326_; 
wire _abc_44694_new_n2327_; 
wire _abc_44694_new_n2328_; 
wire _abc_44694_new_n2329_; 
wire _abc_44694_new_n2330_; 
wire _abc_44694_new_n2331_; 
wire _abc_44694_new_n2332_; 
wire _abc_44694_new_n2333_; 
wire _abc_44694_new_n2334_; 
wire _abc_44694_new_n2335_; 
wire _abc_44694_new_n2336_; 
wire _abc_44694_new_n2337_; 
wire _abc_44694_new_n2338_; 
wire _abc_44694_new_n2339_; 
wire _abc_44694_new_n2340_; 
wire _abc_44694_new_n2341_; 
wire _abc_44694_new_n2342_; 
wire _abc_44694_new_n2343_; 
wire _abc_44694_new_n2344_; 
wire _abc_44694_new_n2345_; 
wire _abc_44694_new_n2346_; 
wire _abc_44694_new_n2347_; 
wire _abc_44694_new_n2348_; 
wire _abc_44694_new_n2349_; 
wire _abc_44694_new_n2350_; 
wire _abc_44694_new_n2351_; 
wire _abc_44694_new_n2352_; 
wire _abc_44694_new_n2353_; 
wire _abc_44694_new_n2354_; 
wire _abc_44694_new_n2355_; 
wire _abc_44694_new_n2356_; 
wire _abc_44694_new_n2358_; 
wire _abc_44694_new_n2359_; 
wire _abc_44694_new_n2360_; 
wire _abc_44694_new_n2361_; 
wire _abc_44694_new_n2362_; 
wire _abc_44694_new_n2363_; 
wire _abc_44694_new_n2364_; 
wire _abc_44694_new_n2365_; 
wire _abc_44694_new_n2366_; 
wire _abc_44694_new_n2367_; 
wire _abc_44694_new_n2368_; 
wire _abc_44694_new_n2369_; 
wire _abc_44694_new_n2370_; 
wire _abc_44694_new_n2371_; 
wire _abc_44694_new_n2372_; 
wire _abc_44694_new_n2373_; 
wire _abc_44694_new_n2374_; 
wire _abc_44694_new_n2375_; 
wire _abc_44694_new_n2376_; 
wire _abc_44694_new_n2377_; 
wire _abc_44694_new_n2378_; 
wire _abc_44694_new_n2379_; 
wire _abc_44694_new_n2380_; 
wire _abc_44694_new_n2381_; 
wire _abc_44694_new_n2382_; 
wire _abc_44694_new_n2383_; 
wire _abc_44694_new_n2384_; 
wire _abc_44694_new_n2385_; 
wire _abc_44694_new_n2386_; 
wire _abc_44694_new_n2387_; 
wire _abc_44694_new_n2388_; 
wire _abc_44694_new_n2389_; 
wire _abc_44694_new_n2390_; 
wire _abc_44694_new_n2391_; 
wire _abc_44694_new_n2392_; 
wire _abc_44694_new_n2393_; 
wire _abc_44694_new_n2394_; 
wire _abc_44694_new_n2395_; 
wire _abc_44694_new_n2397_; 
wire _abc_44694_new_n2398_; 
wire _abc_44694_new_n2399_; 
wire _abc_44694_new_n2400_; 
wire _abc_44694_new_n2401_; 
wire _abc_44694_new_n2402_; 
wire _abc_44694_new_n2403_; 
wire _abc_44694_new_n2404_; 
wire _abc_44694_new_n2405_; 
wire _abc_44694_new_n2406_; 
wire _abc_44694_new_n2407_; 
wire _abc_44694_new_n2408_; 
wire _abc_44694_new_n2409_; 
wire _abc_44694_new_n2410_; 
wire _abc_44694_new_n2411_; 
wire _abc_44694_new_n2412_; 
wire _abc_44694_new_n2413_; 
wire _abc_44694_new_n2414_; 
wire _abc_44694_new_n2415_; 
wire _abc_44694_new_n2416_; 
wire _abc_44694_new_n2417_; 
wire _abc_44694_new_n2418_; 
wire _abc_44694_new_n2419_; 
wire _abc_44694_new_n2420_; 
wire _abc_44694_new_n2421_; 
wire _abc_44694_new_n2422_; 
wire _abc_44694_new_n2423_; 
wire _abc_44694_new_n2424_; 
wire _abc_44694_new_n2425_; 
wire _abc_44694_new_n2426_; 
wire _abc_44694_new_n2427_; 
wire _abc_44694_new_n2428_; 
wire _abc_44694_new_n2429_; 
wire _abc_44694_new_n2430_; 
wire _abc_44694_new_n2431_; 
wire _abc_44694_new_n2432_; 
wire _abc_44694_new_n2434_; 
wire _abc_44694_new_n2435_; 
wire _abc_44694_new_n2436_; 
wire _abc_44694_new_n2437_; 
wire _abc_44694_new_n2438_; 
wire _abc_44694_new_n2439_; 
wire _abc_44694_new_n2440_; 
wire _abc_44694_new_n2441_; 
wire _abc_44694_new_n2442_; 
wire _abc_44694_new_n2443_; 
wire _abc_44694_new_n2444_; 
wire _abc_44694_new_n2445_; 
wire _abc_44694_new_n2446_; 
wire _abc_44694_new_n2447_; 
wire _abc_44694_new_n2448_; 
wire _abc_44694_new_n2449_; 
wire _abc_44694_new_n2450_; 
wire _abc_44694_new_n2451_; 
wire _abc_44694_new_n2452_; 
wire _abc_44694_new_n2453_; 
wire _abc_44694_new_n2454_; 
wire _abc_44694_new_n2455_; 
wire _abc_44694_new_n2456_; 
wire _abc_44694_new_n2457_; 
wire _abc_44694_new_n2458_; 
wire _abc_44694_new_n2459_; 
wire _abc_44694_new_n2460_; 
wire _abc_44694_new_n2461_; 
wire _abc_44694_new_n2462_; 
wire _abc_44694_new_n2463_; 
wire _abc_44694_new_n2464_; 
wire _abc_44694_new_n2465_; 
wire _abc_44694_new_n2466_; 
wire _abc_44694_new_n2467_; 
wire _abc_44694_new_n2468_; 
wire _abc_44694_new_n2470_; 
wire _abc_44694_new_n2471_; 
wire _abc_44694_new_n2472_; 
wire _abc_44694_new_n2473_; 
wire _abc_44694_new_n2474_; 
wire _abc_44694_new_n2475_; 
wire _abc_44694_new_n2476_; 
wire _abc_44694_new_n2477_; 
wire _abc_44694_new_n2478_; 
wire _abc_44694_new_n2479_; 
wire _abc_44694_new_n2480_; 
wire _abc_44694_new_n2481_; 
wire _abc_44694_new_n2482_; 
wire _abc_44694_new_n2483_; 
wire _abc_44694_new_n2484_; 
wire _abc_44694_new_n2485_; 
wire _abc_44694_new_n2486_; 
wire _abc_44694_new_n2487_; 
wire _abc_44694_new_n2488_; 
wire _abc_44694_new_n2489_; 
wire _abc_44694_new_n2490_; 
wire _abc_44694_new_n2491_; 
wire _abc_44694_new_n2492_; 
wire _abc_44694_new_n2493_; 
wire _abc_44694_new_n2494_; 
wire _abc_44694_new_n2495_; 
wire _abc_44694_new_n2496_; 
wire _abc_44694_new_n2497_; 
wire _abc_44694_new_n2498_; 
wire _abc_44694_new_n2499_; 
wire _abc_44694_new_n2500_; 
wire _abc_44694_new_n2501_; 
wire _abc_44694_new_n2502_; 
wire _abc_44694_new_n2503_; 
wire _abc_44694_new_n2504_; 
wire _abc_44694_new_n2505_; 
wire _abc_44694_new_n2506_; 
wire _abc_44694_new_n2507_; 
wire _abc_44694_new_n2508_; 
wire _abc_44694_new_n2509_; 
wire _abc_44694_new_n2511_; 
wire _abc_44694_new_n2512_; 
wire _abc_44694_new_n2513_; 
wire _abc_44694_new_n2514_; 
wire _abc_44694_new_n2515_; 
wire _abc_44694_new_n2516_; 
wire _abc_44694_new_n2517_; 
wire _abc_44694_new_n2518_; 
wire _abc_44694_new_n2519_; 
wire _abc_44694_new_n2520_; 
wire _abc_44694_new_n2521_; 
wire _abc_44694_new_n2522_; 
wire _abc_44694_new_n2523_; 
wire _abc_44694_new_n2524_; 
wire _abc_44694_new_n2525_; 
wire _abc_44694_new_n2526_; 
wire _abc_44694_new_n2527_; 
wire _abc_44694_new_n2528_; 
wire _abc_44694_new_n2529_; 
wire _abc_44694_new_n2530_; 
wire _abc_44694_new_n2531_; 
wire _abc_44694_new_n2532_; 
wire _abc_44694_new_n2533_; 
wire _abc_44694_new_n2534_; 
wire _abc_44694_new_n2535_; 
wire _abc_44694_new_n2536_; 
wire _abc_44694_new_n2537_; 
wire _abc_44694_new_n2538_; 
wire _abc_44694_new_n2539_; 
wire _abc_44694_new_n2540_; 
wire _abc_44694_new_n2541_; 
wire _abc_44694_new_n2542_; 
wire _abc_44694_new_n2543_; 
wire _abc_44694_new_n2544_; 
wire _abc_44694_new_n2546_; 
wire _abc_44694_new_n2546__bF_buf0; 
wire _abc_44694_new_n2546__bF_buf1; 
wire _abc_44694_new_n2546__bF_buf2; 
wire _abc_44694_new_n2546__bF_buf3; 
wire _abc_44694_new_n2546__bF_buf4; 
wire _abc_44694_new_n2547_; 
wire _abc_44694_new_n2548_; 
wire _abc_44694_new_n2549_; 
wire _abc_44694_new_n2550_; 
wire _abc_44694_new_n2552_; 
wire _abc_44694_new_n2553_; 
wire _abc_44694_new_n2554_; 
wire _abc_44694_new_n2555_; 
wire _abc_44694_new_n2557_; 
wire _abc_44694_new_n2558_; 
wire _abc_44694_new_n2559_; 
wire _abc_44694_new_n2560_; 
wire _abc_44694_new_n2562_; 
wire _abc_44694_new_n2563_; 
wire _abc_44694_new_n2564_; 
wire _abc_44694_new_n2565_; 
wire _abc_44694_new_n2567_; 
wire _abc_44694_new_n2568_; 
wire _abc_44694_new_n2569_; 
wire _abc_44694_new_n2570_; 
wire _abc_44694_new_n2572_; 
wire _abc_44694_new_n2573_; 
wire _abc_44694_new_n2574_; 
wire _abc_44694_new_n2575_; 
wire _abc_44694_new_n2577_; 
wire _abc_44694_new_n2578_; 
wire _abc_44694_new_n2579_; 
wire _abc_44694_new_n2580_; 
wire _abc_44694_new_n2582_; 
wire _abc_44694_new_n2583_; 
wire _abc_44694_new_n2584_; 
wire _abc_44694_new_n2585_; 
wire _abc_44694_new_n2587_; 
wire _abc_44694_new_n2588_; 
wire _abc_44694_new_n2589_; 
wire _abc_44694_new_n2590_; 
wire _abc_44694_new_n2592_; 
wire _abc_44694_new_n2593_; 
wire _abc_44694_new_n2594_; 
wire _abc_44694_new_n2595_; 
wire _abc_44694_new_n2596_; 
wire _abc_44694_new_n2597_; 
wire _abc_44694_new_n2598_; 
wire _abc_44694_new_n2600_; 
wire _abc_44694_new_n2601_; 
wire _abc_44694_new_n2602_; 
wire _abc_44694_new_n2603_; 
wire _abc_44694_new_n2604_; 
wire _abc_44694_new_n2605_; 
wire _abc_44694_new_n2606_; 
wire _abc_44694_new_n2608_; 
wire _abc_44694_new_n2609_; 
wire _abc_44694_new_n2610_; 
wire _abc_44694_new_n2611_; 
wire _abc_44694_new_n2612_; 
wire _abc_44694_new_n2613_; 
wire _abc_44694_new_n2614_; 
wire _abc_44694_new_n2616_; 
wire _abc_44694_new_n2617_; 
wire _abc_44694_new_n2618_; 
wire _abc_44694_new_n2619_; 
wire _abc_44694_new_n2621_; 
wire _abc_44694_new_n2622_; 
wire _abc_44694_new_n2623_; 
wire _abc_44694_new_n2624_; 
wire _abc_44694_new_n2626_; 
wire _abc_44694_new_n2627_; 
wire _abc_44694_new_n2628_; 
wire _abc_44694_new_n2629_; 
wire _abc_44694_new_n2631_; 
wire _abc_44694_new_n2632_; 
wire _abc_44694_new_n2633_; 
wire _abc_44694_new_n2634_; 
wire _abc_44694_new_n2636_; 
wire _abc_44694_new_n2637_; 
wire _abc_44694_new_n2638_; 
wire _abc_44694_new_n2639_; 
wire _abc_44694_new_n2641_; 
wire _abc_44694_new_n2642_; 
wire _abc_44694_new_n2643_; 
wire _abc_44694_new_n2644_; 
wire _abc_44694_new_n2646_; 
wire _abc_44694_new_n2647_; 
wire _abc_44694_new_n2648_; 
wire _abc_44694_new_n2649_; 
wire _abc_44694_new_n2651_; 
wire _abc_44694_new_n2652_; 
wire _abc_44694_new_n2653_; 
wire _abc_44694_new_n2654_; 
wire _abc_44694_new_n2656_; 
wire _abc_44694_new_n2657_; 
wire _abc_44694_new_n2658_; 
wire _abc_44694_new_n2659_; 
wire _abc_44694_new_n2661_; 
wire _abc_44694_new_n2662_; 
wire _abc_44694_new_n2663_; 
wire _abc_44694_new_n2664_; 
wire _abc_44694_new_n2666_; 
wire _abc_44694_new_n2667_; 
wire _abc_44694_new_n2668_; 
wire _abc_44694_new_n2669_; 
wire _abc_44694_new_n2671_; 
wire _abc_44694_new_n2672_; 
wire _abc_44694_new_n2673_; 
wire _abc_44694_new_n2674_; 
wire _abc_44694_new_n2676_; 
wire _abc_44694_new_n2677_; 
wire _abc_44694_new_n2678_; 
wire _abc_44694_new_n2679_; 
wire _abc_44694_new_n2681_; 
wire _abc_44694_new_n2682_; 
wire _abc_44694_new_n2683_; 
wire _abc_44694_new_n2684_; 
wire _abc_44694_new_n2686_; 
wire _abc_44694_new_n2687_; 
wire _abc_44694_new_n2688_; 
wire _abc_44694_new_n2689_; 
wire _abc_44694_new_n2691_; 
wire _abc_44694_new_n2692_; 
wire _abc_44694_new_n2693_; 
wire _abc_44694_new_n2694_; 
wire _abc_44694_new_n2696_; 
wire _abc_44694_new_n2697_; 
wire _abc_44694_new_n2698_; 
wire _abc_44694_new_n2699_; 
wire _abc_44694_new_n2701_; 
wire _abc_44694_new_n2702_; 
wire _abc_44694_new_n2703_; 
wire _abc_44694_new_n2704_; 
wire _abc_44694_new_n2706_; 
wire _abc_44694_new_n2707_; 
wire _abc_44694_new_n2708_; 
wire _abc_44694_new_n2709_; 
wire _abc_44694_new_n2711_; 
wire _abc_44694_new_n2712_; 
wire _abc_44694_new_n2713_; 
wire _abc_44694_new_n2714_; 
wire _abc_44694_new_n2716_; 
wire _abc_44694_new_n2717_; 
wire _abc_44694_new_n2718_; 
wire _abc_44694_new_n2719_; 
wire _abc_44694_new_n2720_; 
wire _abc_44694_new_n2721_; 
wire _abc_44694_new_n2722_; 
wire _abc_44694_new_n2723_; 
wire _abc_44694_new_n2724_; 
wire _abc_44694_new_n2725_; 
wire _abc_44694_new_n2726_; 
wire _abc_44694_new_n2727_; 
wire _abc_44694_new_n2728_; 
wire _abc_44694_new_n2729_; 
wire _abc_44694_new_n2730_; 
wire _abc_44694_new_n2731_; 
wire _abc_44694_new_n2732_; 
wire _abc_44694_new_n2733_; 
wire _abc_44694_new_n2735_; 
wire _abc_44694_new_n2737_; 
wire _abc_44694_new_n2739_; 
wire _abc_44694_new_n2741_; 
wire _abc_44694_new_n2743_; 
wire _abc_44694_new_n2744_; 
wire _abc_44694_new_n2745_; 
wire _abc_44694_new_n2746_; 
wire _abc_44694_new_n2747_; 
wire _abc_44694_new_n2748_; 
wire _abc_44694_new_n2749_; 
wire _abc_44694_new_n2750_; 
wire _abc_44694_new_n2751_; 
wire _abc_44694_new_n2752_; 
wire _abc_44694_new_n2753_; 
wire _abc_44694_new_n2754_; 
wire _abc_44694_new_n2755_; 
wire _abc_44694_new_n2756_; 
wire _abc_44694_new_n2758_; 
wire _abc_44694_new_n2759_; 
wire _abc_44694_new_n2761_; 
wire _abc_44694_new_n2762_; 
wire _abc_44694_new_n2764_; 
wire _abc_44694_new_n2765_; 
wire _abc_44694_new_n2767_; 
wire _abc_44694_new_n2768_; 
wire _abc_44694_new_n2770_; 
wire _abc_44694_new_n2771_; 
wire _abc_44694_new_n2773_; 
wire _abc_44694_new_n2774_; 
wire _abc_44694_new_n2775_; 
wire _abc_44694_new_n2776_; 
wire _abc_44694_new_n2777_; 
wire _abc_44694_new_n2778_; 
wire _abc_44694_new_n2779_; 
wire _abc_44694_new_n2779__bF_buf0; 
wire _abc_44694_new_n2779__bF_buf1; 
wire _abc_44694_new_n2779__bF_buf2; 
wire _abc_44694_new_n2779__bF_buf3; 
wire _abc_44694_new_n2779__bF_buf4; 
wire _abc_44694_new_n2780_; 
wire _abc_44694_new_n2782_; 
wire _abc_44694_new_n2783_; 
wire _abc_44694_new_n2784_; 
wire _abc_44694_new_n2785_; 
wire _abc_44694_new_n2787_; 
wire _abc_44694_new_n2788_; 
wire _abc_44694_new_n2789_; 
wire _abc_44694_new_n2790_; 
wire _abc_44694_new_n2792_; 
wire _abc_44694_new_n2793_; 
wire _abc_44694_new_n2794_; 
wire _abc_44694_new_n2795_; 
wire _abc_44694_new_n2797_; 
wire _abc_44694_new_n2798_; 
wire _abc_44694_new_n2799_; 
wire _abc_44694_new_n2800_; 
wire _abc_44694_new_n2802_; 
wire _abc_44694_new_n2803_; 
wire _abc_44694_new_n2804_; 
wire _abc_44694_new_n2805_; 
wire _abc_44694_new_n2807_; 
wire _abc_44694_new_n2808_; 
wire _abc_44694_new_n2809_; 
wire _abc_44694_new_n2810_; 
wire _abc_44694_new_n2812_; 
wire _abc_44694_new_n2813_; 
wire _abc_44694_new_n2814_; 
wire _abc_44694_new_n2815_; 
wire _abc_44694_new_n2817_; 
wire _abc_44694_new_n2818_; 
wire _abc_44694_new_n2819_; 
wire _abc_44694_new_n2820_; 
wire _abc_44694_new_n2822_; 
wire _abc_44694_new_n2823_; 
wire _abc_44694_new_n2824_; 
wire _abc_44694_new_n2825_; 
wire _abc_44694_new_n2826_; 
wire _abc_44694_new_n2826__bF_buf0; 
wire _abc_44694_new_n2826__bF_buf1; 
wire _abc_44694_new_n2826__bF_buf2; 
wire _abc_44694_new_n2826__bF_buf3; 
wire _abc_44694_new_n2827_; 
wire _abc_44694_new_n2828_; 
wire _abc_44694_new_n2829_; 
wire _abc_44694_new_n2831_; 
wire _abc_44694_new_n2832_; 
wire _abc_44694_new_n2833_; 
wire _abc_44694_new_n2834_; 
wire _abc_44694_new_n2835_; 
wire _abc_44694_new_n2836_; 
wire _abc_44694_new_n2837_; 
wire _abc_44694_new_n2838_; 
wire _abc_44694_new_n2839_; 
wire _abc_44694_new_n2840_; 
wire _abc_44694_new_n2841_; 
wire _abc_44694_new_n2842_; 
wire _abc_44694_new_n2844_; 
wire _abc_44694_new_n2845_; 
wire _abc_44694_new_n2846_; 
wire _abc_44694_new_n2847_; 
wire _abc_44694_new_n2848_; 
wire _abc_44694_new_n2849_; 
wire _abc_44694_new_n2850_; 
wire _abc_44694_new_n2852_; 
wire _abc_44694_new_n2853_; 
wire _abc_44694_new_n2854_; 
wire _abc_44694_new_n2855_; 
wire _abc_44694_new_n2856_; 
wire _abc_44694_new_n2857_; 
wire _abc_44694_new_n2858_; 
wire _abc_44694_new_n2860_; 
wire _abc_44694_new_n2861_; 
wire _abc_44694_new_n2862_; 
wire _abc_44694_new_n2863_; 
wire _abc_44694_new_n2864_; 
wire _abc_44694_new_n2865_; 
wire _abc_44694_new_n2866_; 
wire _abc_44694_new_n2868_; 
wire _abc_44694_new_n2869_; 
wire _abc_44694_new_n2870_; 
wire _abc_44694_new_n2871_; 
wire _abc_44694_new_n2872_; 
wire _abc_44694_new_n2873_; 
wire _abc_44694_new_n2874_; 
wire _abc_44694_new_n2876_; 
wire _abc_44694_new_n2877_; 
wire _abc_44694_new_n2878_; 
wire _abc_44694_new_n2879_; 
wire _abc_44694_new_n2880_; 
wire _abc_44694_new_n2881_; 
wire _abc_44694_new_n2882_; 
wire _abc_44694_new_n2884_; 
wire _abc_44694_new_n2885_; 
wire _abc_44694_new_n2886_; 
wire _abc_44694_new_n2887_; 
wire _abc_44694_new_n2888_; 
wire _abc_44694_new_n2889_; 
wire _abc_44694_new_n2890_; 
wire _abc_44694_new_n2892_; 
wire _abc_44694_new_n2893_; 
wire _abc_44694_new_n2894_; 
wire _abc_44694_new_n2895_; 
wire _abc_44694_new_n2896_; 
wire _abc_44694_new_n2897_; 
wire _abc_44694_new_n2898_; 
wire _abc_44694_new_n2900_; 
wire _abc_44694_new_n2901_; 
wire _abc_44694_new_n2902_; 
wire _abc_44694_new_n2903_; 
wire _abc_44694_new_n2904_; 
wire _abc_44694_new_n2905_; 
wire _abc_44694_new_n2906_; 
wire _abc_44694_new_n2908_; 
wire _abc_44694_new_n2909_; 
wire _abc_44694_new_n2910_; 
wire _abc_44694_new_n2911_; 
wire _abc_44694_new_n2912_; 
wire _abc_44694_new_n2913_; 
wire _abc_44694_new_n2914_; 
wire _abc_44694_new_n2916_; 
wire _abc_44694_new_n2917_; 
wire _abc_44694_new_n2918_; 
wire _abc_44694_new_n2919_; 
wire _abc_44694_new_n2920_; 
wire _abc_44694_new_n2921_; 
wire _abc_44694_new_n2922_; 
wire _abc_44694_new_n2924_; 
wire _abc_44694_new_n2925_; 
wire _abc_44694_new_n2926_; 
wire _abc_44694_new_n2927_; 
wire _abc_44694_new_n2928_; 
wire _abc_44694_new_n2929_; 
wire _abc_44694_new_n2930_; 
wire _abc_44694_new_n2932_; 
wire _abc_44694_new_n2933_; 
wire _abc_44694_new_n2934_; 
wire _abc_44694_new_n2935_; 
wire _abc_44694_new_n2936_; 
wire _abc_44694_new_n2937_; 
wire _abc_44694_new_n2938_; 
wire _abc_44694_new_n2940_; 
wire _abc_44694_new_n2941_; 
wire _abc_44694_new_n2942_; 
wire _abc_44694_new_n2943_; 
wire _abc_44694_new_n2944_; 
wire _abc_44694_new_n2945_; 
wire _abc_44694_new_n2946_; 
wire _abc_44694_new_n2948_; 
wire _abc_44694_new_n2949_; 
wire _abc_44694_new_n2950_; 
wire _abc_44694_new_n2951_; 
wire _abc_44694_new_n2952_; 
wire _abc_44694_new_n2953_; 
wire _abc_44694_new_n2954_; 
wire _abc_44694_new_n2956_; 
wire _abc_44694_new_n2957_; 
wire _abc_44694_new_n2958_; 
wire _abc_44694_new_n2959_; 
wire _abc_44694_new_n2960_; 
wire _abc_44694_new_n2961_; 
wire _abc_44694_new_n2962_; 
wire _abc_44694_new_n2964_; 
wire _abc_44694_new_n2965_; 
wire _abc_44694_new_n2965__bF_buf0; 
wire _abc_44694_new_n2965__bF_buf1; 
wire _abc_44694_new_n2965__bF_buf2; 
wire _abc_44694_new_n2965__bF_buf3; 
wire _abc_44694_new_n2965__bF_buf4; 
wire _abc_44694_new_n2966_; 
wire _abc_44694_new_n2967_; 
wire _abc_44694_new_n2968_; 
wire _abc_44694_new_n2969_; 
wire _abc_44694_new_n2970_; 
wire _abc_44694_new_n2971_; 
wire _abc_44694_new_n2972_; 
wire _abc_44694_new_n2972__bF_buf0; 
wire _abc_44694_new_n2972__bF_buf1; 
wire _abc_44694_new_n2972__bF_buf2; 
wire _abc_44694_new_n2972__bF_buf3; 
wire _abc_44694_new_n2972__bF_buf4; 
wire _abc_44694_new_n2973_; 
wire _abc_44694_new_n2975_; 
wire _abc_44694_new_n2976_; 
wire _abc_44694_new_n2977_; 
wire _abc_44694_new_n2978_; 
wire _abc_44694_new_n2979_; 
wire _abc_44694_new_n2980_; 
wire _abc_44694_new_n2981_; 
wire _abc_44694_new_n2983_; 
wire _abc_44694_new_n2984_; 
wire _abc_44694_new_n2985_; 
wire _abc_44694_new_n2986_; 
wire _abc_44694_new_n2987_; 
wire _abc_44694_new_n2988_; 
wire _abc_44694_new_n2989_; 
wire _abc_44694_new_n2990_; 
wire _abc_44694_new_n2991_; 
wire _abc_44694_new_n2992_; 
wire _abc_44694_new_n2993_; 
wire _abc_44694_new_n2994_; 
wire _abc_44694_new_n2996_; 
wire _abc_44694_new_n2997_; 
wire _abc_44694_new_n2998_; 
wire _abc_44694_new_n2999_; 
wire _abc_44694_new_n3000_; 
wire _abc_44694_new_n3001_; 
wire _abc_44694_new_n3002_; 
wire _abc_44694_new_n3004_; 
wire _abc_44694_new_n3005_; 
wire _abc_44694_new_n3006_; 
wire _abc_44694_new_n3007_; 
wire _abc_44694_new_n3008_; 
wire _abc_44694_new_n3009_; 
wire _abc_44694_new_n3010_; 
wire _abc_44694_new_n3011_; 
wire _abc_44694_new_n3013_; 
wire _abc_44694_new_n3014_; 
wire _abc_44694_new_n3015_; 
wire _abc_44694_new_n3016_; 
wire _abc_44694_new_n3017_; 
wire _abc_44694_new_n3018_; 
wire _abc_44694_new_n3019_; 
wire _abc_44694_new_n3021_; 
wire _abc_44694_new_n3022_; 
wire _abc_44694_new_n3023_; 
wire _abc_44694_new_n3024_; 
wire _abc_44694_new_n3025_; 
wire _abc_44694_new_n3026_; 
wire _abc_44694_new_n3027_; 
wire _abc_44694_new_n3028_; 
wire _abc_44694_new_n3030_; 
wire _abc_44694_new_n3031_; 
wire _abc_44694_new_n3032_; 
wire _abc_44694_new_n3033_; 
wire _abc_44694_new_n3034_; 
wire _abc_44694_new_n3035_; 
wire _abc_44694_new_n3036_; 
wire _abc_44694_new_n3038_; 
wire _abc_44694_new_n3039_; 
wire _abc_44694_new_n3040_; 
wire _abc_44694_new_n3041_; 
wire _abc_44694_new_n3042_; 
wire _abc_44694_new_n3043_; 
wire _abc_44694_new_n3044_; 
wire _abc_44694_new_n3045_; 
wire _abc_44694_new_n3047_; 
wire _abc_44694_new_n3048_; 
wire _abc_44694_new_n3049_; 
wire _abc_44694_new_n3050_; 
wire _abc_44694_new_n3051_; 
wire _abc_44694_new_n3052_; 
wire _abc_44694_new_n3053_; 
wire _abc_44694_new_n3054_; 
wire _abc_44694_new_n3055_; 
wire _abc_44694_new_n3056_; 
wire _abc_44694_new_n3057_; 
wire _abc_44694_new_n3058_; 
wire _abc_44694_new_n3060_; 
wire _abc_44694_new_n3061_; 
wire _abc_44694_new_n3062_; 
wire _abc_44694_new_n3063_; 
wire _abc_44694_new_n3064_; 
wire _abc_44694_new_n3065_; 
wire _abc_44694_new_n3066_; 
wire _abc_44694_new_n3067_; 
wire _abc_44694_new_n3068_; 
wire _abc_44694_new_n3069_; 
wire _abc_44694_new_n3070_; 
wire _abc_44694_new_n3072_; 
wire _abc_44694_new_n3073_; 
wire _abc_44694_new_n3074_; 
wire _abc_44694_new_n3075_; 
wire _abc_44694_new_n3076_; 
wire _abc_44694_new_n3077_; 
wire _abc_44694_new_n3078_; 
wire _abc_44694_new_n3079_; 
wire _abc_44694_new_n3080_; 
wire _abc_44694_new_n3082_; 
wire _abc_44694_new_n3083_; 
wire _abc_44694_new_n3084_; 
wire _abc_44694_new_n3085_; 
wire _abc_44694_new_n3086_; 
wire _abc_44694_new_n3087_; 
wire _abc_44694_new_n3088_; 
wire _abc_44694_new_n3090_; 
wire _abc_44694_new_n3091_; 
wire _abc_44694_new_n3092_; 
wire _abc_44694_new_n3093_; 
wire _abc_44694_new_n3094_; 
wire _abc_44694_new_n3095_; 
wire _abc_44694_new_n3096_; 
wire _abc_44694_new_n3098_; 
wire _abc_44694_new_n3099_; 
wire _abc_44694_new_n3100_; 
wire _abc_44694_new_n3101_; 
wire _abc_44694_new_n3102_; 
wire _abc_44694_new_n3103_; 
wire _abc_44694_new_n3104_; 
wire _abc_44694_new_n3106_; 
wire _abc_44694_new_n3107_; 
wire _abc_44694_new_n3108_; 
wire _abc_44694_new_n3109_; 
wire _abc_44694_new_n3110_; 
wire _abc_44694_new_n3111_; 
wire _abc_44694_new_n3112_; 
wire _abc_44694_new_n3114_; 
wire _abc_44694_new_n3115_; 
wire _abc_44694_new_n3116_; 
wire _abc_44694_new_n3117_; 
wire _abc_44694_new_n3118_; 
wire _abc_44694_new_n3119_; 
wire _abc_44694_new_n3120_; 
wire _abc_44694_new_n3121_; 
wire _abc_44694_new_n3122_; 
wire _abc_44694_new_n3123_; 
wire _abc_44694_new_n3124_; 
wire _abc_44694_new_n3126_; 
wire _abc_44694_new_n3127_; 
wire _abc_44694_new_n3128_; 
wire _abc_44694_new_n3129_; 
wire _abc_44694_new_n3130_; 
wire _abc_44694_new_n3131_; 
wire _abc_44694_new_n3132_; 
wire _abc_44694_new_n3133_; 
wire _abc_44694_new_n3134_; 
wire _abc_44694_new_n3135_; 
wire _abc_44694_new_n3136_; 
wire _abc_44694_new_n3138_; 
wire _abc_44694_new_n3139_; 
wire _abc_44694_new_n3140_; 
wire _abc_44694_new_n3141_; 
wire _abc_44694_new_n3142_; 
wire _abc_44694_new_n3143_; 
wire _abc_44694_new_n3144_; 
wire _abc_44694_new_n3145_; 
wire _abc_44694_new_n3146_; 
wire _abc_44694_new_n3147_; 
wire _abc_44694_new_n3148_; 
wire _abc_44694_new_n3150_; 
wire _abc_44694_new_n3151_; 
wire _abc_44694_new_n3152_; 
wire _abc_44694_new_n3153_; 
wire _abc_44694_new_n3154_; 
wire _abc_44694_new_n3155_; 
wire _abc_44694_new_n3156_; 
wire _abc_44694_new_n3157_; 
wire _abc_44694_new_n3158_; 
wire _abc_44694_new_n3159_; 
wire _abc_44694_new_n3160_; 
wire _abc_44694_new_n3162_; 
wire _abc_44694_new_n3163_; 
wire _abc_44694_new_n3164_; 
wire _abc_44694_new_n3165_; 
wire _abc_44694_new_n3166_; 
wire _abc_44694_new_n3167_; 
wire _abc_44694_new_n3168_; 
wire _abc_44694_new_n3169_; 
wire _abc_44694_new_n3170_; 
wire _abc_44694_new_n3171_; 
wire _abc_44694_new_n3172_; 
wire _abc_44694_new_n3174_; 
wire _abc_44694_new_n3175_; 
wire _abc_44694_new_n3176_; 
wire _abc_44694_new_n3177_; 
wire _abc_44694_new_n3178_; 
wire _abc_44694_new_n3179_; 
wire _abc_44694_new_n3180_; 
wire _abc_44694_new_n3181_; 
wire _abc_44694_new_n3182_; 
wire _abc_44694_new_n3183_; 
wire _abc_44694_new_n3184_; 
wire _abc_44694_new_n3186_; 
wire _abc_44694_new_n3187_; 
wire _abc_44694_new_n3188_; 
wire _abc_44694_new_n3189_; 
wire _abc_44694_new_n3190_; 
wire _abc_44694_new_n3191_; 
wire _abc_44694_new_n3192_; 
wire _abc_44694_new_n3193_; 
wire _abc_44694_new_n3194_; 
wire _abc_44694_new_n3195_; 
wire _abc_44694_new_n3196_; 
wire _abc_44694_new_n3198_; 
wire _abc_44694_new_n3199_; 
wire _abc_44694_new_n3200_; 
wire _abc_44694_new_n3201_; 
wire _abc_44694_new_n3202_; 
wire _abc_44694_new_n3203_; 
wire _abc_44694_new_n3204_; 
wire _abc_44694_new_n3205_; 
wire _abc_44694_new_n3206_; 
wire _abc_44694_new_n3207_; 
wire _abc_44694_new_n3208_; 
wire _abc_44694_new_n3210_; 
wire _abc_44694_new_n3211_; 
wire _abc_44694_new_n3212_; 
wire _abc_44694_new_n3213_; 
wire _abc_44694_new_n3214_; 
wire _abc_44694_new_n3215_; 
wire _abc_44694_new_n3216_; 
wire _abc_44694_new_n3217_; 
wire _abc_44694_new_n3218_; 
wire _abc_44694_new_n3219_; 
wire _abc_44694_new_n3220_; 
wire _abc_44694_new_n3222_; 
wire _abc_44694_new_n3223_; 
wire _abc_44694_new_n3224_; 
wire _abc_44694_new_n3225_; 
wire _abc_44694_new_n3226_; 
wire _abc_44694_new_n3227_; 
wire _abc_44694_new_n3228_; 
wire _abc_44694_new_n3229_; 
wire _abc_44694_new_n3230_; 
wire _abc_44694_new_n3231_; 
wire _abc_44694_new_n3232_; 
wire _abc_44694_new_n3234_; 
wire _abc_44694_new_n3235_; 
wire _abc_44694_new_n3236_; 
wire _abc_44694_new_n3237_; 
wire _abc_44694_new_n3238_; 
wire _abc_44694_new_n3239_; 
wire _abc_44694_new_n3240_; 
wire _abc_44694_new_n3241_; 
wire _abc_44694_new_n3242_; 
wire _abc_44694_new_n3243_; 
wire _abc_44694_new_n3244_; 
wire _abc_44694_new_n3246_; 
wire _abc_44694_new_n3247_; 
wire _abc_44694_new_n3248_; 
wire _abc_44694_new_n3249_; 
wire _abc_44694_new_n3250_; 
wire _abc_44694_new_n3251_; 
wire _abc_44694_new_n3252_; 
wire _abc_44694_new_n3253_; 
wire _abc_44694_new_n3254_; 
wire _abc_44694_new_n3255_; 
wire _abc_44694_new_n3256_; 
wire _abc_44694_new_n3258_; 
wire _abc_44694_new_n3259_; 
wire _abc_44694_new_n3260_; 
wire _abc_44694_new_n3261_; 
wire _abc_44694_new_n3262_; 
wire _abc_44694_new_n3263_; 
wire _abc_44694_new_n3264_; 
wire _abc_44694_new_n3265_; 
wire _abc_44694_new_n3266_; 
wire _abc_44694_new_n3267_; 
wire _abc_44694_new_n3268_; 
wire _abc_44694_new_n3270_; 
wire _abc_44694_new_n3271_; 
wire _abc_44694_new_n3272_; 
wire _abc_44694_new_n3273_; 
wire _abc_44694_new_n3274_; 
wire _abc_44694_new_n3275_; 
wire _abc_44694_new_n3276_; 
wire _abc_44694_new_n3277_; 
wire _abc_44694_new_n3278_; 
wire _abc_44694_new_n3279_; 
wire _abc_44694_new_n3280_; 
wire _abc_44694_new_n3282_; 
wire _abc_44694_new_n3283_; 
wire _abc_44694_new_n3284_; 
wire _abc_44694_new_n3285_; 
wire _abc_44694_new_n3286_; 
wire _abc_44694_new_n3287_; 
wire _abc_44694_new_n3288_; 
wire _abc_44694_new_n3289_; 
wire _abc_44694_new_n3290_; 
wire _abc_44694_new_n3291_; 
wire _abc_44694_new_n3292_; 
wire _abc_44694_new_n3294_; 
wire _abc_44694_new_n3295_; 
wire _abc_44694_new_n3296_; 
wire _abc_44694_new_n3297_; 
wire _abc_44694_new_n3298_; 
wire _abc_44694_new_n3299_; 
wire _abc_44694_new_n3300_; 
wire _abc_44694_new_n3301_; 
wire _abc_44694_new_n3302_; 
wire _abc_44694_new_n3303_; 
wire _abc_44694_new_n3304_; 
wire _abc_44694_new_n3306_; 
wire _abc_44694_new_n3307_; 
wire _abc_44694_new_n3308_; 
wire _abc_44694_new_n3309_; 
wire _abc_44694_new_n3310_; 
wire _abc_44694_new_n3312_; 
wire _abc_44694_new_n3313_; 
wire _abc_44694_new_n3314_; 
wire _abc_44694_new_n3315_; 
wire _abc_44694_new_n3316_; 
wire _abc_44694_new_n3317_; 
wire _abc_44694_new_n3318_; 
wire _abc_44694_new_n3319_; 
wire _abc_44694_new_n3320_; 
wire _abc_44694_new_n3321_; 
wire _abc_44694_new_n3322_; 
wire _abc_44694_new_n3323_; 
wire _abc_44694_new_n3325_; 
wire _abc_44694_new_n3326_; 
wire _abc_44694_new_n3328_; 
wire _abc_44694_new_n3329_; 
wire _abc_44694_new_n3331_; 
wire _abc_44694_new_n3332_; 
wire _abc_44694_new_n3333_; 
wire _abc_44694_new_n3334_; 
wire _abc_44694_new_n3334__bF_buf0; 
wire _abc_44694_new_n3334__bF_buf1; 
wire _abc_44694_new_n3334__bF_buf2; 
wire _abc_44694_new_n3334__bF_buf3; 
wire _abc_44694_new_n3334__bF_buf4; 
wire _abc_44694_new_n3334__bF_buf5; 
wire _abc_44694_new_n3335_; 
wire _abc_44694_new_n3336_; 
wire _abc_44694_new_n3338_; 
wire _abc_44694_new_n3339_; 
wire _abc_44694_new_n3340_; 
wire _abc_44694_new_n3341_; 
wire _abc_44694_new_n3342_; 
wire _abc_44694_new_n3343_; 
wire _abc_44694_new_n3344_; 
wire _abc_44694_new_n3345_; 
wire _abc_44694_new_n3346_; 
wire _abc_44694_new_n3347_; 
wire _abc_44694_new_n3350_; 
wire _abc_44694_new_n3351_; 
wire _abc_44694_new_n3352_; 
wire _abc_44694_new_n3353_; 
wire _abc_44694_new_n3355_; 
wire _abc_44694_new_n3356_; 
wire _abc_44694_new_n3357_; 
wire _abc_44694_new_n3358_; 
wire _abc_44694_new_n3360_; 
wire _abc_44694_new_n3361_; 
wire _abc_44694_new_n3362_; 
wire _abc_44694_new_n3363_; 
wire _abc_44694_new_n3365_; 
wire _abc_44694_new_n3366_; 
wire _abc_44694_new_n3367_; 
wire _abc_44694_new_n3368_; 
wire _abc_44694_new_n3370_; 
wire _abc_44694_new_n3371_; 
wire _abc_44694_new_n3372_; 
wire _abc_44694_new_n3373_; 
wire _abc_44694_new_n3375_; 
wire _abc_44694_new_n3376_; 
wire _abc_44694_new_n3377_; 
wire _abc_44694_new_n3378_; 
wire _abc_44694_new_n3380_; 
wire _abc_44694_new_n3381_; 
wire _abc_44694_new_n3382_; 
wire _abc_44694_new_n3383_; 
wire _abc_44694_new_n3385_; 
wire _abc_44694_new_n3386_; 
wire _abc_44694_new_n3387_; 
wire _abc_44694_new_n3388_; 
wire _abc_44694_new_n3390_; 
wire _abc_44694_new_n3391_; 
wire _abc_44694_new_n3392_; 
wire _abc_44694_new_n3393_; 
wire _abc_44694_new_n3395_; 
wire _abc_44694_new_n3396_; 
wire _abc_44694_new_n3397_; 
wire _abc_44694_new_n3398_; 
wire _abc_44694_new_n3400_; 
wire _abc_44694_new_n3401_; 
wire _abc_44694_new_n3402_; 
wire _abc_44694_new_n3403_; 
wire _abc_44694_new_n3405_; 
wire _abc_44694_new_n3406_; 
wire _abc_44694_new_n3407_; 
wire _abc_44694_new_n3408_; 
wire _abc_44694_new_n3410_; 
wire _abc_44694_new_n3411_; 
wire _abc_44694_new_n3412_; 
wire _abc_44694_new_n3413_; 
wire _abc_44694_new_n3415_; 
wire _abc_44694_new_n3416_; 
wire _abc_44694_new_n3417_; 
wire _abc_44694_new_n3418_; 
wire _abc_44694_new_n3420_; 
wire _abc_44694_new_n3421_; 
wire _abc_44694_new_n3422_; 
wire _abc_44694_new_n3423_; 
wire _abc_44694_new_n3425_; 
wire _abc_44694_new_n3426_; 
wire _abc_44694_new_n3427_; 
wire _abc_44694_new_n3428_; 
wire _abc_44694_new_n3430_; 
wire _abc_44694_new_n3431_; 
wire _abc_44694_new_n3432_; 
wire _abc_44694_new_n3433_; 
wire _abc_44694_new_n3435_; 
wire _abc_44694_new_n3436_; 
wire _abc_44694_new_n3437_; 
wire _abc_44694_new_n3438_; 
wire _abc_44694_new_n3440_; 
wire _abc_44694_new_n3441_; 
wire _abc_44694_new_n3442_; 
wire _abc_44694_new_n3443_; 
wire _abc_44694_new_n3445_; 
wire _abc_44694_new_n3446_; 
wire _abc_44694_new_n3447_; 
wire _abc_44694_new_n3448_; 
wire _abc_44694_new_n3450_; 
wire _abc_44694_new_n3451_; 
wire _abc_44694_new_n3452_; 
wire _abc_44694_new_n3453_; 
wire _abc_44694_new_n3455_; 
wire _abc_44694_new_n3456_; 
wire _abc_44694_new_n3457_; 
wire _abc_44694_new_n3458_; 
wire _abc_44694_new_n3460_; 
wire _abc_44694_new_n3461_; 
wire _abc_44694_new_n3462_; 
wire _abc_44694_new_n3463_; 
wire _abc_44694_new_n3465_; 
wire _abc_44694_new_n3466_; 
wire _abc_44694_new_n3467_; 
wire _abc_44694_new_n3468_; 
wire _abc_44694_new_n3470_; 
wire _abc_44694_new_n3471_; 
wire _abc_44694_new_n3472_; 
wire _abc_44694_new_n3473_; 
wire _abc_44694_new_n3475_; 
wire _abc_44694_new_n3476_; 
wire _abc_44694_new_n3477_; 
wire _abc_44694_new_n3478_; 
wire _abc_44694_new_n3480_; 
wire _abc_44694_new_n3481_; 
wire _abc_44694_new_n3482_; 
wire _abc_44694_new_n3483_; 
wire _abc_44694_new_n3485_; 
wire _abc_44694_new_n3486_; 
wire _abc_44694_new_n3487_; 
wire _abc_44694_new_n3488_; 
wire _abc_44694_new_n3490_; 
wire _abc_44694_new_n3491_; 
wire _abc_44694_new_n3492_; 
wire _abc_44694_new_n3493_; 
wire _abc_44694_new_n3495_; 
wire _abc_44694_new_n3496_; 
wire _abc_44694_new_n3497_; 
wire _abc_44694_new_n3498_; 
wire _abc_44694_new_n3500_; 
wire _abc_44694_new_n3501_; 
wire _abc_44694_new_n3502_; 
wire _abc_44694_new_n3503_; 
wire _abc_44694_new_n3505_; 
wire _abc_44694_new_n3506_; 
wire _abc_44694_new_n3507_; 
wire _abc_44694_new_n3508_; 
wire _abc_44694_new_n3510_; 
wire _abc_44694_new_n3511_; 
wire _abc_44694_new_n3512_; 
wire _abc_44694_new_n3512__bF_buf0; 
wire _abc_44694_new_n3512__bF_buf1; 
wire _abc_44694_new_n3512__bF_buf2; 
wire _abc_44694_new_n3512__bF_buf3; 
wire _abc_44694_new_n3512__bF_buf4; 
wire _abc_44694_new_n3513_; 
wire _abc_44694_new_n3513__bF_buf0; 
wire _abc_44694_new_n3513__bF_buf1; 
wire _abc_44694_new_n3513__bF_buf2; 
wire _abc_44694_new_n3513__bF_buf3; 
wire _abc_44694_new_n3513__bF_buf4; 
wire _abc_44694_new_n3514_; 
wire _abc_44694_new_n3515_; 
wire _abc_44694_new_n3515__bF_buf0; 
wire _abc_44694_new_n3515__bF_buf1; 
wire _abc_44694_new_n3515__bF_buf2; 
wire _abc_44694_new_n3515__bF_buf3; 
wire _abc_44694_new_n3516_; 
wire _abc_44694_new_n3517_; 
wire _abc_44694_new_n3518_; 
wire _abc_44694_new_n3518__bF_buf0; 
wire _abc_44694_new_n3518__bF_buf1; 
wire _abc_44694_new_n3518__bF_buf2; 
wire _abc_44694_new_n3518__bF_buf3; 
wire _abc_44694_new_n3519_; 
wire _abc_44694_new_n3519__bF_buf0; 
wire _abc_44694_new_n3519__bF_buf1; 
wire _abc_44694_new_n3519__bF_buf2; 
wire _abc_44694_new_n3519__bF_buf3; 
wire _abc_44694_new_n3519__bF_buf4; 
wire _abc_44694_new_n3520_; 
wire _abc_44694_new_n3520__bF_buf0; 
wire _abc_44694_new_n3520__bF_buf1; 
wire _abc_44694_new_n3520__bF_buf2; 
wire _abc_44694_new_n3520__bF_buf3; 
wire _abc_44694_new_n3520__bF_buf4; 
wire _abc_44694_new_n3521_; 
wire _abc_44694_new_n3521__bF_buf0; 
wire _abc_44694_new_n3521__bF_buf1; 
wire _abc_44694_new_n3521__bF_buf2; 
wire _abc_44694_new_n3521__bF_buf3; 
wire _abc_44694_new_n3521__bF_buf4; 
wire _abc_44694_new_n3522_; 
wire _abc_44694_new_n3523_; 
wire _abc_44694_new_n3524_; 
wire _abc_44694_new_n3525_; 
wire _abc_44694_new_n3526_; 
wire _abc_44694_new_n3527_; 
wire _abc_44694_new_n3527__bF_buf0; 
wire _abc_44694_new_n3527__bF_buf1; 
wire _abc_44694_new_n3527__bF_buf2; 
wire _abc_44694_new_n3527__bF_buf3; 
wire _abc_44694_new_n3527__bF_buf4; 
wire _abc_44694_new_n3528_; 
wire _abc_44694_new_n3529_; 
wire _abc_44694_new_n3530_; 
wire _abc_44694_new_n3531_; 
wire _abc_44694_new_n3532_; 
wire _abc_44694_new_n3534_; 
wire _abc_44694_new_n3535_; 
wire _abc_44694_new_n3536_; 
wire _abc_44694_new_n3537_; 
wire _abc_44694_new_n3538_; 
wire _abc_44694_new_n3539_; 
wire _abc_44694_new_n3540_; 
wire _abc_44694_new_n3541_; 
wire _abc_44694_new_n3542_; 
wire _abc_44694_new_n3544_; 
wire _abc_44694_new_n3545_; 
wire _abc_44694_new_n3546_; 
wire _abc_44694_new_n3546__bF_buf0; 
wire _abc_44694_new_n3546__bF_buf1; 
wire _abc_44694_new_n3546__bF_buf2; 
wire _abc_44694_new_n3546__bF_buf3; 
wire _abc_44694_new_n3547_; 
wire _abc_44694_new_n3548_; 
wire _abc_44694_new_n3549_; 
wire _abc_44694_new_n3550_; 
wire _abc_44694_new_n3551_; 
wire _abc_44694_new_n3552_; 
wire _abc_44694_new_n3553_; 
wire _abc_44694_new_n3554_; 
wire _abc_44694_new_n3556_; 
wire _abc_44694_new_n3557_; 
wire _abc_44694_new_n3558_; 
wire _abc_44694_new_n3559_; 
wire _abc_44694_new_n3560_; 
wire _abc_44694_new_n3561_; 
wire _abc_44694_new_n3563_; 
wire _abc_44694_new_n3563__bF_buf0; 
wire _abc_44694_new_n3563__bF_buf1; 
wire _abc_44694_new_n3563__bF_buf2; 
wire _abc_44694_new_n3563__bF_buf3; 
wire _abc_44694_new_n3563__bF_buf4; 
wire _abc_44694_new_n3564_; 
wire _abc_44694_new_n3565_; 
wire _abc_44694_new_n3566_; 
wire _abc_44694_new_n3567_; 
wire _abc_44694_new_n3568_; 
wire _abc_44694_new_n3569_; 
wire _abc_44694_new_n3570_; 
wire _abc_44694_new_n3571_; 
wire _abc_44694_new_n3572_; 
wire _abc_44694_new_n3573_; 
wire _abc_44694_new_n3574_; 
wire _abc_44694_new_n3575_; 
wire _abc_44694_new_n3576_; 
wire _abc_44694_new_n3577_; 
wire _abc_44694_new_n3579_; 
wire _abc_44694_new_n3580_; 
wire _abc_44694_new_n3581_; 
wire _abc_44694_new_n3582_; 
wire _abc_44694_new_n3583_; 
wire _abc_44694_new_n3584_; 
wire _abc_44694_new_n3585_; 
wire _abc_44694_new_n3586_; 
wire _abc_44694_new_n3587_; 
wire _abc_44694_new_n3588_; 
wire _abc_44694_new_n3589_; 
wire _abc_44694_new_n3590_; 
wire _abc_44694_new_n3591_; 
wire _abc_44694_new_n3592_; 
wire _abc_44694_new_n3594_; 
wire _abc_44694_new_n3595_; 
wire _abc_44694_new_n3596_; 
wire _abc_44694_new_n3597_; 
wire _abc_44694_new_n3598_; 
wire _abc_44694_new_n3599_; 
wire _abc_44694_new_n3600_; 
wire _abc_44694_new_n3601_; 
wire _abc_44694_new_n3602_; 
wire _abc_44694_new_n3603_; 
wire _abc_44694_new_n3604_; 
wire _abc_44694_new_n3605_; 
wire _abc_44694_new_n3606_; 
wire _abc_44694_new_n3607_; 
wire _abc_44694_new_n3609_; 
wire _abc_44694_new_n3610_; 
wire _abc_44694_new_n3611_; 
wire _abc_44694_new_n3612_; 
wire _abc_44694_new_n3613_; 
wire _abc_44694_new_n3614_; 
wire _abc_44694_new_n3615_; 
wire _abc_44694_new_n3616_; 
wire _abc_44694_new_n3617_; 
wire _abc_44694_new_n3618_; 
wire _abc_44694_new_n3619_; 
wire _abc_44694_new_n3620_; 
wire _abc_44694_new_n3621_; 
wire _abc_44694_new_n3622_; 
wire _abc_44694_new_n3624_; 
wire _abc_44694_new_n3625_; 
wire _abc_44694_new_n3626_; 
wire _abc_44694_new_n3627_; 
wire _abc_44694_new_n3628_; 
wire _abc_44694_new_n3629_; 
wire _abc_44694_new_n3630_; 
wire _abc_44694_new_n3631_; 
wire _abc_44694_new_n3632_; 
wire _abc_44694_new_n3633_; 
wire _abc_44694_new_n3634_; 
wire _abc_44694_new_n3635_; 
wire _abc_44694_new_n3636_; 
wire _abc_44694_new_n3637_; 
wire _abc_44694_new_n3639_; 
wire _abc_44694_new_n3640_; 
wire _abc_44694_new_n3641_; 
wire _abc_44694_new_n3642_; 
wire _abc_44694_new_n3643_; 
wire _abc_44694_new_n3644_; 
wire _abc_44694_new_n3645_; 
wire _abc_44694_new_n3646_; 
wire _abc_44694_new_n3647_; 
wire _abc_44694_new_n3648_; 
wire _abc_44694_new_n3649_; 
wire _abc_44694_new_n3650_; 
wire _abc_44694_new_n3651_; 
wire _abc_44694_new_n3652_; 
wire _abc_44694_new_n3654_; 
wire _abc_44694_new_n3655_; 
wire _abc_44694_new_n3656_; 
wire _abc_44694_new_n3657_; 
wire _abc_44694_new_n3658_; 
wire _abc_44694_new_n3659_; 
wire _abc_44694_new_n3660_; 
wire _abc_44694_new_n3661_; 
wire _abc_44694_new_n3662_; 
wire _abc_44694_new_n3663_; 
wire _abc_44694_new_n3664_; 
wire _abc_44694_new_n3665_; 
wire _abc_44694_new_n3666_; 
wire _abc_44694_new_n3667_; 
wire _abc_44694_new_n3669_; 
wire _abc_44694_new_n3670_; 
wire _abc_44694_new_n3671_; 
wire _abc_44694_new_n3672_; 
wire _abc_44694_new_n3673_; 
wire _abc_44694_new_n3674_; 
wire _abc_44694_new_n3675_; 
wire _abc_44694_new_n3676_; 
wire _abc_44694_new_n3677_; 
wire _abc_44694_new_n3678_; 
wire _abc_44694_new_n3679_; 
wire _abc_44694_new_n3680_; 
wire _abc_44694_new_n3681_; 
wire _abc_44694_new_n3682_; 
wire _abc_44694_new_n3684_; 
wire _abc_44694_new_n3685_; 
wire _abc_44694_new_n3686_; 
wire _abc_44694_new_n3687_; 
wire _abc_44694_new_n3688_; 
wire _abc_44694_new_n3689_; 
wire _abc_44694_new_n3690_; 
wire _abc_44694_new_n3691_; 
wire _abc_44694_new_n3692_; 
wire _abc_44694_new_n3693_; 
wire _abc_44694_new_n3694_; 
wire _abc_44694_new_n3695_; 
wire _abc_44694_new_n3696_; 
wire _abc_44694_new_n3697_; 
wire _abc_44694_new_n3699_; 
wire _abc_44694_new_n3700_; 
wire _abc_44694_new_n3701_; 
wire _abc_44694_new_n3702_; 
wire _abc_44694_new_n3703_; 
wire _abc_44694_new_n3704_; 
wire _abc_44694_new_n3705_; 
wire _abc_44694_new_n3706_; 
wire _abc_44694_new_n3707_; 
wire _abc_44694_new_n3708_; 
wire _abc_44694_new_n3709_; 
wire _abc_44694_new_n3710_; 
wire _abc_44694_new_n3711_; 
wire _abc_44694_new_n3712_; 
wire _abc_44694_new_n3714_; 
wire _abc_44694_new_n3715_; 
wire _abc_44694_new_n3716_; 
wire _abc_44694_new_n3717_; 
wire _abc_44694_new_n3718_; 
wire _abc_44694_new_n3719_; 
wire _abc_44694_new_n3720_; 
wire _abc_44694_new_n3721_; 
wire _abc_44694_new_n3722_; 
wire _abc_44694_new_n3723_; 
wire _abc_44694_new_n3724_; 
wire _abc_44694_new_n3725_; 
wire _abc_44694_new_n3726_; 
wire _abc_44694_new_n3727_; 
wire _abc_44694_new_n3729_; 
wire _abc_44694_new_n3730_; 
wire _abc_44694_new_n3731_; 
wire _abc_44694_new_n3732_; 
wire _abc_44694_new_n3733_; 
wire _abc_44694_new_n3734_; 
wire _abc_44694_new_n3735_; 
wire _abc_44694_new_n3736_; 
wire _abc_44694_new_n3737_; 
wire _abc_44694_new_n3738_; 
wire _abc_44694_new_n3739_; 
wire _abc_44694_new_n3740_; 
wire _abc_44694_new_n3741_; 
wire _abc_44694_new_n3742_; 
wire _abc_44694_new_n3744_; 
wire _abc_44694_new_n3745_; 
wire _abc_44694_new_n3746_; 
wire _abc_44694_new_n3747_; 
wire _abc_44694_new_n3748_; 
wire _abc_44694_new_n3749_; 
wire _abc_44694_new_n3750_; 
wire _abc_44694_new_n3751_; 
wire _abc_44694_new_n3752_; 
wire _abc_44694_new_n3753_; 
wire _abc_44694_new_n3754_; 
wire _abc_44694_new_n3755_; 
wire _abc_44694_new_n3756_; 
wire _abc_44694_new_n3757_; 
wire _abc_44694_new_n3759_; 
wire _abc_44694_new_n3760_; 
wire _abc_44694_new_n3761_; 
wire _abc_44694_new_n3762_; 
wire _abc_44694_new_n3763_; 
wire _abc_44694_new_n3764_; 
wire _abc_44694_new_n3765_; 
wire _abc_44694_new_n3766_; 
wire _abc_44694_new_n3767_; 
wire _abc_44694_new_n3768_; 
wire _abc_44694_new_n3769_; 
wire _abc_44694_new_n3770_; 
wire _abc_44694_new_n3771_; 
wire _abc_44694_new_n3772_; 
wire _abc_44694_new_n3774_; 
wire _abc_44694_new_n3775_; 
wire _abc_44694_new_n3776_; 
wire _abc_44694_new_n3777_; 
wire _abc_44694_new_n3778_; 
wire _abc_44694_new_n3779_; 
wire _abc_44694_new_n3780_; 
wire _abc_44694_new_n3781_; 
wire _abc_44694_new_n3782_; 
wire _abc_44694_new_n3783_; 
wire _abc_44694_new_n3784_; 
wire _abc_44694_new_n3785_; 
wire _abc_44694_new_n3786_; 
wire _abc_44694_new_n3787_; 
wire _abc_44694_new_n3789_; 
wire _abc_44694_new_n3790_; 
wire _abc_44694_new_n3791_; 
wire _abc_44694_new_n3792_; 
wire _abc_44694_new_n3793_; 
wire _abc_44694_new_n3794_; 
wire _abc_44694_new_n3795_; 
wire _abc_44694_new_n3796_; 
wire _abc_44694_new_n3797_; 
wire _abc_44694_new_n3798_; 
wire _abc_44694_new_n3799_; 
wire _abc_44694_new_n3800_; 
wire _abc_44694_new_n3801_; 
wire _abc_44694_new_n3802_; 
wire _abc_44694_new_n3804_; 
wire _abc_44694_new_n3805_; 
wire _abc_44694_new_n3806_; 
wire _abc_44694_new_n3807_; 
wire _abc_44694_new_n3808_; 
wire _abc_44694_new_n3809_; 
wire _abc_44694_new_n3810_; 
wire _abc_44694_new_n3811_; 
wire _abc_44694_new_n3812_; 
wire _abc_44694_new_n3813_; 
wire _abc_44694_new_n3814_; 
wire _abc_44694_new_n3815_; 
wire _abc_44694_new_n3816_; 
wire _abc_44694_new_n3817_; 
wire _abc_44694_new_n3819_; 
wire _abc_44694_new_n3820_; 
wire _abc_44694_new_n3821_; 
wire _abc_44694_new_n3822_; 
wire _abc_44694_new_n3823_; 
wire _abc_44694_new_n3824_; 
wire _abc_44694_new_n3825_; 
wire _abc_44694_new_n3826_; 
wire _abc_44694_new_n3827_; 
wire _abc_44694_new_n3828_; 
wire _abc_44694_new_n3829_; 
wire _abc_44694_new_n3830_; 
wire _abc_44694_new_n3831_; 
wire _abc_44694_new_n3832_; 
wire _abc_44694_new_n3834_; 
wire _abc_44694_new_n3835_; 
wire _abc_44694_new_n3836_; 
wire _abc_44694_new_n3837_; 
wire _abc_44694_new_n3838_; 
wire _abc_44694_new_n3839_; 
wire _abc_44694_new_n3840_; 
wire _abc_44694_new_n3841_; 
wire _abc_44694_new_n3842_; 
wire _abc_44694_new_n3843_; 
wire _abc_44694_new_n3844_; 
wire _abc_44694_new_n3845_; 
wire _abc_44694_new_n3846_; 
wire _abc_44694_new_n3847_; 
wire _abc_44694_new_n3849_; 
wire _abc_44694_new_n3850_; 
wire _abc_44694_new_n3851_; 
wire _abc_44694_new_n3852_; 
wire _abc_44694_new_n3853_; 
wire _abc_44694_new_n3854_; 
wire _abc_44694_new_n3855_; 
wire _abc_44694_new_n3856_; 
wire _abc_44694_new_n3857_; 
wire _abc_44694_new_n3858_; 
wire _abc_44694_new_n3859_; 
wire _abc_44694_new_n3860_; 
wire _abc_44694_new_n3861_; 
wire _abc_44694_new_n3862_; 
wire _abc_44694_new_n3864_; 
wire _abc_44694_new_n3865_; 
wire _abc_44694_new_n3866_; 
wire _abc_44694_new_n3867_; 
wire _abc_44694_new_n3868_; 
wire _abc_44694_new_n3869_; 
wire _abc_44694_new_n3870_; 
wire _abc_44694_new_n3871_; 
wire _abc_44694_new_n3872_; 
wire _abc_44694_new_n3873_; 
wire _abc_44694_new_n3874_; 
wire _abc_44694_new_n3875_; 
wire _abc_44694_new_n3876_; 
wire _abc_44694_new_n3877_; 
wire _abc_44694_new_n3879_; 
wire _abc_44694_new_n3880_; 
wire _abc_44694_new_n3881_; 
wire _abc_44694_new_n3882_; 
wire _abc_44694_new_n3883_; 
wire _abc_44694_new_n3884_; 
wire _abc_44694_new_n3885_; 
wire _abc_44694_new_n3886_; 
wire _abc_44694_new_n3887_; 
wire _abc_44694_new_n3888_; 
wire _abc_44694_new_n3889_; 
wire _abc_44694_new_n3890_; 
wire _abc_44694_new_n3891_; 
wire _abc_44694_new_n3892_; 
wire _abc_44694_new_n3894_; 
wire _abc_44694_new_n3895_; 
wire _abc_44694_new_n3896_; 
wire _abc_44694_new_n3897_; 
wire _abc_44694_new_n3898_; 
wire _abc_44694_new_n3899_; 
wire _abc_44694_new_n3900_; 
wire _abc_44694_new_n3901_; 
wire _abc_44694_new_n3902_; 
wire _abc_44694_new_n3903_; 
wire _abc_44694_new_n3904_; 
wire _abc_44694_new_n3905_; 
wire _abc_44694_new_n3906_; 
wire _abc_44694_new_n3907_; 
wire _abc_44694_new_n3909_; 
wire _abc_44694_new_n3910_; 
wire _abc_44694_new_n3911_; 
wire _abc_44694_new_n3912_; 
wire _abc_44694_new_n3913_; 
wire _abc_44694_new_n3914_; 
wire _abc_44694_new_n3915_; 
wire _abc_44694_new_n3916_; 
wire _abc_44694_new_n3917_; 
wire _abc_44694_new_n3918_; 
wire _abc_44694_new_n3919_; 
wire _abc_44694_new_n3920_; 
wire _abc_44694_new_n3921_; 
wire _abc_44694_new_n3922_; 
wire _abc_44694_new_n3924_; 
wire _abc_44694_new_n3925_; 
wire _abc_44694_new_n3926_; 
wire _abc_44694_new_n3927_; 
wire _abc_44694_new_n3928_; 
wire _abc_44694_new_n3929_; 
wire _abc_44694_new_n3930_; 
wire _abc_44694_new_n3931_; 
wire _abc_44694_new_n3932_; 
wire _abc_44694_new_n3933_; 
wire _abc_44694_new_n3934_; 
wire _abc_44694_new_n3935_; 
wire _abc_44694_new_n3936_; 
wire _abc_44694_new_n3937_; 
wire _abc_44694_new_n3939_; 
wire _abc_44694_new_n3940_; 
wire _abc_44694_new_n3941_; 
wire _abc_44694_new_n3942_; 
wire _abc_44694_new_n3943_; 
wire _abc_44694_new_n3944_; 
wire _abc_44694_new_n3945_; 
wire _abc_44694_new_n3946_; 
wire _abc_44694_new_n3947_; 
wire _abc_44694_new_n3948_; 
wire _abc_44694_new_n3949_; 
wire _abc_44694_new_n3950_; 
wire _abc_44694_new_n3951_; 
wire _abc_44694_new_n3952_; 
wire _abc_44694_new_n3954_; 
wire _abc_44694_new_n3955_; 
wire _abc_44694_new_n3956_; 
wire _abc_44694_new_n3957_; 
wire _abc_44694_new_n3958_; 
wire _abc_44694_new_n3959_; 
wire _abc_44694_new_n3960_; 
wire _abc_44694_new_n3961_; 
wire _abc_44694_new_n3962_; 
wire _abc_44694_new_n3963_; 
wire _abc_44694_new_n3964_; 
wire _abc_44694_new_n3965_; 
wire _abc_44694_new_n3966_; 
wire _abc_44694_new_n3967_; 
wire _abc_44694_new_n3969_; 
wire _abc_44694_new_n3970_; 
wire _abc_44694_new_n3971_; 
wire _abc_44694_new_n3972_; 
wire _abc_44694_new_n3973_; 
wire _abc_44694_new_n3974_; 
wire _abc_44694_new_n3975_; 
wire _abc_44694_new_n3976_; 
wire _abc_44694_new_n3977_; 
wire _abc_44694_new_n3978_; 
wire _abc_44694_new_n3979_; 
wire _abc_44694_new_n3980_; 
wire _abc_44694_new_n3981_; 
wire _abc_44694_new_n3982_; 
wire _abc_44694_new_n3984_; 
wire _abc_44694_new_n3985_; 
wire _abc_44694_new_n3986_; 
wire _abc_44694_new_n3987_; 
wire _abc_44694_new_n3988_; 
wire _abc_44694_new_n3989_; 
wire _abc_44694_new_n3990_; 
wire _abc_44694_new_n3991_; 
wire _abc_44694_new_n3992_; 
wire _abc_44694_new_n3993_; 
wire _abc_44694_new_n3994_; 
wire _abc_44694_new_n3995_; 
wire _abc_44694_new_n3996_; 
wire _abc_44694_new_n3997_; 
wire _abc_44694_new_n3999_; 
wire _abc_44694_new_n4000_; 
wire _abc_44694_new_n4001_; 
wire _abc_44694_new_n4002_; 
wire _abc_44694_new_n4003_; 
wire _abc_44694_new_n4004_; 
wire _abc_44694_new_n4005_; 
wire _abc_44694_new_n4006_; 
wire _abc_44694_new_n4007_; 
wire _abc_44694_new_n4008_; 
wire _abc_44694_new_n4009_; 
wire _abc_44694_new_n4010_; 
wire _abc_44694_new_n4011_; 
wire _abc_44694_new_n4012_; 
wire _abc_44694_new_n4014_; 
wire _abc_44694_new_n4015_; 
wire _abc_44694_new_n4016_; 
wire _abc_44694_new_n4017_; 
wire _abc_44694_new_n4018_; 
wire _abc_44694_new_n4019_; 
wire _abc_44694_new_n4020_; 
wire _abc_44694_new_n4021_; 
wire _abc_44694_new_n4022_; 
wire _abc_44694_new_n4023_; 
wire _abc_44694_new_n4024_; 
wire _abc_44694_new_n4025_; 
wire _abc_44694_new_n4026_; 
wire _abc_44694_new_n4027_; 
wire _abc_44694_new_n4029_; 
wire _abc_44694_new_n4030_; 
wire _abc_44694_new_n4031_; 
wire _abc_44694_new_n4032_; 
wire _abc_44694_new_n4033_; 
wire _abc_44694_new_n4034_; 
wire _abc_44694_new_n4035_; 
wire _abc_44694_new_n4036_; 
wire _abc_44694_new_n4037_; 
wire _abc_44694_new_n4038_; 
wire _abc_44694_new_n4039_; 
wire _abc_44694_new_n4040_; 
wire _abc_44694_new_n4041_; 
wire _abc_44694_new_n4042_; 
wire _abc_44694_new_n4044_; 
wire _abc_44694_new_n4045_; 
wire _abc_44694_new_n4046_; 
wire _abc_44694_new_n4047_; 
wire _abc_44694_new_n4048_; 
wire _abc_44694_new_n4049_; 
wire _abc_44694_new_n4051_; 
wire _abc_44694_new_n4052_; 
wire _abc_44694_new_n4053_; 
wire _abc_44694_new_n4054_; 
wire _abc_44694_new_n4056_; 
wire _abc_44694_new_n4057_; 
wire _abc_44694_new_n4058_; 
wire _abc_44694_new_n4059_; 
wire _abc_44694_new_n4060_; 
wire _abc_44694_new_n4061_; 
wire _abc_44694_new_n4063_; 
wire _abc_44694_new_n4064_; 
wire _abc_44694_new_n4064__bF_buf0; 
wire _abc_44694_new_n4064__bF_buf1; 
wire _abc_44694_new_n4064__bF_buf2; 
wire _abc_44694_new_n4064__bF_buf3; 
wire _abc_44694_new_n4064__bF_buf4; 
wire _abc_44694_new_n4065_; 
wire _abc_44694_new_n4067_; 
wire _abc_44694_new_n4068_; 
wire _abc_44694_new_n4070_; 
wire _abc_44694_new_n4071_; 
wire _abc_44694_new_n4072_; 
wire _abc_44694_new_n4073_; 
wire _abc_44694_new_n4074_; 
wire _abc_44694_new_n4075_; 
wire _abc_44694_new_n4076_; 
wire _abc_44694_new_n4077_; 
wire _abc_44694_new_n4078_; 
wire _abc_44694_new_n4079_; 
wire _abc_44694_new_n4080_; 
wire _abc_44694_new_n4081_; 
wire _abc_44694_new_n4083_; 
wire _abc_44694_new_n4084_; 
wire _abc_44694_new_n4085_; 
wire _abc_44694_new_n4086_; 
wire _abc_44694_new_n4087_; 
wire _abc_44694_new_n4088_; 
wire _abc_44694_new_n4089_; 
wire _abc_44694_new_n4090_; 
wire _abc_44694_new_n4091_; 
wire _abc_44694_new_n4092_; 
wire _abc_44694_new_n4093_; 
wire _abc_44694_new_n4094_; 
wire _abc_44694_new_n4095_; 
wire _abc_44694_new_n4097_; 
wire _abc_44694_new_n4098_; 
wire _abc_44694_new_n4099_; 
wire _abc_44694_new_n4100_; 
wire _abc_44694_new_n4101_; 
wire _abc_44694_new_n4102_; 
wire _abc_44694_new_n4103_; 
wire _abc_44694_new_n4104_; 
wire _abc_44694_new_n4105_; 
wire _abc_44694_new_n4106_; 
wire _abc_44694_new_n4107_; 
wire _abc_44694_new_n4108_; 
wire _abc_44694_new_n4109_; 
wire _abc_44694_new_n4110_; 
wire _abc_44694_new_n4112_; 
wire _abc_44694_new_n4113_; 
wire _abc_44694_new_n4114_; 
wire _abc_44694_new_n4115_; 
wire _abc_44694_new_n4116_; 
wire _abc_44694_new_n4117_; 
wire _abc_44694_new_n4118_; 
wire _abc_44694_new_n4119_; 
wire _abc_44694_new_n4120_; 
wire _abc_44694_new_n4121_; 
wire _abc_44694_new_n4122_; 
wire _abc_44694_new_n4123_; 
wire _abc_44694_new_n4124_; 
wire _abc_44694_new_n4126_; 
wire _abc_44694_new_n4127_; 
wire _abc_44694_new_n4128_; 
wire _abc_44694_new_n4129_; 
wire _abc_44694_new_n4130_; 
wire _abc_44694_new_n4131_; 
wire _abc_44694_new_n4132_; 
wire _abc_44694_new_n4133_; 
wire _abc_44694_new_n4134_; 
wire _abc_44694_new_n4135_; 
wire _abc_44694_new_n4136_; 
wire _abc_44694_new_n4137_; 
wire _abc_44694_new_n4138_; 
wire _abc_44694_new_n4140_; 
wire _abc_44694_new_n4141_; 
wire _abc_44694_new_n4142_; 
wire _abc_44694_new_n4143_; 
wire _abc_44694_new_n4144_; 
wire _abc_44694_new_n4145_; 
wire _abc_44694_new_n4146_; 
wire _abc_44694_new_n4147_; 
wire _abc_44694_new_n4148_; 
wire _abc_44694_new_n4149_; 
wire _abc_44694_new_n4150_; 
wire _abc_44694_new_n4151_; 
wire _abc_44694_new_n4152_; 
wire _abc_44694_new_n4153_; 
wire _abc_44694_new_n4154_; 
wire _abc_44694_new_n4155_; 
wire _abc_44694_new_n4157_; 
wire _abc_44694_new_n4158_; 
wire _abc_44694_new_n4159_; 
wire _abc_44694_new_n4160_; 
wire _abc_44694_new_n4161_; 
wire _abc_44694_new_n4162_; 
wire _abc_44694_new_n4163_; 
wire _abc_44694_new_n4164_; 
wire _abc_44694_new_n4165_; 
wire _abc_44694_new_n4166_; 
wire _abc_44694_new_n4167_; 
wire _abc_44694_new_n4168_; 
wire _abc_44694_new_n4169_; 
wire _abc_44694_new_n4170_; 
wire _abc_44694_new_n4171_; 
wire _abc_44694_new_n4172_; 
wire _abc_44694_new_n4173_; 
wire _abc_44694_new_n4174_; 
wire _abc_44694_new_n4175_; 
wire _abc_44694_new_n4177_; 
wire _abc_44694_new_n4178_; 
wire _abc_44694_new_n4179_; 
wire _abc_44694_new_n4180_; 
wire _abc_44694_new_n4181_; 
wire _abc_44694_new_n4182_; 
wire _abc_44694_new_n4183_; 
wire _abc_44694_new_n4184_; 
wire _abc_44694_new_n4185_; 
wire _abc_44694_new_n4186_; 
wire _abc_44694_new_n4187_; 
wire _abc_44694_new_n4188_; 
wire _abc_44694_new_n4189_; 
wire _abc_44694_new_n4191_; 
wire _abc_44694_new_n4192_; 
wire _abc_44694_new_n4193_; 
wire _abc_44694_new_n4194_; 
wire _abc_44694_new_n4195_; 
wire _abc_44694_new_n4196_; 
wire _abc_44694_new_n4197_; 
wire _abc_44694_new_n4198_; 
wire _abc_44694_new_n4199_; 
wire _abc_44694_new_n4200_; 
wire _abc_44694_new_n4201_; 
wire _abc_44694_new_n4202_; 
wire _abc_44694_new_n4203_; 
wire _abc_44694_new_n4204_; 
wire _abc_44694_new_n4205_; 
wire _abc_44694_new_n4206_; 
wire _abc_44694_new_n4207_; 
wire _abc_44694_new_n4208_; 
wire _abc_44694_new_n4209_; 
wire _abc_44694_new_n4211_; 
wire _abc_44694_new_n4212_; 
wire _abc_44694_new_n4213_; 
wire _abc_44694_new_n4214_; 
wire _abc_44694_new_n4215_; 
wire _abc_44694_new_n4216_; 
wire _abc_44694_new_n4217_; 
wire _abc_44694_new_n4218_; 
wire _abc_44694_new_n4219_; 
wire _abc_44694_new_n4220_; 
wire _abc_44694_new_n4221_; 
wire _abc_44694_new_n4222_; 
wire _abc_44694_new_n4223_; 
wire _abc_44694_new_n4224_; 
wire _abc_44694_new_n4225_; 
wire _abc_44694_new_n4226_; 
wire _abc_44694_new_n4227_; 
wire _abc_44694_new_n4229_; 
wire _abc_44694_new_n4230_; 
wire _abc_44694_new_n4231_; 
wire _abc_44694_new_n4232_; 
wire _abc_44694_new_n4233_; 
wire _abc_44694_new_n4234_; 
wire _abc_44694_new_n4235_; 
wire _abc_44694_new_n4236_; 
wire _abc_44694_new_n4237_; 
wire _abc_44694_new_n4238_; 
wire _abc_44694_new_n4239_; 
wire _abc_44694_new_n4240_; 
wire _abc_44694_new_n4241_; 
wire _abc_44694_new_n4242_; 
wire _abc_44694_new_n4243_; 
wire _abc_44694_new_n4244_; 
wire _abc_44694_new_n4245_; 
wire _abc_44694_new_n4246_; 
wire _abc_44694_new_n4247_; 
wire _abc_44694_new_n4248_; 
wire _abc_44694_new_n4249_; 
wire _abc_44694_new_n4250_; 
wire _abc_44694_new_n4251_; 
wire _abc_44694_new_n4253_; 
wire _abc_44694_new_n4254_; 
wire _abc_44694_new_n4255_; 
wire _abc_44694_new_n4256_; 
wire _abc_44694_new_n4257_; 
wire _abc_44694_new_n4258_; 
wire _abc_44694_new_n4259_; 
wire _abc_44694_new_n4260_; 
wire _abc_44694_new_n4261_; 
wire _abc_44694_new_n4262_; 
wire _abc_44694_new_n4263_; 
wire _abc_44694_new_n4264_; 
wire _abc_44694_new_n4265_; 
wire _abc_44694_new_n4266_; 
wire _abc_44694_new_n4267_; 
wire _abc_44694_new_n4268_; 
wire _abc_44694_new_n4269_; 
wire _abc_44694_new_n4270_; 
wire _abc_44694_new_n4271_; 
wire _abc_44694_new_n4272_; 
wire _abc_44694_new_n4274_; 
wire _abc_44694_new_n4275_; 
wire _abc_44694_new_n4276_; 
wire _abc_44694_new_n4277_; 
wire _abc_44694_new_n4278_; 
wire _abc_44694_new_n4279_; 
wire _abc_44694_new_n4280_; 
wire _abc_44694_new_n4281_; 
wire _abc_44694_new_n4282_; 
wire _abc_44694_new_n4283_; 
wire _abc_44694_new_n4284_; 
wire _abc_44694_new_n4285_; 
wire _abc_44694_new_n4286_; 
wire _abc_44694_new_n4287_; 
wire _abc_44694_new_n4288_; 
wire _abc_44694_new_n4289_; 
wire _abc_44694_new_n4290_; 
wire _abc_44694_new_n4291_; 
wire _abc_44694_new_n4293_; 
wire _abc_44694_new_n4294_; 
wire _abc_44694_new_n4295_; 
wire _abc_44694_new_n4296_; 
wire _abc_44694_new_n4297_; 
wire _abc_44694_new_n4297__bF_buf0; 
wire _abc_44694_new_n4297__bF_buf1; 
wire _abc_44694_new_n4297__bF_buf2; 
wire _abc_44694_new_n4297__bF_buf3; 
wire _abc_44694_new_n4297__bF_buf4; 
wire _abc_44694_new_n4298_; 
wire _abc_44694_new_n4299_; 
wire _abc_44694_new_n4300_; 
wire _abc_44694_new_n4301_; 
wire _abc_44694_new_n4302_; 
wire _abc_44694_new_n4303_; 
wire _abc_44694_new_n4304_; 
wire _abc_44694_new_n4305_; 
wire _abc_44694_new_n4306_; 
wire _abc_44694_new_n4307_; 
wire _abc_44694_new_n4308_; 
wire _abc_44694_new_n4309_; 
wire _abc_44694_new_n4310_; 
wire _abc_44694_new_n4311_; 
wire _abc_44694_new_n4312_; 
wire _abc_44694_new_n4313_; 
wire _abc_44694_new_n4314_; 
wire _abc_44694_new_n4316_; 
wire _abc_44694_new_n4317_; 
wire _abc_44694_new_n4318_; 
wire _abc_44694_new_n4319_; 
wire _abc_44694_new_n4320_; 
wire _abc_44694_new_n4321_; 
wire _abc_44694_new_n4322_; 
wire _abc_44694_new_n4323_; 
wire _abc_44694_new_n4324_; 
wire _abc_44694_new_n4325_; 
wire _abc_44694_new_n4326_; 
wire _abc_44694_new_n4327_; 
wire _abc_44694_new_n4328_; 
wire _abc_44694_new_n4329_; 
wire _abc_44694_new_n4330_; 
wire _abc_44694_new_n4331_; 
wire _abc_44694_new_n4332_; 
wire _abc_44694_new_n4333_; 
wire _abc_44694_new_n4334_; 
wire _abc_44694_new_n4335_; 
wire _abc_44694_new_n4336_; 
wire _abc_44694_new_n4338_; 
wire _abc_44694_new_n4339_; 
wire _abc_44694_new_n4340_; 
wire _abc_44694_new_n4341_; 
wire _abc_44694_new_n4342_; 
wire _abc_44694_new_n4343_; 
wire _abc_44694_new_n4344_; 
wire _abc_44694_new_n4345_; 
wire _abc_44694_new_n4346_; 
wire _abc_44694_new_n4347_; 
wire _abc_44694_new_n4348_; 
wire _abc_44694_new_n4349_; 
wire _abc_44694_new_n4350_; 
wire _abc_44694_new_n4351_; 
wire _abc_44694_new_n4352_; 
wire _abc_44694_new_n4353_; 
wire _abc_44694_new_n4354_; 
wire _abc_44694_new_n4356_; 
wire _abc_44694_new_n4357_; 
wire _abc_44694_new_n4358_; 
wire _abc_44694_new_n4359_; 
wire _abc_44694_new_n4360_; 
wire _abc_44694_new_n4361_; 
wire _abc_44694_new_n4362_; 
wire _abc_44694_new_n4363_; 
wire _abc_44694_new_n4364_; 
wire _abc_44694_new_n4365_; 
wire _abc_44694_new_n4366_; 
wire _abc_44694_new_n4367_; 
wire _abc_44694_new_n4368_; 
wire _abc_44694_new_n4369_; 
wire _abc_44694_new_n4370_; 
wire _abc_44694_new_n4371_; 
wire _abc_44694_new_n4372_; 
wire _abc_44694_new_n4374_; 
wire _abc_44694_new_n4375_; 
wire _abc_44694_new_n4376_; 
wire _abc_44694_new_n4377_; 
wire _abc_44694_new_n4378_; 
wire _abc_44694_new_n4379_; 
wire _abc_44694_new_n4380_; 
wire _abc_44694_new_n4381_; 
wire _abc_44694_new_n4382_; 
wire _abc_44694_new_n4383_; 
wire _abc_44694_new_n4384_; 
wire _abc_44694_new_n4385_; 
wire _abc_44694_new_n4386_; 
wire _abc_44694_new_n4387_; 
wire _abc_44694_new_n4388_; 
wire _abc_44694_new_n4389_; 
wire _abc_44694_new_n4390_; 
wire _abc_44694_new_n4392_; 
wire _abc_44694_new_n4393_; 
wire _abc_44694_new_n4394_; 
wire _abc_44694_new_n4395_; 
wire _abc_44694_new_n4396_; 
wire _abc_44694_new_n4397_; 
wire _abc_44694_new_n4398_; 
wire _abc_44694_new_n4399_; 
wire _abc_44694_new_n4400_; 
wire _abc_44694_new_n4401_; 
wire _abc_44694_new_n4402_; 
wire _abc_44694_new_n4403_; 
wire _abc_44694_new_n4404_; 
wire _abc_44694_new_n4405_; 
wire _abc_44694_new_n4406_; 
wire _abc_44694_new_n4407_; 
wire _abc_44694_new_n4408_; 
wire _abc_44694_new_n4409_; 
wire _abc_44694_new_n4410_; 
wire _abc_44694_new_n4411_; 
wire _abc_44694_new_n4412_; 
wire _abc_44694_new_n4414_; 
wire _abc_44694_new_n4415_; 
wire _abc_44694_new_n4416_; 
wire _abc_44694_new_n4417_; 
wire _abc_44694_new_n4418_; 
wire _abc_44694_new_n4419_; 
wire _abc_44694_new_n4420_; 
wire _abc_44694_new_n4421_; 
wire _abc_44694_new_n4422_; 
wire _abc_44694_new_n4423_; 
wire _abc_44694_new_n4424_; 
wire _abc_44694_new_n4425_; 
wire _abc_44694_new_n4426_; 
wire _abc_44694_new_n4427_; 
wire _abc_44694_new_n4429_; 
wire _abc_44694_new_n4430_; 
wire _abc_44694_new_n4431_; 
wire _abc_44694_new_n4432_; 
wire _abc_44694_new_n4433_; 
wire _abc_44694_new_n4434_; 
wire _abc_44694_new_n4435_; 
wire _abc_44694_new_n4436_; 
wire _abc_44694_new_n4437_; 
wire _abc_44694_new_n4438_; 
wire _abc_44694_new_n4439_; 
wire _abc_44694_new_n4440_; 
wire _abc_44694_new_n4441_; 
wire _abc_44694_new_n4442_; 
wire _abc_44694_new_n4443_; 
wire _abc_44694_new_n4444_; 
wire _abc_44694_new_n4445_; 
wire _abc_44694_new_n4447_; 
wire _abc_44694_new_n4448_; 
wire _abc_44694_new_n4449_; 
wire _abc_44694_new_n4450_; 
wire _abc_44694_new_n4451_; 
wire _abc_44694_new_n4452_; 
wire _abc_44694_new_n4453_; 
wire _abc_44694_new_n4454_; 
wire _abc_44694_new_n4455_; 
wire _abc_44694_new_n4456_; 
wire _abc_44694_new_n4457_; 
wire _abc_44694_new_n4458_; 
wire _abc_44694_new_n4459_; 
wire _abc_44694_new_n4460_; 
wire _abc_44694_new_n4461_; 
wire _abc_44694_new_n4462_; 
wire _abc_44694_new_n4463_; 
wire _abc_44694_new_n4465_; 
wire _abc_44694_new_n4466_; 
wire _abc_44694_new_n4467_; 
wire _abc_44694_new_n4468_; 
wire _abc_44694_new_n4469_; 
wire _abc_44694_new_n4470_; 
wire _abc_44694_new_n4471_; 
wire _abc_44694_new_n4472_; 
wire _abc_44694_new_n4473_; 
wire _abc_44694_new_n4474_; 
wire _abc_44694_new_n4475_; 
wire _abc_44694_new_n4476_; 
wire _abc_44694_new_n4477_; 
wire _abc_44694_new_n4478_; 
wire _abc_44694_new_n4479_; 
wire _abc_44694_new_n4480_; 
wire _abc_44694_new_n4481_; 
wire _abc_44694_new_n4482_; 
wire _abc_44694_new_n4483_; 
wire _abc_44694_new_n4484_; 
wire _abc_44694_new_n4485_; 
wire _abc_44694_new_n4486_; 
wire _abc_44694_new_n4487_; 
wire _abc_44694_new_n4488_; 
wire _abc_44694_new_n4489_; 
wire _abc_44694_new_n4490_; 
wire _abc_44694_new_n4491_; 
wire _abc_44694_new_n4493_; 
wire _abc_44694_new_n4494_; 
wire _abc_44694_new_n4495_; 
wire _abc_44694_new_n4496_; 
wire _abc_44694_new_n4497_; 
wire _abc_44694_new_n4498_; 
wire _abc_44694_new_n4499_; 
wire _abc_44694_new_n4500_; 
wire _abc_44694_new_n4501_; 
wire _abc_44694_new_n4502_; 
wire _abc_44694_new_n4503_; 
wire _abc_44694_new_n4504_; 
wire _abc_44694_new_n4505_; 
wire _abc_44694_new_n4506_; 
wire _abc_44694_new_n4507_; 
wire _abc_44694_new_n4508_; 
wire _abc_44694_new_n4509_; 
wire _abc_44694_new_n4511_; 
wire _abc_44694_new_n4512_; 
wire _abc_44694_new_n4513_; 
wire _abc_44694_new_n4514_; 
wire _abc_44694_new_n4515_; 
wire _abc_44694_new_n4516_; 
wire _abc_44694_new_n4517_; 
wire _abc_44694_new_n4518_; 
wire _abc_44694_new_n4519_; 
wire _abc_44694_new_n4520_; 
wire _abc_44694_new_n4521_; 
wire _abc_44694_new_n4522_; 
wire _abc_44694_new_n4523_; 
wire _abc_44694_new_n4524_; 
wire _abc_44694_new_n4525_; 
wire _abc_44694_new_n4526_; 
wire _abc_44694_new_n4527_; 
wire _abc_44694_new_n4528_; 
wire _abc_44694_new_n4530_; 
wire _abc_44694_new_n4531_; 
wire _abc_44694_new_n4532_; 
wire _abc_44694_new_n4533_; 
wire _abc_44694_new_n4534_; 
wire _abc_44694_new_n4535_; 
wire _abc_44694_new_n4536_; 
wire _abc_44694_new_n4537_; 
wire _abc_44694_new_n4538_; 
wire _abc_44694_new_n4539_; 
wire _abc_44694_new_n4540_; 
wire _abc_44694_new_n4541_; 
wire _abc_44694_new_n4542_; 
wire _abc_44694_new_n4543_; 
wire _abc_44694_new_n4545_; 
wire _abc_44694_new_n4546_; 
wire _abc_44694_new_n4547_; 
wire _abc_44694_new_n4548_; 
wire _abc_44694_new_n4549_; 
wire _abc_44694_new_n4550_; 
wire _abc_44694_new_n4551_; 
wire _abc_44694_new_n4552_; 
wire _abc_44694_new_n4553_; 
wire _abc_44694_new_n4554_; 
wire _abc_44694_new_n4555_; 
wire _abc_44694_new_n4556_; 
wire _abc_44694_new_n4557_; 
wire _abc_44694_new_n4558_; 
wire _abc_44694_new_n4559_; 
wire _abc_44694_new_n4560_; 
wire _abc_44694_new_n4561_; 
wire _abc_44694_new_n4562_; 
wire _abc_44694_new_n4563_; 
wire _abc_44694_new_n4564_; 
wire _abc_44694_new_n4565_; 
wire _abc_44694_new_n4566_; 
wire _abc_44694_new_n4567_; 
wire _abc_44694_new_n4569_; 
wire _abc_44694_new_n4570_; 
wire _abc_44694_new_n4571_; 
wire _abc_44694_new_n4572_; 
wire _abc_44694_new_n4573_; 
wire _abc_44694_new_n4574_; 
wire _abc_44694_new_n4575_; 
wire _abc_44694_new_n4576_; 
wire _abc_44694_new_n4577_; 
wire _abc_44694_new_n4578_; 
wire _abc_44694_new_n4579_; 
wire _abc_44694_new_n4580_; 
wire _abc_44694_new_n4581_; 
wire _abc_44694_new_n4582_; 
wire _abc_44694_new_n4583_; 
wire _abc_44694_new_n4584_; 
wire _abc_44694_new_n4585_; 
wire _abc_44694_new_n4587_; 
wire _abc_44694_new_n4588_; 
wire _abc_44694_new_n4589_; 
wire _abc_44694_new_n4590_; 
wire _abc_44694_new_n4591_; 
wire _abc_44694_new_n4592_; 
wire _abc_44694_new_n4593_; 
wire _abc_44694_new_n4594_; 
wire _abc_44694_new_n4595_; 
wire _abc_44694_new_n4596_; 
wire _abc_44694_new_n4597_; 
wire _abc_44694_new_n4598_; 
wire _abc_44694_new_n4599_; 
wire _abc_44694_new_n4600_; 
wire _abc_44694_new_n4601_; 
wire _abc_44694_new_n4602_; 
wire _abc_44694_new_n4603_; 
wire _abc_44694_new_n4604_; 
wire _abc_44694_new_n4605_; 
wire _abc_44694_new_n4607_; 
wire _abc_44694_new_n4608_; 
wire _abc_44694_new_n4609_; 
wire _abc_44694_new_n4610_; 
wire _abc_44694_new_n4611_; 
wire _abc_44694_new_n4612_; 
wire _abc_44694_new_n4613_; 
wire _abc_44694_new_n4614_; 
wire _abc_44694_new_n4615_; 
wire _abc_44694_new_n4616_; 
wire _abc_44694_new_n4617_; 
wire _abc_44694_new_n4618_; 
wire _abc_44694_new_n4619_; 
wire _abc_44694_new_n4620_; 
wire _abc_44694_new_n4623_; 
wire _abc_44694_new_n4625_; 
wire _abc_44694_new_n4626_; 
wire _abc_44694_new_n617_; 
wire _abc_44694_new_n618_; 
wire _abc_44694_new_n619_; 
wire _abc_44694_new_n620_; 
wire _abc_44694_new_n621_; 
wire _abc_44694_new_n622_; 
wire _abc_44694_new_n623_; 
wire _abc_44694_new_n624_; 
wire _abc_44694_new_n625_; 
wire _abc_44694_new_n626_; 
wire _abc_44694_new_n627_; 
wire _abc_44694_new_n628_; 
wire _abc_44694_new_n630_; 
wire _abc_44694_new_n631_; 
wire _abc_44694_new_n632_; 
wire _abc_44694_new_n633_; 
wire _abc_44694_new_n634_; 
wire _abc_44694_new_n635_; 
wire _abc_44694_new_n636_; 
wire _abc_44694_new_n637_; 
wire _abc_44694_new_n638_; 
wire _abc_44694_new_n639_; 
wire _abc_44694_new_n640_; 
wire _abc_44694_new_n641_; 
wire _abc_44694_new_n642_; 
wire _abc_44694_new_n643_; 
wire _abc_44694_new_n644_; 
wire _abc_44694_new_n645_; 
wire _abc_44694_new_n646_; 
wire _abc_44694_new_n647_; 
wire _abc_44694_new_n648_; 
wire _abc_44694_new_n649_; 
wire _abc_44694_new_n650_; 
wire _abc_44694_new_n651_; 
wire _abc_44694_new_n652_; 
wire _abc_44694_new_n653_; 
wire _abc_44694_new_n654_; 
wire _abc_44694_new_n655_; 
wire _abc_44694_new_n656_; 
wire _abc_44694_new_n657_; 
wire _abc_44694_new_n658_; 
wire _abc_44694_new_n660_; 
wire _abc_44694_new_n661_; 
wire _abc_44694_new_n662_; 
wire _abc_44694_new_n664_; 
wire _abc_44694_new_n665_; 
wire _abc_44694_new_n667_; 
wire _abc_44694_new_n668_; 
wire _abc_44694_new_n668__bF_buf0; 
wire _abc_44694_new_n668__bF_buf1; 
wire _abc_44694_new_n668__bF_buf2; 
wire _abc_44694_new_n668__bF_buf3; 
wire _abc_44694_new_n668__bF_buf4; 
wire _abc_44694_new_n669_; 
wire _abc_44694_new_n671_; 
wire _abc_44694_new_n672_; 
wire _abc_44694_new_n673_; 
wire _abc_44694_new_n673__bF_buf0; 
wire _abc_44694_new_n673__bF_buf1; 
wire _abc_44694_new_n673__bF_buf2; 
wire _abc_44694_new_n673__bF_buf3; 
wire _abc_44694_new_n673__bF_buf4; 
wire _abc_44694_new_n674_; 
wire _abc_44694_new_n675_; 
wire _abc_44694_new_n676_; 
wire _abc_44694_new_n677_; 
wire _abc_44694_new_n677__bF_buf0; 
wire _abc_44694_new_n677__bF_buf1; 
wire _abc_44694_new_n677__bF_buf2; 
wire _abc_44694_new_n677__bF_buf3; 
wire _abc_44694_new_n678_; 
wire _abc_44694_new_n679_; 
wire _abc_44694_new_n680_; 
wire _abc_44694_new_n681_; 
wire _abc_44694_new_n682_; 
wire _abc_44694_new_n683_; 
wire _abc_44694_new_n684_; 
wire _abc_44694_new_n685_; 
wire _abc_44694_new_n686_; 
wire _abc_44694_new_n687_; 
wire _abc_44694_new_n688_; 
wire _abc_44694_new_n689_; 
wire _abc_44694_new_n690_; 
wire _abc_44694_new_n691_; 
wire _abc_44694_new_n692_; 
wire _abc_44694_new_n693_; 
wire _abc_44694_new_n694_; 
wire _abc_44694_new_n695_; 
wire _abc_44694_new_n696_; 
wire _abc_44694_new_n697_; 
wire _abc_44694_new_n699_; 
wire _abc_44694_new_n700_; 
wire _abc_44694_new_n701_; 
wire _abc_44694_new_n702_; 
wire _abc_44694_new_n703_; 
wire _abc_44694_new_n704_; 
wire _abc_44694_new_n705_; 
wire _abc_44694_new_n706_; 
wire _abc_44694_new_n707_; 
wire _abc_44694_new_n708_; 
wire _abc_44694_new_n709_; 
wire _abc_44694_new_n710_; 
wire _abc_44694_new_n711_; 
wire _abc_44694_new_n712_; 
wire _abc_44694_new_n713_; 
wire _abc_44694_new_n715_; 
wire _abc_44694_new_n716_; 
wire _abc_44694_new_n717_; 
wire _abc_44694_new_n718_; 
wire _abc_44694_new_n719_; 
wire _abc_44694_new_n720_; 
wire _abc_44694_new_n721_; 
wire _abc_44694_new_n722_; 
wire _abc_44694_new_n723_; 
wire _abc_44694_new_n724_; 
wire _abc_44694_new_n725_; 
wire _abc_44694_new_n726_; 
wire _abc_44694_new_n727_; 
wire _abc_44694_new_n728_; 
wire _abc_44694_new_n729_; 
wire _abc_44694_new_n731_; 
wire _abc_44694_new_n732_; 
wire _abc_44694_new_n733_; 
wire _abc_44694_new_n734_; 
wire _abc_44694_new_n735_; 
wire _abc_44694_new_n736_; 
wire _abc_44694_new_n737_; 
wire _abc_44694_new_n738_; 
wire _abc_44694_new_n739_; 
wire _abc_44694_new_n740_; 
wire _abc_44694_new_n741_; 
wire _abc_44694_new_n742_; 
wire _abc_44694_new_n743_; 
wire _abc_44694_new_n744_; 
wire _abc_44694_new_n745_; 
wire _abc_44694_new_n747_; 
wire _abc_44694_new_n748_; 
wire _abc_44694_new_n749_; 
wire _abc_44694_new_n750_; 
wire _abc_44694_new_n751_; 
wire _abc_44694_new_n752_; 
wire _abc_44694_new_n753_; 
wire _abc_44694_new_n754_; 
wire _abc_44694_new_n755_; 
wire _abc_44694_new_n756_; 
wire _abc_44694_new_n757_; 
wire _abc_44694_new_n758_; 
wire _abc_44694_new_n759_; 
wire _abc_44694_new_n760_; 
wire _abc_44694_new_n761_; 
wire _abc_44694_new_n763_; 
wire _abc_44694_new_n764_; 
wire _abc_44694_new_n765_; 
wire _abc_44694_new_n766_; 
wire _abc_44694_new_n767_; 
wire _abc_44694_new_n768_; 
wire _abc_44694_new_n769_; 
wire _abc_44694_new_n770_; 
wire _abc_44694_new_n771_; 
wire _abc_44694_new_n772_; 
wire _abc_44694_new_n773_; 
wire _abc_44694_new_n774_; 
wire _abc_44694_new_n775_; 
wire _abc_44694_new_n776_; 
wire _abc_44694_new_n777_; 
wire _abc_44694_new_n779_; 
wire _abc_44694_new_n780_; 
wire _abc_44694_new_n781_; 
wire _abc_44694_new_n782_; 
wire _abc_44694_new_n783_; 
wire _abc_44694_new_n784_; 
wire _abc_44694_new_n785_; 
wire _abc_44694_new_n786_; 
wire _abc_44694_new_n787_; 
wire _abc_44694_new_n788_; 
wire _abc_44694_new_n789_; 
wire _abc_44694_new_n790_; 
wire _abc_44694_new_n791_; 
wire _abc_44694_new_n792_; 
wire _abc_44694_new_n793_; 
wire _abc_44694_new_n795_; 
wire _abc_44694_new_n796_; 
wire _abc_44694_new_n797_; 
wire _abc_44694_new_n798_; 
wire _abc_44694_new_n799_; 
wire _abc_44694_new_n800_; 
wire _abc_44694_new_n801_; 
wire _abc_44694_new_n802_; 
wire _abc_44694_new_n803_; 
wire _abc_44694_new_n804_; 
wire _abc_44694_new_n805_; 
wire _abc_44694_new_n806_; 
wire _abc_44694_new_n807_; 
wire _abc_44694_new_n808_; 
wire _abc_44694_new_n809_; 
wire _abc_44694_new_n811_; 
wire _abc_44694_new_n812_; 
wire _abc_44694_new_n813_; 
wire _abc_44694_new_n814_; 
wire _abc_44694_new_n815_; 
wire _abc_44694_new_n816_; 
wire _abc_44694_new_n817_; 
wire _abc_44694_new_n817__bF_buf0; 
wire _abc_44694_new_n817__bF_buf1; 
wire _abc_44694_new_n817__bF_buf2; 
wire _abc_44694_new_n817__bF_buf3; 
wire _abc_44694_new_n818_; 
wire _abc_44694_new_n820_; 
wire _abc_44694_new_n821_; 
wire _abc_44694_new_n822_; 
wire _abc_44694_new_n823_; 
wire _abc_44694_new_n824_; 
wire _abc_44694_new_n825_; 
wire _abc_44694_new_n827_; 
wire _abc_44694_new_n828_; 
wire _abc_44694_new_n829_; 
wire _abc_44694_new_n830_; 
wire _abc_44694_new_n831_; 
wire _abc_44694_new_n832_; 
wire _abc_44694_new_n834_; 
wire _abc_44694_new_n835_; 
wire _abc_44694_new_n836_; 
wire _abc_44694_new_n837_; 
wire _abc_44694_new_n838_; 
wire _abc_44694_new_n839_; 
wire _abc_44694_new_n841_; 
wire _abc_44694_new_n842_; 
wire _abc_44694_new_n843_; 
wire _abc_44694_new_n844_; 
wire _abc_44694_new_n845_; 
wire _abc_44694_new_n846_; 
wire _abc_44694_new_n848_; 
wire _abc_44694_new_n849_; 
wire _abc_44694_new_n850_; 
wire _abc_44694_new_n851_; 
wire _abc_44694_new_n852_; 
wire _abc_44694_new_n853_; 
wire _abc_44694_new_n855_; 
wire _abc_44694_new_n856_; 
wire _abc_44694_new_n857_; 
wire _abc_44694_new_n858_; 
wire _abc_44694_new_n859_; 
wire _abc_44694_new_n860_; 
wire _abc_44694_new_n862_; 
wire _abc_44694_new_n863_; 
wire _abc_44694_new_n864_; 
wire _abc_44694_new_n865_; 
wire _abc_44694_new_n866_; 
wire _abc_44694_new_n867_; 
wire _abc_44694_new_n869_; 
wire _abc_44694_new_n870_; 
wire _abc_44694_new_n871_; 
wire _abc_44694_new_n872_; 
wire _abc_44694_new_n873_; 
wire _abc_44694_new_n874_; 
wire _abc_44694_new_n875_; 
wire _abc_44694_new_n876_; 
wire _abc_44694_new_n878_; 
wire _abc_44694_new_n879_; 
wire _abc_44694_new_n880_; 
wire _abc_44694_new_n881_; 
wire _abc_44694_new_n882_; 
wire _abc_44694_new_n884_; 
wire _abc_44694_new_n885_; 
wire _abc_44694_new_n886_; 
wire _abc_44694_new_n887_; 
wire _abc_44694_new_n888_; 
wire _abc_44694_new_n890_; 
wire _abc_44694_new_n891_; 
wire _abc_44694_new_n892_; 
wire _abc_44694_new_n893_; 
wire _abc_44694_new_n894_; 
wire _abc_44694_new_n896_; 
wire _abc_44694_new_n897_; 
wire _abc_44694_new_n898_; 
wire _abc_44694_new_n899_; 
wire _abc_44694_new_n900_; 
wire _abc_44694_new_n902_; 
wire _abc_44694_new_n903_; 
wire _abc_44694_new_n904_; 
wire _abc_44694_new_n905_; 
wire _abc_44694_new_n906_; 
wire _abc_44694_new_n908_; 
wire _abc_44694_new_n909_; 
wire _abc_44694_new_n910_; 
wire _abc_44694_new_n911_; 
wire _abc_44694_new_n912_; 
wire _abc_44694_new_n914_; 
wire _abc_44694_new_n915_; 
wire _abc_44694_new_n916_; 
wire _abc_44694_new_n917_; 
wire _abc_44694_new_n918_; 
wire _abc_44694_new_n920_; 
wire _abc_44694_new_n921_; 
wire _abc_44694_new_n922_; 
wire _abc_44694_new_n923_; 
wire _abc_44694_new_n924_; 
wire _abc_44694_new_n926_; 
wire _abc_44694_new_n927_; 
wire _abc_44694_new_n928_; 
wire _abc_44694_new_n929_; 
wire _abc_44694_new_n930_; 
wire _abc_44694_new_n932_; 
wire _abc_44694_new_n933_; 
wire _abc_44694_new_n934_; 
wire _abc_44694_new_n935_; 
wire _abc_44694_new_n936_; 
wire _abc_44694_new_n938_; 
wire _abc_44694_new_n939_; 
wire _abc_44694_new_n940_; 
wire _abc_44694_new_n941_; 
wire _abc_44694_new_n942_; 
wire _abc_44694_new_n944_; 
wire _abc_44694_new_n945_; 
wire _abc_44694_new_n946_; 
wire _abc_44694_new_n947_; 
wire _abc_44694_new_n948_; 
wire _abc_44694_new_n950_; 
wire _abc_44694_new_n951_; 
wire _abc_44694_new_n952_; 
wire _abc_44694_new_n953_; 
wire _abc_44694_new_n954_; 
wire _abc_44694_new_n956_; 
wire _abc_44694_new_n957_; 
wire _abc_44694_new_n958_; 
wire _abc_44694_new_n959_; 
wire _abc_44694_new_n960_; 
wire _abc_44694_new_n962_; 
wire _abc_44694_new_n963_; 
wire _abc_44694_new_n964_; 
wire _abc_44694_new_n965_; 
wire _abc_44694_new_n966_; 
wire _abc_44694_new_n969_; 
wire _abc_44694_new_n970_; 
wire _abc_44694_new_n971_; 
wire _abc_44694_new_n972_; 
wire _abc_44694_new_n973_; 
wire _abc_44694_new_n974_; 
wire _abc_44694_new_n975_; 
wire _abc_44694_new_n976_; 
wire _abc_44694_new_n977_; 
wire _abc_44694_new_n978_; 
wire _abc_44694_new_n979_; 
wire _abc_44694_new_n980_; 
wire _abc_44694_new_n981_; 
wire _abc_44694_new_n982_; 
wire _abc_44694_new_n983_; 
wire _abc_44694_new_n984_; 
wire _abc_44694_new_n985_; 
wire _abc_44694_new_n986_; 
wire _abc_44694_new_n987_; 
wire _abc_44694_new_n988_; 
wire _abc_44694_new_n989_; 
wire _abc_44694_new_n990_; 
wire _abc_44694_new_n991_; 
wire _abc_44694_new_n992_; 
wire _abc_44694_new_n993_; 
wire _abc_44694_new_n994_; 
wire _abc_44694_new_n995_; 
wire _abc_44694_new_n996_; 
wire _abc_44694_new_n997_; 
wire _abc_44694_new_n998_; 
wire _abc_44694_new_n999_; 
wire _auto_iopadmap_cc_368_execute_48707; 
wire _auto_iopadmap_cc_368_execute_48709; 
wire _auto_iopadmap_cc_368_execute_48711_0_; 
wire _auto_iopadmap_cc_368_execute_48711_10_; 
wire _auto_iopadmap_cc_368_execute_48711_11_; 
wire _auto_iopadmap_cc_368_execute_48711_12_; 
wire _auto_iopadmap_cc_368_execute_48711_13_; 
wire _auto_iopadmap_cc_368_execute_48711_14_; 
wire _auto_iopadmap_cc_368_execute_48711_15_; 
wire _auto_iopadmap_cc_368_execute_48711_16_; 
wire _auto_iopadmap_cc_368_execute_48711_17_; 
wire _auto_iopadmap_cc_368_execute_48711_18_; 
wire _auto_iopadmap_cc_368_execute_48711_19_; 
wire _auto_iopadmap_cc_368_execute_48711_1_; 
wire _auto_iopadmap_cc_368_execute_48711_20_; 
wire _auto_iopadmap_cc_368_execute_48711_21_; 
wire _auto_iopadmap_cc_368_execute_48711_22_; 
wire _auto_iopadmap_cc_368_execute_48711_23_; 
wire _auto_iopadmap_cc_368_execute_48711_24_; 
wire _auto_iopadmap_cc_368_execute_48711_25_; 
wire _auto_iopadmap_cc_368_execute_48711_26_; 
wire _auto_iopadmap_cc_368_execute_48711_27_; 
wire _auto_iopadmap_cc_368_execute_48711_28_; 
wire _auto_iopadmap_cc_368_execute_48711_29_; 
wire _auto_iopadmap_cc_368_execute_48711_2_; 
wire _auto_iopadmap_cc_368_execute_48711_30_; 
wire _auto_iopadmap_cc_368_execute_48711_31_; 
wire _auto_iopadmap_cc_368_execute_48711_3_; 
wire _auto_iopadmap_cc_368_execute_48711_4_; 
wire _auto_iopadmap_cc_368_execute_48711_5_; 
wire _auto_iopadmap_cc_368_execute_48711_6_; 
wire _auto_iopadmap_cc_368_execute_48711_7_; 
wire _auto_iopadmap_cc_368_execute_48711_8_; 
wire _auto_iopadmap_cc_368_execute_48711_9_; 
wire _auto_iopadmap_cc_368_execute_48748; 
wire _auto_iopadmap_cc_368_execute_48750_0_; 
wire _auto_iopadmap_cc_368_execute_48750_10_; 
wire _auto_iopadmap_cc_368_execute_48750_11_; 
wire _auto_iopadmap_cc_368_execute_48750_12_; 
wire _auto_iopadmap_cc_368_execute_48750_13_; 
wire _auto_iopadmap_cc_368_execute_48750_14_; 
wire _auto_iopadmap_cc_368_execute_48750_15_; 
wire _auto_iopadmap_cc_368_execute_48750_16_; 
wire _auto_iopadmap_cc_368_execute_48750_17_; 
wire _auto_iopadmap_cc_368_execute_48750_18_; 
wire _auto_iopadmap_cc_368_execute_48750_19_; 
wire _auto_iopadmap_cc_368_execute_48750_1_; 
wire _auto_iopadmap_cc_368_execute_48750_20_; 
wire _auto_iopadmap_cc_368_execute_48750_21_; 
wire _auto_iopadmap_cc_368_execute_48750_22_; 
wire _auto_iopadmap_cc_368_execute_48750_23_; 
wire _auto_iopadmap_cc_368_execute_48750_24_; 
wire _auto_iopadmap_cc_368_execute_48750_25_; 
wire _auto_iopadmap_cc_368_execute_48750_26_; 
wire _auto_iopadmap_cc_368_execute_48750_27_; 
wire _auto_iopadmap_cc_368_execute_48750_28_; 
wire _auto_iopadmap_cc_368_execute_48750_29_; 
wire _auto_iopadmap_cc_368_execute_48750_2_; 
wire _auto_iopadmap_cc_368_execute_48750_30_; 
wire _auto_iopadmap_cc_368_execute_48750_31_; 
wire _auto_iopadmap_cc_368_execute_48750_3_; 
wire _auto_iopadmap_cc_368_execute_48750_4_; 
wire _auto_iopadmap_cc_368_execute_48750_5_; 
wire _auto_iopadmap_cc_368_execute_48750_6_; 
wire _auto_iopadmap_cc_368_execute_48750_7_; 
wire _auto_iopadmap_cc_368_execute_48750_8_; 
wire _auto_iopadmap_cc_368_execute_48750_9_; 
wire _auto_iopadmap_cc_368_execute_48783_0_; 
wire _auto_iopadmap_cc_368_execute_48783_1_; 
wire _auto_iopadmap_cc_368_execute_48783_2_; 
wire _auto_iopadmap_cc_368_execute_48783_3_; 
wire _auto_iopadmap_cc_368_execute_48788; 
wire _auto_iopadmap_cc_368_execute_48790; 
wire alu__abc_42281_new_n1000_; 
wire alu__abc_42281_new_n1001_; 
wire alu__abc_42281_new_n1002_; 
wire alu__abc_42281_new_n1003_; 
wire alu__abc_42281_new_n1004_; 
wire alu__abc_42281_new_n1005_; 
wire alu__abc_42281_new_n1006_; 
wire alu__abc_42281_new_n1007_; 
wire alu__abc_42281_new_n1008_; 
wire alu__abc_42281_new_n1009_; 
wire alu__abc_42281_new_n1010_; 
wire alu__abc_42281_new_n1011_; 
wire alu__abc_42281_new_n1012_; 
wire alu__abc_42281_new_n1013_; 
wire alu__abc_42281_new_n1014_; 
wire alu__abc_42281_new_n1015_; 
wire alu__abc_42281_new_n1016_; 
wire alu__abc_42281_new_n1017_; 
wire alu__abc_42281_new_n1018_; 
wire alu__abc_42281_new_n1019_; 
wire alu__abc_42281_new_n1020_; 
wire alu__abc_42281_new_n1021_; 
wire alu__abc_42281_new_n1022_; 
wire alu__abc_42281_new_n1023_; 
wire alu__abc_42281_new_n1024_; 
wire alu__abc_42281_new_n1025_; 
wire alu__abc_42281_new_n1026_; 
wire alu__abc_42281_new_n1027_; 
wire alu__abc_42281_new_n1028_; 
wire alu__abc_42281_new_n1029_; 
wire alu__abc_42281_new_n1030_; 
wire alu__abc_42281_new_n1031_; 
wire alu__abc_42281_new_n1032_; 
wire alu__abc_42281_new_n1033_; 
wire alu__abc_42281_new_n1034_; 
wire alu__abc_42281_new_n1035_; 
wire alu__abc_42281_new_n1036_; 
wire alu__abc_42281_new_n1037_; 
wire alu__abc_42281_new_n1038_; 
wire alu__abc_42281_new_n1039_; 
wire alu__abc_42281_new_n1040_; 
wire alu__abc_42281_new_n1041_; 
wire alu__abc_42281_new_n1042_; 
wire alu__abc_42281_new_n1043_; 
wire alu__abc_42281_new_n1044_; 
wire alu__abc_42281_new_n1045_; 
wire alu__abc_42281_new_n1046_; 
wire alu__abc_42281_new_n1047_; 
wire alu__abc_42281_new_n1048_; 
wire alu__abc_42281_new_n1049_; 
wire alu__abc_42281_new_n1050_; 
wire alu__abc_42281_new_n1051_; 
wire alu__abc_42281_new_n1052_; 
wire alu__abc_42281_new_n1053_; 
wire alu__abc_42281_new_n1054_; 
wire alu__abc_42281_new_n1055_; 
wire alu__abc_42281_new_n1056_; 
wire alu__abc_42281_new_n1057_; 
wire alu__abc_42281_new_n1058_; 
wire alu__abc_42281_new_n1059_; 
wire alu__abc_42281_new_n1060_; 
wire alu__abc_42281_new_n1061_; 
wire alu__abc_42281_new_n1062_; 
wire alu__abc_42281_new_n1063_; 
wire alu__abc_42281_new_n1064_; 
wire alu__abc_42281_new_n1065_; 
wire alu__abc_42281_new_n1066_; 
wire alu__abc_42281_new_n1067_; 
wire alu__abc_42281_new_n1068_; 
wire alu__abc_42281_new_n1069_; 
wire alu__abc_42281_new_n1070_; 
wire alu__abc_42281_new_n1071_; 
wire alu__abc_42281_new_n1072_; 
wire alu__abc_42281_new_n1073_; 
wire alu__abc_42281_new_n1074_; 
wire alu__abc_42281_new_n1075_; 
wire alu__abc_42281_new_n1076_; 
wire alu__abc_42281_new_n1077_; 
wire alu__abc_42281_new_n1078_; 
wire alu__abc_42281_new_n1079_; 
wire alu__abc_42281_new_n1080_; 
wire alu__abc_42281_new_n1081_; 
wire alu__abc_42281_new_n1083_; 
wire alu__abc_42281_new_n1084_; 
wire alu__abc_42281_new_n1085_; 
wire alu__abc_42281_new_n1086_; 
wire alu__abc_42281_new_n1087_; 
wire alu__abc_42281_new_n1088_; 
wire alu__abc_42281_new_n1089_; 
wire alu__abc_42281_new_n1090_; 
wire alu__abc_42281_new_n1091_; 
wire alu__abc_42281_new_n1092_; 
wire alu__abc_42281_new_n1093_; 
wire alu__abc_42281_new_n1094_; 
wire alu__abc_42281_new_n1095_; 
wire alu__abc_42281_new_n1096_; 
wire alu__abc_42281_new_n1097_; 
wire alu__abc_42281_new_n1098_; 
wire alu__abc_42281_new_n1099_; 
wire alu__abc_42281_new_n1100_; 
wire alu__abc_42281_new_n1101_; 
wire alu__abc_42281_new_n1102_; 
wire alu__abc_42281_new_n1103_; 
wire alu__abc_42281_new_n1104_; 
wire alu__abc_42281_new_n1105_; 
wire alu__abc_42281_new_n1106_; 
wire alu__abc_42281_new_n1107_; 
wire alu__abc_42281_new_n1108_; 
wire alu__abc_42281_new_n1109_; 
wire alu__abc_42281_new_n110_; 
wire alu__abc_42281_new_n1110_; 
wire alu__abc_42281_new_n1111_; 
wire alu__abc_42281_new_n1112_; 
wire alu__abc_42281_new_n1113_; 
wire alu__abc_42281_new_n1114_; 
wire alu__abc_42281_new_n1115_; 
wire alu__abc_42281_new_n1116_; 
wire alu__abc_42281_new_n1117_; 
wire alu__abc_42281_new_n1118_; 
wire alu__abc_42281_new_n1119_; 
wire alu__abc_42281_new_n111_; 
wire alu__abc_42281_new_n1120_; 
wire alu__abc_42281_new_n1121_; 
wire alu__abc_42281_new_n1122_; 
wire alu__abc_42281_new_n1123_; 
wire alu__abc_42281_new_n1124_; 
wire alu__abc_42281_new_n1125_; 
wire alu__abc_42281_new_n1126_; 
wire alu__abc_42281_new_n1127_; 
wire alu__abc_42281_new_n1128_; 
wire alu__abc_42281_new_n1129_; 
wire alu__abc_42281_new_n112_; 
wire alu__abc_42281_new_n1130_; 
wire alu__abc_42281_new_n1131_; 
wire alu__abc_42281_new_n1132_; 
wire alu__abc_42281_new_n1133_; 
wire alu__abc_42281_new_n1134_; 
wire alu__abc_42281_new_n1135_; 
wire alu__abc_42281_new_n1136_; 
wire alu__abc_42281_new_n1137_; 
wire alu__abc_42281_new_n1138_; 
wire alu__abc_42281_new_n1139_; 
wire alu__abc_42281_new_n113_; 
wire alu__abc_42281_new_n1140_; 
wire alu__abc_42281_new_n1141_; 
wire alu__abc_42281_new_n1142_; 
wire alu__abc_42281_new_n1143_; 
wire alu__abc_42281_new_n1144_; 
wire alu__abc_42281_new_n1145_; 
wire alu__abc_42281_new_n1146_; 
wire alu__abc_42281_new_n1147_; 
wire alu__abc_42281_new_n1148_; 
wire alu__abc_42281_new_n1149_; 
wire alu__abc_42281_new_n114_; 
wire alu__abc_42281_new_n1150_; 
wire alu__abc_42281_new_n1151_; 
wire alu__abc_42281_new_n1152_; 
wire alu__abc_42281_new_n1153_; 
wire alu__abc_42281_new_n1154_; 
wire alu__abc_42281_new_n1155_; 
wire alu__abc_42281_new_n1156_; 
wire alu__abc_42281_new_n1157_; 
wire alu__abc_42281_new_n1159_; 
wire alu__abc_42281_new_n115_; 
wire alu__abc_42281_new_n1160_; 
wire alu__abc_42281_new_n1161_; 
wire alu__abc_42281_new_n1162_; 
wire alu__abc_42281_new_n1163_; 
wire alu__abc_42281_new_n1164_; 
wire alu__abc_42281_new_n1165_; 
wire alu__abc_42281_new_n1166_; 
wire alu__abc_42281_new_n1167_; 
wire alu__abc_42281_new_n1168_; 
wire alu__abc_42281_new_n1169_; 
wire alu__abc_42281_new_n116_; 
wire alu__abc_42281_new_n1170_; 
wire alu__abc_42281_new_n1171_; 
wire alu__abc_42281_new_n1172_; 
wire alu__abc_42281_new_n1173_; 
wire alu__abc_42281_new_n1174_; 
wire alu__abc_42281_new_n1175_; 
wire alu__abc_42281_new_n1176_; 
wire alu__abc_42281_new_n1177_; 
wire alu__abc_42281_new_n1178_; 
wire alu__abc_42281_new_n1179_; 
wire alu__abc_42281_new_n117_; 
wire alu__abc_42281_new_n1180_; 
wire alu__abc_42281_new_n1181_; 
wire alu__abc_42281_new_n1182_; 
wire alu__abc_42281_new_n1183_; 
wire alu__abc_42281_new_n1184_; 
wire alu__abc_42281_new_n1185_; 
wire alu__abc_42281_new_n1186_; 
wire alu__abc_42281_new_n1187_; 
wire alu__abc_42281_new_n1188_; 
wire alu__abc_42281_new_n1189_; 
wire alu__abc_42281_new_n118_; 
wire alu__abc_42281_new_n1190_; 
wire alu__abc_42281_new_n1191_; 
wire alu__abc_42281_new_n1192_; 
wire alu__abc_42281_new_n1193_; 
wire alu__abc_42281_new_n1194_; 
wire alu__abc_42281_new_n1195_; 
wire alu__abc_42281_new_n1196_; 
wire alu__abc_42281_new_n1197_; 
wire alu__abc_42281_new_n1198_; 
wire alu__abc_42281_new_n1199_; 
wire alu__abc_42281_new_n119_; 
wire alu__abc_42281_new_n1200_; 
wire alu__abc_42281_new_n1201_; 
wire alu__abc_42281_new_n1202_; 
wire alu__abc_42281_new_n1203_; 
wire alu__abc_42281_new_n1204_; 
wire alu__abc_42281_new_n1205_; 
wire alu__abc_42281_new_n1206_; 
wire alu__abc_42281_new_n1207_; 
wire alu__abc_42281_new_n1208_; 
wire alu__abc_42281_new_n1209_; 
wire alu__abc_42281_new_n120_; 
wire alu__abc_42281_new_n1210_; 
wire alu__abc_42281_new_n1211_; 
wire alu__abc_42281_new_n1212_; 
wire alu__abc_42281_new_n1213_; 
wire alu__abc_42281_new_n1214_; 
wire alu__abc_42281_new_n1215_; 
wire alu__abc_42281_new_n1216_; 
wire alu__abc_42281_new_n1217_; 
wire alu__abc_42281_new_n1218_; 
wire alu__abc_42281_new_n1219_; 
wire alu__abc_42281_new_n121_; 
wire alu__abc_42281_new_n1220_; 
wire alu__abc_42281_new_n1221_; 
wire alu__abc_42281_new_n1222_; 
wire alu__abc_42281_new_n1223_; 
wire alu__abc_42281_new_n1224_; 
wire alu__abc_42281_new_n1225_; 
wire alu__abc_42281_new_n1226_; 
wire alu__abc_42281_new_n1227_; 
wire alu__abc_42281_new_n1228_; 
wire alu__abc_42281_new_n1229_; 
wire alu__abc_42281_new_n122_; 
wire alu__abc_42281_new_n1230_; 
wire alu__abc_42281_new_n1231_; 
wire alu__abc_42281_new_n1233_; 
wire alu__abc_42281_new_n1234_; 
wire alu__abc_42281_new_n1235_; 
wire alu__abc_42281_new_n1236_; 
wire alu__abc_42281_new_n1237_; 
wire alu__abc_42281_new_n1238_; 
wire alu__abc_42281_new_n1239_; 
wire alu__abc_42281_new_n123_; 
wire alu__abc_42281_new_n1240_; 
wire alu__abc_42281_new_n1241_; 
wire alu__abc_42281_new_n1242_; 
wire alu__abc_42281_new_n1243_; 
wire alu__abc_42281_new_n1244_; 
wire alu__abc_42281_new_n1245_; 
wire alu__abc_42281_new_n1246_; 
wire alu__abc_42281_new_n1247_; 
wire alu__abc_42281_new_n1248_; 
wire alu__abc_42281_new_n1249_; 
wire alu__abc_42281_new_n124_; 
wire alu__abc_42281_new_n1250_; 
wire alu__abc_42281_new_n1251_; 
wire alu__abc_42281_new_n1252_; 
wire alu__abc_42281_new_n1253_; 
wire alu__abc_42281_new_n1254_; 
wire alu__abc_42281_new_n1255_; 
wire alu__abc_42281_new_n1256_; 
wire alu__abc_42281_new_n1257_; 
wire alu__abc_42281_new_n1258_; 
wire alu__abc_42281_new_n1259_; 
wire alu__abc_42281_new_n125_; 
wire alu__abc_42281_new_n1260_; 
wire alu__abc_42281_new_n1261_; 
wire alu__abc_42281_new_n1262_; 
wire alu__abc_42281_new_n1263_; 
wire alu__abc_42281_new_n1264_; 
wire alu__abc_42281_new_n1265_; 
wire alu__abc_42281_new_n1266_; 
wire alu__abc_42281_new_n1267_; 
wire alu__abc_42281_new_n1268_; 
wire alu__abc_42281_new_n1269_; 
wire alu__abc_42281_new_n126_; 
wire alu__abc_42281_new_n1270_; 
wire alu__abc_42281_new_n1271_; 
wire alu__abc_42281_new_n1272_; 
wire alu__abc_42281_new_n1273_; 
wire alu__abc_42281_new_n1274_; 
wire alu__abc_42281_new_n1275_; 
wire alu__abc_42281_new_n1276_; 
wire alu__abc_42281_new_n1277_; 
wire alu__abc_42281_new_n1278_; 
wire alu__abc_42281_new_n1279_; 
wire alu__abc_42281_new_n127_; 
wire alu__abc_42281_new_n1280_; 
wire alu__abc_42281_new_n1281_; 
wire alu__abc_42281_new_n1282_; 
wire alu__abc_42281_new_n1283_; 
wire alu__abc_42281_new_n1285_; 
wire alu__abc_42281_new_n1286_; 
wire alu__abc_42281_new_n1287_; 
wire alu__abc_42281_new_n1288_; 
wire alu__abc_42281_new_n1289_; 
wire alu__abc_42281_new_n128_; 
wire alu__abc_42281_new_n1290_; 
wire alu__abc_42281_new_n1291_; 
wire alu__abc_42281_new_n1292_; 
wire alu__abc_42281_new_n1293_; 
wire alu__abc_42281_new_n1294_; 
wire alu__abc_42281_new_n1295_; 
wire alu__abc_42281_new_n1296_; 
wire alu__abc_42281_new_n1297_; 
wire alu__abc_42281_new_n1298_; 
wire alu__abc_42281_new_n1299_; 
wire alu__abc_42281_new_n129_; 
wire alu__abc_42281_new_n1300_; 
wire alu__abc_42281_new_n1301_; 
wire alu__abc_42281_new_n1302_; 
wire alu__abc_42281_new_n1303_; 
wire alu__abc_42281_new_n1304_; 
wire alu__abc_42281_new_n1305_; 
wire alu__abc_42281_new_n1306_; 
wire alu__abc_42281_new_n1307_; 
wire alu__abc_42281_new_n1308_; 
wire alu__abc_42281_new_n1309_; 
wire alu__abc_42281_new_n130_; 
wire alu__abc_42281_new_n1310_; 
wire alu__abc_42281_new_n1311_; 
wire alu__abc_42281_new_n1312_; 
wire alu__abc_42281_new_n1313_; 
wire alu__abc_42281_new_n1314_; 
wire alu__abc_42281_new_n1315_; 
wire alu__abc_42281_new_n1316_; 
wire alu__abc_42281_new_n1317_; 
wire alu__abc_42281_new_n1318_; 
wire alu__abc_42281_new_n1319_; 
wire alu__abc_42281_new_n131_; 
wire alu__abc_42281_new_n1320_; 
wire alu__abc_42281_new_n1321_; 
wire alu__abc_42281_new_n1322_; 
wire alu__abc_42281_new_n1323_; 
wire alu__abc_42281_new_n1324_; 
wire alu__abc_42281_new_n1325_; 
wire alu__abc_42281_new_n1326_; 
wire alu__abc_42281_new_n1327_; 
wire alu__abc_42281_new_n1328_; 
wire alu__abc_42281_new_n1329_; 
wire alu__abc_42281_new_n132_; 
wire alu__abc_42281_new_n1330_; 
wire alu__abc_42281_new_n1331_; 
wire alu__abc_42281_new_n1332_; 
wire alu__abc_42281_new_n1333_; 
wire alu__abc_42281_new_n1334_; 
wire alu__abc_42281_new_n1335_; 
wire alu__abc_42281_new_n1337_; 
wire alu__abc_42281_new_n1338_; 
wire alu__abc_42281_new_n1339_; 
wire alu__abc_42281_new_n133_; 
wire alu__abc_42281_new_n1340_; 
wire alu__abc_42281_new_n1341_; 
wire alu__abc_42281_new_n1342_; 
wire alu__abc_42281_new_n1343_; 
wire alu__abc_42281_new_n1344_; 
wire alu__abc_42281_new_n1345_; 
wire alu__abc_42281_new_n1346_; 
wire alu__abc_42281_new_n1347_; 
wire alu__abc_42281_new_n1348_; 
wire alu__abc_42281_new_n1349_; 
wire alu__abc_42281_new_n134_; 
wire alu__abc_42281_new_n1350_; 
wire alu__abc_42281_new_n1351_; 
wire alu__abc_42281_new_n1352_; 
wire alu__abc_42281_new_n1353_; 
wire alu__abc_42281_new_n1354_; 
wire alu__abc_42281_new_n1355_; 
wire alu__abc_42281_new_n1356_; 
wire alu__abc_42281_new_n1357_; 
wire alu__abc_42281_new_n1358_; 
wire alu__abc_42281_new_n1359_; 
wire alu__abc_42281_new_n135_; 
wire alu__abc_42281_new_n1360_; 
wire alu__abc_42281_new_n1361_; 
wire alu__abc_42281_new_n1362_; 
wire alu__abc_42281_new_n1363_; 
wire alu__abc_42281_new_n1364_; 
wire alu__abc_42281_new_n1365_; 
wire alu__abc_42281_new_n1366_; 
wire alu__abc_42281_new_n1367_; 
wire alu__abc_42281_new_n1368_; 
wire alu__abc_42281_new_n1369_; 
wire alu__abc_42281_new_n136_; 
wire alu__abc_42281_new_n1370_; 
wire alu__abc_42281_new_n1371_; 
wire alu__abc_42281_new_n1372_; 
wire alu__abc_42281_new_n1373_; 
wire alu__abc_42281_new_n1374_; 
wire alu__abc_42281_new_n1375_; 
wire alu__abc_42281_new_n1376_; 
wire alu__abc_42281_new_n1377_; 
wire alu__abc_42281_new_n1378_; 
wire alu__abc_42281_new_n1379_; 
wire alu__abc_42281_new_n137_; 
wire alu__abc_42281_new_n1380_; 
wire alu__abc_42281_new_n1381_; 
wire alu__abc_42281_new_n1382_; 
wire alu__abc_42281_new_n1383_; 
wire alu__abc_42281_new_n1384_; 
wire alu__abc_42281_new_n1385_; 
wire alu__abc_42281_new_n1386_; 
wire alu__abc_42281_new_n1388_; 
wire alu__abc_42281_new_n1389_; 
wire alu__abc_42281_new_n138_; 
wire alu__abc_42281_new_n1390_; 
wire alu__abc_42281_new_n1391_; 
wire alu__abc_42281_new_n1392_; 
wire alu__abc_42281_new_n1393_; 
wire alu__abc_42281_new_n1394_; 
wire alu__abc_42281_new_n1395_; 
wire alu__abc_42281_new_n1396_; 
wire alu__abc_42281_new_n1397_; 
wire alu__abc_42281_new_n1398_; 
wire alu__abc_42281_new_n1399_; 
wire alu__abc_42281_new_n139_; 
wire alu__abc_42281_new_n1400_; 
wire alu__abc_42281_new_n1401_; 
wire alu__abc_42281_new_n1402_; 
wire alu__abc_42281_new_n1403_; 
wire alu__abc_42281_new_n1404_; 
wire alu__abc_42281_new_n1405_; 
wire alu__abc_42281_new_n1406_; 
wire alu__abc_42281_new_n1407_; 
wire alu__abc_42281_new_n1408_; 
wire alu__abc_42281_new_n1409_; 
wire alu__abc_42281_new_n140_; 
wire alu__abc_42281_new_n1410_; 
wire alu__abc_42281_new_n1411_; 
wire alu__abc_42281_new_n1412_; 
wire alu__abc_42281_new_n1413_; 
wire alu__abc_42281_new_n1414_; 
wire alu__abc_42281_new_n1415_; 
wire alu__abc_42281_new_n1416_; 
wire alu__abc_42281_new_n1417_; 
wire alu__abc_42281_new_n1418_; 
wire alu__abc_42281_new_n1419_; 
wire alu__abc_42281_new_n141_; 
wire alu__abc_42281_new_n1420_; 
wire alu__abc_42281_new_n1421_; 
wire alu__abc_42281_new_n1422_; 
wire alu__abc_42281_new_n1423_; 
wire alu__abc_42281_new_n1424_; 
wire alu__abc_42281_new_n1425_; 
wire alu__abc_42281_new_n1426_; 
wire alu__abc_42281_new_n1427_; 
wire alu__abc_42281_new_n1428_; 
wire alu__abc_42281_new_n1429_; 
wire alu__abc_42281_new_n142_; 
wire alu__abc_42281_new_n1430_; 
wire alu__abc_42281_new_n1431_; 
wire alu__abc_42281_new_n1432_; 
wire alu__abc_42281_new_n1433_; 
wire alu__abc_42281_new_n1434_; 
wire alu__abc_42281_new_n1435_; 
wire alu__abc_42281_new_n1436_; 
wire alu__abc_42281_new_n1437_; 
wire alu__abc_42281_new_n1438_; 
wire alu__abc_42281_new_n143_; 
wire alu__abc_42281_new_n1440_; 
wire alu__abc_42281_new_n1441_; 
wire alu__abc_42281_new_n1442_; 
wire alu__abc_42281_new_n1443_; 
wire alu__abc_42281_new_n1444_; 
wire alu__abc_42281_new_n1445_; 
wire alu__abc_42281_new_n1446_; 
wire alu__abc_42281_new_n1447_; 
wire alu__abc_42281_new_n1448_; 
wire alu__abc_42281_new_n1449_; 
wire alu__abc_42281_new_n144_; 
wire alu__abc_42281_new_n1450_; 
wire alu__abc_42281_new_n1451_; 
wire alu__abc_42281_new_n1452_; 
wire alu__abc_42281_new_n1453_; 
wire alu__abc_42281_new_n1454_; 
wire alu__abc_42281_new_n1455_; 
wire alu__abc_42281_new_n1456_; 
wire alu__abc_42281_new_n1457_; 
wire alu__abc_42281_new_n1458_; 
wire alu__abc_42281_new_n1459_; 
wire alu__abc_42281_new_n145_; 
wire alu__abc_42281_new_n1460_; 
wire alu__abc_42281_new_n1461_; 
wire alu__abc_42281_new_n1462_; 
wire alu__abc_42281_new_n1463_; 
wire alu__abc_42281_new_n1464_; 
wire alu__abc_42281_new_n1465_; 
wire alu__abc_42281_new_n1466_; 
wire alu__abc_42281_new_n1467_; 
wire alu__abc_42281_new_n1468_; 
wire alu__abc_42281_new_n1469_; 
wire alu__abc_42281_new_n146_; 
wire alu__abc_42281_new_n1470_; 
wire alu__abc_42281_new_n1471_; 
wire alu__abc_42281_new_n1472_; 
wire alu__abc_42281_new_n1473_; 
wire alu__abc_42281_new_n1474_; 
wire alu__abc_42281_new_n1475_; 
wire alu__abc_42281_new_n1476_; 
wire alu__abc_42281_new_n1477_; 
wire alu__abc_42281_new_n1478_; 
wire alu__abc_42281_new_n1479_; 
wire alu__abc_42281_new_n147_; 
wire alu__abc_42281_new_n1480_; 
wire alu__abc_42281_new_n1481_; 
wire alu__abc_42281_new_n1483_; 
wire alu__abc_42281_new_n1484_; 
wire alu__abc_42281_new_n1485_; 
wire alu__abc_42281_new_n1486_; 
wire alu__abc_42281_new_n1487_; 
wire alu__abc_42281_new_n1488_; 
wire alu__abc_42281_new_n1489_; 
wire alu__abc_42281_new_n148_; 
wire alu__abc_42281_new_n1490_; 
wire alu__abc_42281_new_n1491_; 
wire alu__abc_42281_new_n1492_; 
wire alu__abc_42281_new_n1493_; 
wire alu__abc_42281_new_n1494_; 
wire alu__abc_42281_new_n1495_; 
wire alu__abc_42281_new_n1496_; 
wire alu__abc_42281_new_n1497_; 
wire alu__abc_42281_new_n1498_; 
wire alu__abc_42281_new_n1499_; 
wire alu__abc_42281_new_n149_; 
wire alu__abc_42281_new_n1500_; 
wire alu__abc_42281_new_n1501_; 
wire alu__abc_42281_new_n1502_; 
wire alu__abc_42281_new_n1503_; 
wire alu__abc_42281_new_n1504_; 
wire alu__abc_42281_new_n1505_; 
wire alu__abc_42281_new_n1506_; 
wire alu__abc_42281_new_n1507_; 
wire alu__abc_42281_new_n1508_; 
wire alu__abc_42281_new_n1509_; 
wire alu__abc_42281_new_n150_; 
wire alu__abc_42281_new_n1510_; 
wire alu__abc_42281_new_n1511_; 
wire alu__abc_42281_new_n1512_; 
wire alu__abc_42281_new_n1513_; 
wire alu__abc_42281_new_n1514_; 
wire alu__abc_42281_new_n1515_; 
wire alu__abc_42281_new_n1516_; 
wire alu__abc_42281_new_n1517_; 
wire alu__abc_42281_new_n1518_; 
wire alu__abc_42281_new_n1519_; 
wire alu__abc_42281_new_n151_; 
wire alu__abc_42281_new_n1520_; 
wire alu__abc_42281_new_n1521_; 
wire alu__abc_42281_new_n1522_; 
wire alu__abc_42281_new_n1523_; 
wire alu__abc_42281_new_n1524_; 
wire alu__abc_42281_new_n1526_; 
wire alu__abc_42281_new_n1527_; 
wire alu__abc_42281_new_n1528_; 
wire alu__abc_42281_new_n1529_; 
wire alu__abc_42281_new_n152_; 
wire alu__abc_42281_new_n1530_; 
wire alu__abc_42281_new_n1531_; 
wire alu__abc_42281_new_n1532_; 
wire alu__abc_42281_new_n1533_; 
wire alu__abc_42281_new_n1534_; 
wire alu__abc_42281_new_n1535_; 
wire alu__abc_42281_new_n1536_; 
wire alu__abc_42281_new_n1537_; 
wire alu__abc_42281_new_n1538_; 
wire alu__abc_42281_new_n1539_; 
wire alu__abc_42281_new_n153_; 
wire alu__abc_42281_new_n1540_; 
wire alu__abc_42281_new_n1541_; 
wire alu__abc_42281_new_n1542_; 
wire alu__abc_42281_new_n1543_; 
wire alu__abc_42281_new_n1544_; 
wire alu__abc_42281_new_n1545_; 
wire alu__abc_42281_new_n1546_; 
wire alu__abc_42281_new_n1547_; 
wire alu__abc_42281_new_n1548_; 
wire alu__abc_42281_new_n1549_; 
wire alu__abc_42281_new_n154_; 
wire alu__abc_42281_new_n1550_; 
wire alu__abc_42281_new_n1551_; 
wire alu__abc_42281_new_n1552_; 
wire alu__abc_42281_new_n1553_; 
wire alu__abc_42281_new_n1554_; 
wire alu__abc_42281_new_n1555_; 
wire alu__abc_42281_new_n1556_; 
wire alu__abc_42281_new_n1557_; 
wire alu__abc_42281_new_n1558_; 
wire alu__abc_42281_new_n1559_; 
wire alu__abc_42281_new_n155_; 
wire alu__abc_42281_new_n1560_; 
wire alu__abc_42281_new_n1561_; 
wire alu__abc_42281_new_n1562_; 
wire alu__abc_42281_new_n1563_; 
wire alu__abc_42281_new_n1564_; 
wire alu__abc_42281_new_n1565_; 
wire alu__abc_42281_new_n1566_; 
wire alu__abc_42281_new_n1567_; 
wire alu__abc_42281_new_n1568_; 
wire alu__abc_42281_new_n1569_; 
wire alu__abc_42281_new_n156_; 
wire alu__abc_42281_new_n1571_; 
wire alu__abc_42281_new_n1572_; 
wire alu__abc_42281_new_n1573_; 
wire alu__abc_42281_new_n1574_; 
wire alu__abc_42281_new_n1575_; 
wire alu__abc_42281_new_n1576_; 
wire alu__abc_42281_new_n1577_; 
wire alu__abc_42281_new_n1578_; 
wire alu__abc_42281_new_n1579_; 
wire alu__abc_42281_new_n157_; 
wire alu__abc_42281_new_n1580_; 
wire alu__abc_42281_new_n1581_; 
wire alu__abc_42281_new_n1582_; 
wire alu__abc_42281_new_n1583_; 
wire alu__abc_42281_new_n1584_; 
wire alu__abc_42281_new_n1585_; 
wire alu__abc_42281_new_n1586_; 
wire alu__abc_42281_new_n1587_; 
wire alu__abc_42281_new_n1588_; 
wire alu__abc_42281_new_n1589_; 
wire alu__abc_42281_new_n158_; 
wire alu__abc_42281_new_n1590_; 
wire alu__abc_42281_new_n1591_; 
wire alu__abc_42281_new_n1592_; 
wire alu__abc_42281_new_n1593_; 
wire alu__abc_42281_new_n1594_; 
wire alu__abc_42281_new_n1595_; 
wire alu__abc_42281_new_n1596_; 
wire alu__abc_42281_new_n1597_; 
wire alu__abc_42281_new_n1598_; 
wire alu__abc_42281_new_n1599_; 
wire alu__abc_42281_new_n159_; 
wire alu__abc_42281_new_n1600_; 
wire alu__abc_42281_new_n1601_; 
wire alu__abc_42281_new_n1602_; 
wire alu__abc_42281_new_n1603_; 
wire alu__abc_42281_new_n1604_; 
wire alu__abc_42281_new_n1605_; 
wire alu__abc_42281_new_n1606_; 
wire alu__abc_42281_new_n1607_; 
wire alu__abc_42281_new_n1608_; 
wire alu__abc_42281_new_n1609_; 
wire alu__abc_42281_new_n160_; 
wire alu__abc_42281_new_n1610_; 
wire alu__abc_42281_new_n1611_; 
wire alu__abc_42281_new_n1612_; 
wire alu__abc_42281_new_n1613_; 
wire alu__abc_42281_new_n1615_; 
wire alu__abc_42281_new_n1616_; 
wire alu__abc_42281_new_n1617_; 
wire alu__abc_42281_new_n1618_; 
wire alu__abc_42281_new_n1619_; 
wire alu__abc_42281_new_n161_; 
wire alu__abc_42281_new_n1620_; 
wire alu__abc_42281_new_n1621_; 
wire alu__abc_42281_new_n1622_; 
wire alu__abc_42281_new_n1623_; 
wire alu__abc_42281_new_n1624_; 
wire alu__abc_42281_new_n1625_; 
wire alu__abc_42281_new_n1626_; 
wire alu__abc_42281_new_n1627_; 
wire alu__abc_42281_new_n1628_; 
wire alu__abc_42281_new_n1629_; 
wire alu__abc_42281_new_n162_; 
wire alu__abc_42281_new_n1630_; 
wire alu__abc_42281_new_n1631_; 
wire alu__abc_42281_new_n1632_; 
wire alu__abc_42281_new_n1633_; 
wire alu__abc_42281_new_n1634_; 
wire alu__abc_42281_new_n1635_; 
wire alu__abc_42281_new_n1636_; 
wire alu__abc_42281_new_n1637_; 
wire alu__abc_42281_new_n1638_; 
wire alu__abc_42281_new_n1639_; 
wire alu__abc_42281_new_n163_; 
wire alu__abc_42281_new_n1640_; 
wire alu__abc_42281_new_n1641_; 
wire alu__abc_42281_new_n1642_; 
wire alu__abc_42281_new_n1643_; 
wire alu__abc_42281_new_n1644_; 
wire alu__abc_42281_new_n1645_; 
wire alu__abc_42281_new_n1646_; 
wire alu__abc_42281_new_n1647_; 
wire alu__abc_42281_new_n1648_; 
wire alu__abc_42281_new_n1649_; 
wire alu__abc_42281_new_n164_; 
wire alu__abc_42281_new_n1650_; 
wire alu__abc_42281_new_n1651_; 
wire alu__abc_42281_new_n1652_; 
wire alu__abc_42281_new_n1653_; 
wire alu__abc_42281_new_n1654_; 
wire alu__abc_42281_new_n1655_; 
wire alu__abc_42281_new_n1656_; 
wire alu__abc_42281_new_n1657_; 
wire alu__abc_42281_new_n1658_; 
wire alu__abc_42281_new_n165_; 
wire alu__abc_42281_new_n1660_; 
wire alu__abc_42281_new_n1661_; 
wire alu__abc_42281_new_n1662_; 
wire alu__abc_42281_new_n1663_; 
wire alu__abc_42281_new_n1664_; 
wire alu__abc_42281_new_n1665_; 
wire alu__abc_42281_new_n1666_; 
wire alu__abc_42281_new_n1667_; 
wire alu__abc_42281_new_n1668_; 
wire alu__abc_42281_new_n1669_; 
wire alu__abc_42281_new_n166_; 
wire alu__abc_42281_new_n1670_; 
wire alu__abc_42281_new_n1671_; 
wire alu__abc_42281_new_n1672_; 
wire alu__abc_42281_new_n1673_; 
wire alu__abc_42281_new_n1674_; 
wire alu__abc_42281_new_n1675_; 
wire alu__abc_42281_new_n1676_; 
wire alu__abc_42281_new_n1677_; 
wire alu__abc_42281_new_n1678_; 
wire alu__abc_42281_new_n1679_; 
wire alu__abc_42281_new_n167_; 
wire alu__abc_42281_new_n1680_; 
wire alu__abc_42281_new_n1681_; 
wire alu__abc_42281_new_n1682_; 
wire alu__abc_42281_new_n1683_; 
wire alu__abc_42281_new_n1684_; 
wire alu__abc_42281_new_n1685_; 
wire alu__abc_42281_new_n1686_; 
wire alu__abc_42281_new_n1687_; 
wire alu__abc_42281_new_n1688_; 
wire alu__abc_42281_new_n1689_; 
wire alu__abc_42281_new_n168_; 
wire alu__abc_42281_new_n1690_; 
wire alu__abc_42281_new_n1691_; 
wire alu__abc_42281_new_n1692_; 
wire alu__abc_42281_new_n1693_; 
wire alu__abc_42281_new_n1694_; 
wire alu__abc_42281_new_n1695_; 
wire alu__abc_42281_new_n1696_; 
wire alu__abc_42281_new_n1697_; 
wire alu__abc_42281_new_n1698_; 
wire alu__abc_42281_new_n1699_; 
wire alu__abc_42281_new_n169_; 
wire alu__abc_42281_new_n1700_; 
wire alu__abc_42281_new_n1701_; 
wire alu__abc_42281_new_n1702_; 
wire alu__abc_42281_new_n1704_; 
wire alu__abc_42281_new_n1705_; 
wire alu__abc_42281_new_n1706_; 
wire alu__abc_42281_new_n1707_; 
wire alu__abc_42281_new_n1708_; 
wire alu__abc_42281_new_n1709_; 
wire alu__abc_42281_new_n170_; 
wire alu__abc_42281_new_n1710_; 
wire alu__abc_42281_new_n1711_; 
wire alu__abc_42281_new_n1712_; 
wire alu__abc_42281_new_n1713_; 
wire alu__abc_42281_new_n1714_; 
wire alu__abc_42281_new_n1715_; 
wire alu__abc_42281_new_n1716_; 
wire alu__abc_42281_new_n1717_; 
wire alu__abc_42281_new_n1718_; 
wire alu__abc_42281_new_n1719_; 
wire alu__abc_42281_new_n171_; 
wire alu__abc_42281_new_n1720_; 
wire alu__abc_42281_new_n1721_; 
wire alu__abc_42281_new_n1722_; 
wire alu__abc_42281_new_n1723_; 
wire alu__abc_42281_new_n1724_; 
wire alu__abc_42281_new_n1725_; 
wire alu__abc_42281_new_n1726_; 
wire alu__abc_42281_new_n1727_; 
wire alu__abc_42281_new_n1728_; 
wire alu__abc_42281_new_n1729_; 
wire alu__abc_42281_new_n172_; 
wire alu__abc_42281_new_n1730_; 
wire alu__abc_42281_new_n1731_; 
wire alu__abc_42281_new_n1732_; 
wire alu__abc_42281_new_n1733_; 
wire alu__abc_42281_new_n1734_; 
wire alu__abc_42281_new_n1735_; 
wire alu__abc_42281_new_n1736_; 
wire alu__abc_42281_new_n1737_; 
wire alu__abc_42281_new_n1738_; 
wire alu__abc_42281_new_n1739_; 
wire alu__abc_42281_new_n173_; 
wire alu__abc_42281_new_n1740_; 
wire alu__abc_42281_new_n1741_; 
wire alu__abc_42281_new_n1742_; 
wire alu__abc_42281_new_n1743_; 
wire alu__abc_42281_new_n1744_; 
wire alu__abc_42281_new_n1745_; 
wire alu__abc_42281_new_n1746_; 
wire alu__abc_42281_new_n1747_; 
wire alu__abc_42281_new_n1749_; 
wire alu__abc_42281_new_n174_; 
wire alu__abc_42281_new_n1750_; 
wire alu__abc_42281_new_n1751_; 
wire alu__abc_42281_new_n1752_; 
wire alu__abc_42281_new_n1753_; 
wire alu__abc_42281_new_n1754_; 
wire alu__abc_42281_new_n1755_; 
wire alu__abc_42281_new_n1756_; 
wire alu__abc_42281_new_n1757_; 
wire alu__abc_42281_new_n1758_; 
wire alu__abc_42281_new_n1759_; 
wire alu__abc_42281_new_n175_; 
wire alu__abc_42281_new_n1760_; 
wire alu__abc_42281_new_n1761_; 
wire alu__abc_42281_new_n1762_; 
wire alu__abc_42281_new_n1763_; 
wire alu__abc_42281_new_n1764_; 
wire alu__abc_42281_new_n1765_; 
wire alu__abc_42281_new_n1766_; 
wire alu__abc_42281_new_n1767_; 
wire alu__abc_42281_new_n1768_; 
wire alu__abc_42281_new_n1769_; 
wire alu__abc_42281_new_n176_; 
wire alu__abc_42281_new_n1770_; 
wire alu__abc_42281_new_n1771_; 
wire alu__abc_42281_new_n1772_; 
wire alu__abc_42281_new_n1773_; 
wire alu__abc_42281_new_n1774_; 
wire alu__abc_42281_new_n1775_; 
wire alu__abc_42281_new_n1776_; 
wire alu__abc_42281_new_n1777_; 
wire alu__abc_42281_new_n1778_; 
wire alu__abc_42281_new_n1779_; 
wire alu__abc_42281_new_n177_; 
wire alu__abc_42281_new_n1780_; 
wire alu__abc_42281_new_n1781_; 
wire alu__abc_42281_new_n1782_; 
wire alu__abc_42281_new_n1783_; 
wire alu__abc_42281_new_n1784_; 
wire alu__abc_42281_new_n1785_; 
wire alu__abc_42281_new_n1786_; 
wire alu__abc_42281_new_n1787_; 
wire alu__abc_42281_new_n1788_; 
wire alu__abc_42281_new_n1789_; 
wire alu__abc_42281_new_n178_; 
wire alu__abc_42281_new_n1790_; 
wire alu__abc_42281_new_n1792_; 
wire alu__abc_42281_new_n1793_; 
wire alu__abc_42281_new_n1794_; 
wire alu__abc_42281_new_n1795_; 
wire alu__abc_42281_new_n1796_; 
wire alu__abc_42281_new_n1797_; 
wire alu__abc_42281_new_n1798_; 
wire alu__abc_42281_new_n1799_; 
wire alu__abc_42281_new_n179_; 
wire alu__abc_42281_new_n1800_; 
wire alu__abc_42281_new_n1801_; 
wire alu__abc_42281_new_n1802_; 
wire alu__abc_42281_new_n1803_; 
wire alu__abc_42281_new_n1804_; 
wire alu__abc_42281_new_n1805_; 
wire alu__abc_42281_new_n1806_; 
wire alu__abc_42281_new_n1807_; 
wire alu__abc_42281_new_n1808_; 
wire alu__abc_42281_new_n1809_; 
wire alu__abc_42281_new_n180_; 
wire alu__abc_42281_new_n1810_; 
wire alu__abc_42281_new_n1811_; 
wire alu__abc_42281_new_n1812_; 
wire alu__abc_42281_new_n1813_; 
wire alu__abc_42281_new_n1814_; 
wire alu__abc_42281_new_n1815_; 
wire alu__abc_42281_new_n1816_; 
wire alu__abc_42281_new_n1817_; 
wire alu__abc_42281_new_n1818_; 
wire alu__abc_42281_new_n1819_; 
wire alu__abc_42281_new_n181_; 
wire alu__abc_42281_new_n1820_; 
wire alu__abc_42281_new_n1821_; 
wire alu__abc_42281_new_n1822_; 
wire alu__abc_42281_new_n1823_; 
wire alu__abc_42281_new_n1824_; 
wire alu__abc_42281_new_n1825_; 
wire alu__abc_42281_new_n1826_; 
wire alu__abc_42281_new_n1827_; 
wire alu__abc_42281_new_n1828_; 
wire alu__abc_42281_new_n1829_; 
wire alu__abc_42281_new_n182_; 
wire alu__abc_42281_new_n1830_; 
wire alu__abc_42281_new_n1832_; 
wire alu__abc_42281_new_n1833_; 
wire alu__abc_42281_new_n1834_; 
wire alu__abc_42281_new_n1835_; 
wire alu__abc_42281_new_n1836_; 
wire alu__abc_42281_new_n1837_; 
wire alu__abc_42281_new_n1838_; 
wire alu__abc_42281_new_n1839_; 
wire alu__abc_42281_new_n183_; 
wire alu__abc_42281_new_n1840_; 
wire alu__abc_42281_new_n1841_; 
wire alu__abc_42281_new_n1842_; 
wire alu__abc_42281_new_n1843_; 
wire alu__abc_42281_new_n1844_; 
wire alu__abc_42281_new_n1845_; 
wire alu__abc_42281_new_n1846_; 
wire alu__abc_42281_new_n1847_; 
wire alu__abc_42281_new_n1848_; 
wire alu__abc_42281_new_n1849_; 
wire alu__abc_42281_new_n184_; 
wire alu__abc_42281_new_n1850_; 
wire alu__abc_42281_new_n1851_; 
wire alu__abc_42281_new_n1852_; 
wire alu__abc_42281_new_n1853_; 
wire alu__abc_42281_new_n1854_; 
wire alu__abc_42281_new_n1855_; 
wire alu__abc_42281_new_n1856_; 
wire alu__abc_42281_new_n1857_; 
wire alu__abc_42281_new_n1858_; 
wire alu__abc_42281_new_n1859_; 
wire alu__abc_42281_new_n185_; 
wire alu__abc_42281_new_n1860_; 
wire alu__abc_42281_new_n1861_; 
wire alu__abc_42281_new_n1862_; 
wire alu__abc_42281_new_n1863_; 
wire alu__abc_42281_new_n1864_; 
wire alu__abc_42281_new_n1865_; 
wire alu__abc_42281_new_n1866_; 
wire alu__abc_42281_new_n1867_; 
wire alu__abc_42281_new_n1868_; 
wire alu__abc_42281_new_n1869_; 
wire alu__abc_42281_new_n186_; 
wire alu__abc_42281_new_n1870_; 
wire alu__abc_42281_new_n1871_; 
wire alu__abc_42281_new_n1872_; 
wire alu__abc_42281_new_n1873_; 
wire alu__abc_42281_new_n1874_; 
wire alu__abc_42281_new_n1876_; 
wire alu__abc_42281_new_n1877_; 
wire alu__abc_42281_new_n1878_; 
wire alu__abc_42281_new_n1879_; 
wire alu__abc_42281_new_n187_; 
wire alu__abc_42281_new_n1880_; 
wire alu__abc_42281_new_n1881_; 
wire alu__abc_42281_new_n1882_; 
wire alu__abc_42281_new_n1883_; 
wire alu__abc_42281_new_n1884_; 
wire alu__abc_42281_new_n1885_; 
wire alu__abc_42281_new_n1886_; 
wire alu__abc_42281_new_n1887_; 
wire alu__abc_42281_new_n1888_; 
wire alu__abc_42281_new_n1889_; 
wire alu__abc_42281_new_n188_; 
wire alu__abc_42281_new_n1890_; 
wire alu__abc_42281_new_n1891_; 
wire alu__abc_42281_new_n1892_; 
wire alu__abc_42281_new_n1893_; 
wire alu__abc_42281_new_n1894_; 
wire alu__abc_42281_new_n1895_; 
wire alu__abc_42281_new_n1896_; 
wire alu__abc_42281_new_n1897_; 
wire alu__abc_42281_new_n1898_; 
wire alu__abc_42281_new_n1899_; 
wire alu__abc_42281_new_n189_; 
wire alu__abc_42281_new_n1900_; 
wire alu__abc_42281_new_n1901_; 
wire alu__abc_42281_new_n1902_; 
wire alu__abc_42281_new_n1903_; 
wire alu__abc_42281_new_n1904_; 
wire alu__abc_42281_new_n1905_; 
wire alu__abc_42281_new_n1906_; 
wire alu__abc_42281_new_n1907_; 
wire alu__abc_42281_new_n1908_; 
wire alu__abc_42281_new_n1909_; 
wire alu__abc_42281_new_n190_; 
wire alu__abc_42281_new_n1910_; 
wire alu__abc_42281_new_n1911_; 
wire alu__abc_42281_new_n1912_; 
wire alu__abc_42281_new_n1913_; 
wire alu__abc_42281_new_n1914_; 
wire alu__abc_42281_new_n1915_; 
wire alu__abc_42281_new_n1917_; 
wire alu__abc_42281_new_n1918_; 
wire alu__abc_42281_new_n1919_; 
wire alu__abc_42281_new_n191_; 
wire alu__abc_42281_new_n1920_; 
wire alu__abc_42281_new_n1921_; 
wire alu__abc_42281_new_n1922_; 
wire alu__abc_42281_new_n1923_; 
wire alu__abc_42281_new_n1924_; 
wire alu__abc_42281_new_n1925_; 
wire alu__abc_42281_new_n1926_; 
wire alu__abc_42281_new_n1927_; 
wire alu__abc_42281_new_n1928_; 
wire alu__abc_42281_new_n1929_; 
wire alu__abc_42281_new_n192_; 
wire alu__abc_42281_new_n1930_; 
wire alu__abc_42281_new_n1931_; 
wire alu__abc_42281_new_n1932_; 
wire alu__abc_42281_new_n1933_; 
wire alu__abc_42281_new_n1934_; 
wire alu__abc_42281_new_n1935_; 
wire alu__abc_42281_new_n1936_; 
wire alu__abc_42281_new_n1937_; 
wire alu__abc_42281_new_n1938_; 
wire alu__abc_42281_new_n1939_; 
wire alu__abc_42281_new_n193_; 
wire alu__abc_42281_new_n1940_; 
wire alu__abc_42281_new_n1941_; 
wire alu__abc_42281_new_n1942_; 
wire alu__abc_42281_new_n1943_; 
wire alu__abc_42281_new_n1944_; 
wire alu__abc_42281_new_n1945_; 
wire alu__abc_42281_new_n1946_; 
wire alu__abc_42281_new_n1947_; 
wire alu__abc_42281_new_n1948_; 
wire alu__abc_42281_new_n1949_; 
wire alu__abc_42281_new_n194_; 
wire alu__abc_42281_new_n1950_; 
wire alu__abc_42281_new_n1951_; 
wire alu__abc_42281_new_n1952_; 
wire alu__abc_42281_new_n1953_; 
wire alu__abc_42281_new_n1954_; 
wire alu__abc_42281_new_n1955_; 
wire alu__abc_42281_new_n1957_; 
wire alu__abc_42281_new_n1958_; 
wire alu__abc_42281_new_n1959_; 
wire alu__abc_42281_new_n195_; 
wire alu__abc_42281_new_n1960_; 
wire alu__abc_42281_new_n1961_; 
wire alu__abc_42281_new_n1962_; 
wire alu__abc_42281_new_n1963_; 
wire alu__abc_42281_new_n1964_; 
wire alu__abc_42281_new_n1965_; 
wire alu__abc_42281_new_n1966_; 
wire alu__abc_42281_new_n1967_; 
wire alu__abc_42281_new_n1968_; 
wire alu__abc_42281_new_n1969_; 
wire alu__abc_42281_new_n196_; 
wire alu__abc_42281_new_n1970_; 
wire alu__abc_42281_new_n1971_; 
wire alu__abc_42281_new_n1972_; 
wire alu__abc_42281_new_n1973_; 
wire alu__abc_42281_new_n1974_; 
wire alu__abc_42281_new_n1975_; 
wire alu__abc_42281_new_n1976_; 
wire alu__abc_42281_new_n1977_; 
wire alu__abc_42281_new_n1978_; 
wire alu__abc_42281_new_n1979_; 
wire alu__abc_42281_new_n197_; 
wire alu__abc_42281_new_n1980_; 
wire alu__abc_42281_new_n1981_; 
wire alu__abc_42281_new_n1982_; 
wire alu__abc_42281_new_n1983_; 
wire alu__abc_42281_new_n1984_; 
wire alu__abc_42281_new_n1985_; 
wire alu__abc_42281_new_n1986_; 
wire alu__abc_42281_new_n1987_; 
wire alu__abc_42281_new_n1988_; 
wire alu__abc_42281_new_n1989_; 
wire alu__abc_42281_new_n198_; 
wire alu__abc_42281_new_n1990_; 
wire alu__abc_42281_new_n1991_; 
wire alu__abc_42281_new_n1992_; 
wire alu__abc_42281_new_n1993_; 
wire alu__abc_42281_new_n1994_; 
wire alu__abc_42281_new_n1995_; 
wire alu__abc_42281_new_n1997_; 
wire alu__abc_42281_new_n1998_; 
wire alu__abc_42281_new_n1999_; 
wire alu__abc_42281_new_n199_; 
wire alu__abc_42281_new_n2000_; 
wire alu__abc_42281_new_n2001_; 
wire alu__abc_42281_new_n2002_; 
wire alu__abc_42281_new_n2003_; 
wire alu__abc_42281_new_n2004_; 
wire alu__abc_42281_new_n2005_; 
wire alu__abc_42281_new_n2006_; 
wire alu__abc_42281_new_n2007_; 
wire alu__abc_42281_new_n2008_; 
wire alu__abc_42281_new_n2009_; 
wire alu__abc_42281_new_n200_; 
wire alu__abc_42281_new_n2010_; 
wire alu__abc_42281_new_n2011_; 
wire alu__abc_42281_new_n2012_; 
wire alu__abc_42281_new_n2013_; 
wire alu__abc_42281_new_n2014_; 
wire alu__abc_42281_new_n2015_; 
wire alu__abc_42281_new_n2016_; 
wire alu__abc_42281_new_n2017_; 
wire alu__abc_42281_new_n2018_; 
wire alu__abc_42281_new_n2019_; 
wire alu__abc_42281_new_n201_; 
wire alu__abc_42281_new_n2020_; 
wire alu__abc_42281_new_n2021_; 
wire alu__abc_42281_new_n2022_; 
wire alu__abc_42281_new_n2023_; 
wire alu__abc_42281_new_n2024_; 
wire alu__abc_42281_new_n2025_; 
wire alu__abc_42281_new_n2026_; 
wire alu__abc_42281_new_n2027_; 
wire alu__abc_42281_new_n2028_; 
wire alu__abc_42281_new_n2029_; 
wire alu__abc_42281_new_n202_; 
wire alu__abc_42281_new_n2030_; 
wire alu__abc_42281_new_n2031_; 
wire alu__abc_42281_new_n2032_; 
wire alu__abc_42281_new_n2033_; 
wire alu__abc_42281_new_n2034_; 
wire alu__abc_42281_new_n2035_; 
wire alu__abc_42281_new_n2036_; 
wire alu__abc_42281_new_n2038_; 
wire alu__abc_42281_new_n2039_; 
wire alu__abc_42281_new_n203_; 
wire alu__abc_42281_new_n2040_; 
wire alu__abc_42281_new_n2041_; 
wire alu__abc_42281_new_n2042_; 
wire alu__abc_42281_new_n2043_; 
wire alu__abc_42281_new_n2044_; 
wire alu__abc_42281_new_n2045_; 
wire alu__abc_42281_new_n2046_; 
wire alu__abc_42281_new_n2047_; 
wire alu__abc_42281_new_n2048_; 
wire alu__abc_42281_new_n2049_; 
wire alu__abc_42281_new_n204_; 
wire alu__abc_42281_new_n2050_; 
wire alu__abc_42281_new_n2051_; 
wire alu__abc_42281_new_n2052_; 
wire alu__abc_42281_new_n2053_; 
wire alu__abc_42281_new_n2054_; 
wire alu__abc_42281_new_n2055_; 
wire alu__abc_42281_new_n2056_; 
wire alu__abc_42281_new_n2057_; 
wire alu__abc_42281_new_n2058_; 
wire alu__abc_42281_new_n2059_; 
wire alu__abc_42281_new_n205_; 
wire alu__abc_42281_new_n2060_; 
wire alu__abc_42281_new_n2061_; 
wire alu__abc_42281_new_n2062_; 
wire alu__abc_42281_new_n2063_; 
wire alu__abc_42281_new_n2064_; 
wire alu__abc_42281_new_n2065_; 
wire alu__abc_42281_new_n2066_; 
wire alu__abc_42281_new_n2067_; 
wire alu__abc_42281_new_n2068_; 
wire alu__abc_42281_new_n2069_; 
wire alu__abc_42281_new_n206_; 
wire alu__abc_42281_new_n2070_; 
wire alu__abc_42281_new_n2071_; 
wire alu__abc_42281_new_n2072_; 
wire alu__abc_42281_new_n2073_; 
wire alu__abc_42281_new_n2074_; 
wire alu__abc_42281_new_n2075_; 
wire alu__abc_42281_new_n2076_; 
wire alu__abc_42281_new_n2077_; 
wire alu__abc_42281_new_n2079_; 
wire alu__abc_42281_new_n207_; 
wire alu__abc_42281_new_n2080_; 
wire alu__abc_42281_new_n2081_; 
wire alu__abc_42281_new_n2082_; 
wire alu__abc_42281_new_n2083_; 
wire alu__abc_42281_new_n2084_; 
wire alu__abc_42281_new_n2085_; 
wire alu__abc_42281_new_n2086_; 
wire alu__abc_42281_new_n2087_; 
wire alu__abc_42281_new_n2088_; 
wire alu__abc_42281_new_n2089_; 
wire alu__abc_42281_new_n208_; 
wire alu__abc_42281_new_n2090_; 
wire alu__abc_42281_new_n2091_; 
wire alu__abc_42281_new_n2092_; 
wire alu__abc_42281_new_n2093_; 
wire alu__abc_42281_new_n2094_; 
wire alu__abc_42281_new_n2095_; 
wire alu__abc_42281_new_n2096_; 
wire alu__abc_42281_new_n2097_; 
wire alu__abc_42281_new_n2098_; 
wire alu__abc_42281_new_n2099_; 
wire alu__abc_42281_new_n209_; 
wire alu__abc_42281_new_n2100_; 
wire alu__abc_42281_new_n2101_; 
wire alu__abc_42281_new_n2102_; 
wire alu__abc_42281_new_n2103_; 
wire alu__abc_42281_new_n2104_; 
wire alu__abc_42281_new_n2105_; 
wire alu__abc_42281_new_n2106_; 
wire alu__abc_42281_new_n2107_; 
wire alu__abc_42281_new_n2108_; 
wire alu__abc_42281_new_n2109_; 
wire alu__abc_42281_new_n210_; 
wire alu__abc_42281_new_n2110_; 
wire alu__abc_42281_new_n2111_; 
wire alu__abc_42281_new_n2112_; 
wire alu__abc_42281_new_n2113_; 
wire alu__abc_42281_new_n2114_; 
wire alu__abc_42281_new_n2115_; 
wire alu__abc_42281_new_n2116_; 
wire alu__abc_42281_new_n2117_; 
wire alu__abc_42281_new_n2118_; 
wire alu__abc_42281_new_n211_; 
wire alu__abc_42281_new_n2120_; 
wire alu__abc_42281_new_n2121_; 
wire alu__abc_42281_new_n2122_; 
wire alu__abc_42281_new_n2123_; 
wire alu__abc_42281_new_n2124_; 
wire alu__abc_42281_new_n2125_; 
wire alu__abc_42281_new_n2126_; 
wire alu__abc_42281_new_n2127_; 
wire alu__abc_42281_new_n2128_; 
wire alu__abc_42281_new_n2129_; 
wire alu__abc_42281_new_n212_; 
wire alu__abc_42281_new_n2130_; 
wire alu__abc_42281_new_n2131_; 
wire alu__abc_42281_new_n2132_; 
wire alu__abc_42281_new_n2133_; 
wire alu__abc_42281_new_n2134_; 
wire alu__abc_42281_new_n2135_; 
wire alu__abc_42281_new_n2136_; 
wire alu__abc_42281_new_n2137_; 
wire alu__abc_42281_new_n2138_; 
wire alu__abc_42281_new_n2139_; 
wire alu__abc_42281_new_n213_; 
wire alu__abc_42281_new_n2140_; 
wire alu__abc_42281_new_n2141_; 
wire alu__abc_42281_new_n2142_; 
wire alu__abc_42281_new_n2143_; 
wire alu__abc_42281_new_n2144_; 
wire alu__abc_42281_new_n2145_; 
wire alu__abc_42281_new_n2146_; 
wire alu__abc_42281_new_n2147_; 
wire alu__abc_42281_new_n2148_; 
wire alu__abc_42281_new_n2149_; 
wire alu__abc_42281_new_n214_; 
wire alu__abc_42281_new_n2150_; 
wire alu__abc_42281_new_n2151_; 
wire alu__abc_42281_new_n2152_; 
wire alu__abc_42281_new_n2153_; 
wire alu__abc_42281_new_n2154_; 
wire alu__abc_42281_new_n2155_; 
wire alu__abc_42281_new_n2156_; 
wire alu__abc_42281_new_n2157_; 
wire alu__abc_42281_new_n2159_; 
wire alu__abc_42281_new_n215_; 
wire alu__abc_42281_new_n2160_; 
wire alu__abc_42281_new_n2161_; 
wire alu__abc_42281_new_n2162_; 
wire alu__abc_42281_new_n2163_; 
wire alu__abc_42281_new_n2164_; 
wire alu__abc_42281_new_n2165_; 
wire alu__abc_42281_new_n2166_; 
wire alu__abc_42281_new_n2167_; 
wire alu__abc_42281_new_n2168_; 
wire alu__abc_42281_new_n2169_; 
wire alu__abc_42281_new_n216_; 
wire alu__abc_42281_new_n2170_; 
wire alu__abc_42281_new_n2171_; 
wire alu__abc_42281_new_n2172_; 
wire alu__abc_42281_new_n2173_; 
wire alu__abc_42281_new_n2174_; 
wire alu__abc_42281_new_n2175_; 
wire alu__abc_42281_new_n2176_; 
wire alu__abc_42281_new_n2177_; 
wire alu__abc_42281_new_n2178_; 
wire alu__abc_42281_new_n2179_; 
wire alu__abc_42281_new_n217_; 
wire alu__abc_42281_new_n2180_; 
wire alu__abc_42281_new_n2181_; 
wire alu__abc_42281_new_n2182_; 
wire alu__abc_42281_new_n2183_; 
wire alu__abc_42281_new_n2184_; 
wire alu__abc_42281_new_n2185_; 
wire alu__abc_42281_new_n2186_; 
wire alu__abc_42281_new_n2187_; 
wire alu__abc_42281_new_n2188_; 
wire alu__abc_42281_new_n2189_; 
wire alu__abc_42281_new_n218_; 
wire alu__abc_42281_new_n2190_; 
wire alu__abc_42281_new_n2191_; 
wire alu__abc_42281_new_n2192_; 
wire alu__abc_42281_new_n2193_; 
wire alu__abc_42281_new_n2194_; 
wire alu__abc_42281_new_n2195_; 
wire alu__abc_42281_new_n2196_; 
wire alu__abc_42281_new_n2198_; 
wire alu__abc_42281_new_n2199_; 
wire alu__abc_42281_new_n219_; 
wire alu__abc_42281_new_n2200_; 
wire alu__abc_42281_new_n2201_; 
wire alu__abc_42281_new_n2202_; 
wire alu__abc_42281_new_n2203_; 
wire alu__abc_42281_new_n2204_; 
wire alu__abc_42281_new_n2205_; 
wire alu__abc_42281_new_n2206_; 
wire alu__abc_42281_new_n2207_; 
wire alu__abc_42281_new_n2208_; 
wire alu__abc_42281_new_n2209_; 
wire alu__abc_42281_new_n220_; 
wire alu__abc_42281_new_n2210_; 
wire alu__abc_42281_new_n2211_; 
wire alu__abc_42281_new_n2212_; 
wire alu__abc_42281_new_n2213_; 
wire alu__abc_42281_new_n2214_; 
wire alu__abc_42281_new_n2215_; 
wire alu__abc_42281_new_n2216_; 
wire alu__abc_42281_new_n2217_; 
wire alu__abc_42281_new_n2218_; 
wire alu__abc_42281_new_n2219_; 
wire alu__abc_42281_new_n221_; 
wire alu__abc_42281_new_n2220_; 
wire alu__abc_42281_new_n2221_; 
wire alu__abc_42281_new_n2222_; 
wire alu__abc_42281_new_n2223_; 
wire alu__abc_42281_new_n2224_; 
wire alu__abc_42281_new_n2225_; 
wire alu__abc_42281_new_n2226_; 
wire alu__abc_42281_new_n2227_; 
wire alu__abc_42281_new_n2228_; 
wire alu__abc_42281_new_n2229_; 
wire alu__abc_42281_new_n222_; 
wire alu__abc_42281_new_n2230_; 
wire alu__abc_42281_new_n2231_; 
wire alu__abc_42281_new_n2232_; 
wire alu__abc_42281_new_n2233_; 
wire alu__abc_42281_new_n2234_; 
wire alu__abc_42281_new_n2235_; 
wire alu__abc_42281_new_n2236_; 
wire alu__abc_42281_new_n2237_; 
wire alu__abc_42281_new_n2238_; 
wire alu__abc_42281_new_n223_; 
wire alu__abc_42281_new_n2240_; 
wire alu__abc_42281_new_n2241_; 
wire alu__abc_42281_new_n2242_; 
wire alu__abc_42281_new_n2243_; 
wire alu__abc_42281_new_n2244_; 
wire alu__abc_42281_new_n2245_; 
wire alu__abc_42281_new_n2246_; 
wire alu__abc_42281_new_n2247_; 
wire alu__abc_42281_new_n2248_; 
wire alu__abc_42281_new_n2249_; 
wire alu__abc_42281_new_n224_; 
wire alu__abc_42281_new_n2250_; 
wire alu__abc_42281_new_n2251_; 
wire alu__abc_42281_new_n2252_; 
wire alu__abc_42281_new_n2253_; 
wire alu__abc_42281_new_n2254_; 
wire alu__abc_42281_new_n2255_; 
wire alu__abc_42281_new_n2256_; 
wire alu__abc_42281_new_n2257_; 
wire alu__abc_42281_new_n2258_; 
wire alu__abc_42281_new_n2259_; 
wire alu__abc_42281_new_n225_; 
wire alu__abc_42281_new_n2260_; 
wire alu__abc_42281_new_n2261_; 
wire alu__abc_42281_new_n2262_; 
wire alu__abc_42281_new_n2263_; 
wire alu__abc_42281_new_n2264_; 
wire alu__abc_42281_new_n2265_; 
wire alu__abc_42281_new_n2266_; 
wire alu__abc_42281_new_n2267_; 
wire alu__abc_42281_new_n2268_; 
wire alu__abc_42281_new_n2269_; 
wire alu__abc_42281_new_n226_; 
wire alu__abc_42281_new_n2270_; 
wire alu__abc_42281_new_n2271_; 
wire alu__abc_42281_new_n2272_; 
wire alu__abc_42281_new_n2273_; 
wire alu__abc_42281_new_n2274_; 
wire alu__abc_42281_new_n2275_; 
wire alu__abc_42281_new_n2276_; 
wire alu__abc_42281_new_n2277_; 
wire alu__abc_42281_new_n2278_; 
wire alu__abc_42281_new_n2279_; 
wire alu__abc_42281_new_n227_; 
wire alu__abc_42281_new_n2281_; 
wire alu__abc_42281_new_n2282_; 
wire alu__abc_42281_new_n2283_; 
wire alu__abc_42281_new_n2284_; 
wire alu__abc_42281_new_n2285_; 
wire alu__abc_42281_new_n2286_; 
wire alu__abc_42281_new_n2287_; 
wire alu__abc_42281_new_n2288_; 
wire alu__abc_42281_new_n2289_; 
wire alu__abc_42281_new_n228_; 
wire alu__abc_42281_new_n2290_; 
wire alu__abc_42281_new_n2291_; 
wire alu__abc_42281_new_n2292_; 
wire alu__abc_42281_new_n2293_; 
wire alu__abc_42281_new_n2294_; 
wire alu__abc_42281_new_n2295_; 
wire alu__abc_42281_new_n2296_; 
wire alu__abc_42281_new_n2297_; 
wire alu__abc_42281_new_n2298_; 
wire alu__abc_42281_new_n2299_; 
wire alu__abc_42281_new_n229_; 
wire alu__abc_42281_new_n2300_; 
wire alu__abc_42281_new_n2301_; 
wire alu__abc_42281_new_n2302_; 
wire alu__abc_42281_new_n2303_; 
wire alu__abc_42281_new_n2304_; 
wire alu__abc_42281_new_n2305_; 
wire alu__abc_42281_new_n2306_; 
wire alu__abc_42281_new_n2307_; 
wire alu__abc_42281_new_n2308_; 
wire alu__abc_42281_new_n2309_; 
wire alu__abc_42281_new_n230_; 
wire alu__abc_42281_new_n2310_; 
wire alu__abc_42281_new_n2311_; 
wire alu__abc_42281_new_n2312_; 
wire alu__abc_42281_new_n2313_; 
wire alu__abc_42281_new_n2314_; 
wire alu__abc_42281_new_n2315_; 
wire alu__abc_42281_new_n2316_; 
wire alu__abc_42281_new_n2317_; 
wire alu__abc_42281_new_n2319_; 
wire alu__abc_42281_new_n231_; 
wire alu__abc_42281_new_n2320_; 
wire alu__abc_42281_new_n2321_; 
wire alu__abc_42281_new_n2322_; 
wire alu__abc_42281_new_n2323_; 
wire alu__abc_42281_new_n2324_; 
wire alu__abc_42281_new_n2325_; 
wire alu__abc_42281_new_n2326_; 
wire alu__abc_42281_new_n2327_; 
wire alu__abc_42281_new_n2328_; 
wire alu__abc_42281_new_n2329_; 
wire alu__abc_42281_new_n232_; 
wire alu__abc_42281_new_n2330_; 
wire alu__abc_42281_new_n2331_; 
wire alu__abc_42281_new_n2332_; 
wire alu__abc_42281_new_n2333_; 
wire alu__abc_42281_new_n2334_; 
wire alu__abc_42281_new_n2335_; 
wire alu__abc_42281_new_n2336_; 
wire alu__abc_42281_new_n2337_; 
wire alu__abc_42281_new_n2338_; 
wire alu__abc_42281_new_n2339_; 
wire alu__abc_42281_new_n233_; 
wire alu__abc_42281_new_n2340_; 
wire alu__abc_42281_new_n2341_; 
wire alu__abc_42281_new_n2342_; 
wire alu__abc_42281_new_n2343_; 
wire alu__abc_42281_new_n2344_; 
wire alu__abc_42281_new_n2345_; 
wire alu__abc_42281_new_n2346_; 
wire alu__abc_42281_new_n2347_; 
wire alu__abc_42281_new_n2348_; 
wire alu__abc_42281_new_n2349_; 
wire alu__abc_42281_new_n234_; 
wire alu__abc_42281_new_n2350_; 
wire alu__abc_42281_new_n2351_; 
wire alu__abc_42281_new_n2352_; 
wire alu__abc_42281_new_n2353_; 
wire alu__abc_42281_new_n2354_; 
wire alu__abc_42281_new_n2355_; 
wire alu__abc_42281_new_n2356_; 
wire alu__abc_42281_new_n2357_; 
wire alu__abc_42281_new_n2358_; 
wire alu__abc_42281_new_n235_; 
wire alu__abc_42281_new_n2360_; 
wire alu__abc_42281_new_n2361_; 
wire alu__abc_42281_new_n2362_; 
wire alu__abc_42281_new_n2363_; 
wire alu__abc_42281_new_n2364_; 
wire alu__abc_42281_new_n2365_; 
wire alu__abc_42281_new_n2366_; 
wire alu__abc_42281_new_n2367_; 
wire alu__abc_42281_new_n2368_; 
wire alu__abc_42281_new_n2369_; 
wire alu__abc_42281_new_n236_; 
wire alu__abc_42281_new_n2370_; 
wire alu__abc_42281_new_n2371_; 
wire alu__abc_42281_new_n2372_; 
wire alu__abc_42281_new_n2373_; 
wire alu__abc_42281_new_n2374_; 
wire alu__abc_42281_new_n2375_; 
wire alu__abc_42281_new_n2376_; 
wire alu__abc_42281_new_n2377_; 
wire alu__abc_42281_new_n2378_; 
wire alu__abc_42281_new_n2379_; 
wire alu__abc_42281_new_n237_; 
wire alu__abc_42281_new_n2380_; 
wire alu__abc_42281_new_n2381_; 
wire alu__abc_42281_new_n2382_; 
wire alu__abc_42281_new_n2383_; 
wire alu__abc_42281_new_n2384_; 
wire alu__abc_42281_new_n2385_; 
wire alu__abc_42281_new_n2386_; 
wire alu__abc_42281_new_n2387_; 
wire alu__abc_42281_new_n2388_; 
wire alu__abc_42281_new_n2389_; 
wire alu__abc_42281_new_n238_; 
wire alu__abc_42281_new_n2390_; 
wire alu__abc_42281_new_n2391_; 
wire alu__abc_42281_new_n2392_; 
wire alu__abc_42281_new_n2393_; 
wire alu__abc_42281_new_n2394_; 
wire alu__abc_42281_new_n2395_; 
wire alu__abc_42281_new_n2397_; 
wire alu__abc_42281_new_n2398_; 
wire alu__abc_42281_new_n2399_; 
wire alu__abc_42281_new_n239_; 
wire alu__abc_42281_new_n2400_; 
wire alu__abc_42281_new_n2401_; 
wire alu__abc_42281_new_n2402_; 
wire alu__abc_42281_new_n2403_; 
wire alu__abc_42281_new_n2404_; 
wire alu__abc_42281_new_n2405_; 
wire alu__abc_42281_new_n2406_; 
wire alu__abc_42281_new_n2407_; 
wire alu__abc_42281_new_n2408_; 
wire alu__abc_42281_new_n2409_; 
wire alu__abc_42281_new_n240_; 
wire alu__abc_42281_new_n2410_; 
wire alu__abc_42281_new_n2411_; 
wire alu__abc_42281_new_n2412_; 
wire alu__abc_42281_new_n2413_; 
wire alu__abc_42281_new_n2414_; 
wire alu__abc_42281_new_n2415_; 
wire alu__abc_42281_new_n2416_; 
wire alu__abc_42281_new_n2417_; 
wire alu__abc_42281_new_n2418_; 
wire alu__abc_42281_new_n2419_; 
wire alu__abc_42281_new_n241_; 
wire alu__abc_42281_new_n2420_; 
wire alu__abc_42281_new_n2421_; 
wire alu__abc_42281_new_n2422_; 
wire alu__abc_42281_new_n2423_; 
wire alu__abc_42281_new_n2424_; 
wire alu__abc_42281_new_n2425_; 
wire alu__abc_42281_new_n2426_; 
wire alu__abc_42281_new_n2427_; 
wire alu__abc_42281_new_n2428_; 
wire alu__abc_42281_new_n2429_; 
wire alu__abc_42281_new_n242_; 
wire alu__abc_42281_new_n2430_; 
wire alu__abc_42281_new_n2431_; 
wire alu__abc_42281_new_n2433_; 
wire alu__abc_42281_new_n2434_; 
wire alu__abc_42281_new_n2436_; 
wire alu__abc_42281_new_n2437_; 
wire alu__abc_42281_new_n2438_; 
wire alu__abc_42281_new_n2439_; 
wire alu__abc_42281_new_n243_; 
wire alu__abc_42281_new_n2440_; 
wire alu__abc_42281_new_n2441_; 
wire alu__abc_42281_new_n2442_; 
wire alu__abc_42281_new_n2443_; 
wire alu__abc_42281_new_n2444_; 
wire alu__abc_42281_new_n2445_; 
wire alu__abc_42281_new_n2446_; 
wire alu__abc_42281_new_n2447_; 
wire alu__abc_42281_new_n2448_; 
wire alu__abc_42281_new_n2449_; 
wire alu__abc_42281_new_n244_; 
wire alu__abc_42281_new_n2450_; 
wire alu__abc_42281_new_n2451_; 
wire alu__abc_42281_new_n2452_; 
wire alu__abc_42281_new_n2453_; 
wire alu__abc_42281_new_n2454_; 
wire alu__abc_42281_new_n2455_; 
wire alu__abc_42281_new_n2456_; 
wire alu__abc_42281_new_n2457_; 
wire alu__abc_42281_new_n2458_; 
wire alu__abc_42281_new_n2459_; 
wire alu__abc_42281_new_n245_; 
wire alu__abc_42281_new_n2460_; 
wire alu__abc_42281_new_n2461_; 
wire alu__abc_42281_new_n2462_; 
wire alu__abc_42281_new_n2463_; 
wire alu__abc_42281_new_n2464_; 
wire alu__abc_42281_new_n2465_; 
wire alu__abc_42281_new_n2466_; 
wire alu__abc_42281_new_n2467_; 
wire alu__abc_42281_new_n2468_; 
wire alu__abc_42281_new_n2469_; 
wire alu__abc_42281_new_n246_; 
wire alu__abc_42281_new_n2470_; 
wire alu__abc_42281_new_n2471_; 
wire alu__abc_42281_new_n2472_; 
wire alu__abc_42281_new_n2473_; 
wire alu__abc_42281_new_n2474_; 
wire alu__abc_42281_new_n2475_; 
wire alu__abc_42281_new_n2476_; 
wire alu__abc_42281_new_n2477_; 
wire alu__abc_42281_new_n2478_; 
wire alu__abc_42281_new_n2479_; 
wire alu__abc_42281_new_n247_; 
wire alu__abc_42281_new_n2480_; 
wire alu__abc_42281_new_n2481_; 
wire alu__abc_42281_new_n2482_; 
wire alu__abc_42281_new_n2483_; 
wire alu__abc_42281_new_n2484_; 
wire alu__abc_42281_new_n2485_; 
wire alu__abc_42281_new_n2486_; 
wire alu__abc_42281_new_n2487_; 
wire alu__abc_42281_new_n2488_; 
wire alu__abc_42281_new_n2489_; 
wire alu__abc_42281_new_n248_; 
wire alu__abc_42281_new_n2490_; 
wire alu__abc_42281_new_n2491_; 
wire alu__abc_42281_new_n2492_; 
wire alu__abc_42281_new_n2493_; 
wire alu__abc_42281_new_n2494_; 
wire alu__abc_42281_new_n2495_; 
wire alu__abc_42281_new_n2496_; 
wire alu__abc_42281_new_n2497_; 
wire alu__abc_42281_new_n2498_; 
wire alu__abc_42281_new_n2499_; 
wire alu__abc_42281_new_n249_; 
wire alu__abc_42281_new_n2500_; 
wire alu__abc_42281_new_n2501_; 
wire alu__abc_42281_new_n2502_; 
wire alu__abc_42281_new_n2503_; 
wire alu__abc_42281_new_n2504_; 
wire alu__abc_42281_new_n2505_; 
wire alu__abc_42281_new_n2506_; 
wire alu__abc_42281_new_n2507_; 
wire alu__abc_42281_new_n2508_; 
wire alu__abc_42281_new_n2509_; 
wire alu__abc_42281_new_n250_; 
wire alu__abc_42281_new_n2510_; 
wire alu__abc_42281_new_n2511_; 
wire alu__abc_42281_new_n2512_; 
wire alu__abc_42281_new_n2513_; 
wire alu__abc_42281_new_n2514_; 
wire alu__abc_42281_new_n2515_; 
wire alu__abc_42281_new_n2516_; 
wire alu__abc_42281_new_n2517_; 
wire alu__abc_42281_new_n2518_; 
wire alu__abc_42281_new_n2519_; 
wire alu__abc_42281_new_n251_; 
wire alu__abc_42281_new_n252_; 
wire alu__abc_42281_new_n253_; 
wire alu__abc_42281_new_n254_; 
wire alu__abc_42281_new_n255_; 
wire alu__abc_42281_new_n256_; 
wire alu__abc_42281_new_n257_; 
wire alu__abc_42281_new_n258_; 
wire alu__abc_42281_new_n259_; 
wire alu__abc_42281_new_n260_; 
wire alu__abc_42281_new_n261_; 
wire alu__abc_42281_new_n262_; 
wire alu__abc_42281_new_n263_; 
wire alu__abc_42281_new_n264_; 
wire alu__abc_42281_new_n265_; 
wire alu__abc_42281_new_n266_; 
wire alu__abc_42281_new_n267_; 
wire alu__abc_42281_new_n268_; 
wire alu__abc_42281_new_n269_; 
wire alu__abc_42281_new_n270_; 
wire alu__abc_42281_new_n271_; 
wire alu__abc_42281_new_n271__bF_buf0; 
wire alu__abc_42281_new_n271__bF_buf1; 
wire alu__abc_42281_new_n271__bF_buf2; 
wire alu__abc_42281_new_n271__bF_buf3; 
wire alu__abc_42281_new_n271__bF_buf4; 
wire alu__abc_42281_new_n272_; 
wire alu__abc_42281_new_n273_; 
wire alu__abc_42281_new_n274_; 
wire alu__abc_42281_new_n275_; 
wire alu__abc_42281_new_n276_; 
wire alu__abc_42281_new_n277_; 
wire alu__abc_42281_new_n278_; 
wire alu__abc_42281_new_n279_; 
wire alu__abc_42281_new_n280_; 
wire alu__abc_42281_new_n281_; 
wire alu__abc_42281_new_n281__bF_buf0; 
wire alu__abc_42281_new_n281__bF_buf1; 
wire alu__abc_42281_new_n281__bF_buf2; 
wire alu__abc_42281_new_n281__bF_buf3; 
wire alu__abc_42281_new_n281__bF_buf4; 
wire alu__abc_42281_new_n281__bF_buf5; 
wire alu__abc_42281_new_n281__bF_buf6; 
wire alu__abc_42281_new_n282_; 
wire alu__abc_42281_new_n283_; 
wire alu__abc_42281_new_n284_; 
wire alu__abc_42281_new_n285_; 
wire alu__abc_42281_new_n286_; 
wire alu__abc_42281_new_n287_; 
wire alu__abc_42281_new_n288_; 
wire alu__abc_42281_new_n288__bF_buf0; 
wire alu__abc_42281_new_n288__bF_buf1; 
wire alu__abc_42281_new_n288__bF_buf2; 
wire alu__abc_42281_new_n288__bF_buf3; 
wire alu__abc_42281_new_n288__bF_buf4; 
wire alu__abc_42281_new_n289_; 
wire alu__abc_42281_new_n290_; 
wire alu__abc_42281_new_n291_; 
wire alu__abc_42281_new_n292_; 
wire alu__abc_42281_new_n293_; 
wire alu__abc_42281_new_n294_; 
wire alu__abc_42281_new_n294__bF_buf0; 
wire alu__abc_42281_new_n294__bF_buf1; 
wire alu__abc_42281_new_n294__bF_buf2; 
wire alu__abc_42281_new_n294__bF_buf3; 
wire alu__abc_42281_new_n294__bF_buf4; 
wire alu__abc_42281_new_n294__bF_buf5; 
wire alu__abc_42281_new_n294__bF_buf6; 
wire alu__abc_42281_new_n295_; 
wire alu__abc_42281_new_n296_; 
wire alu__abc_42281_new_n297_; 
wire alu__abc_42281_new_n298_; 
wire alu__abc_42281_new_n299_; 
wire alu__abc_42281_new_n299__bF_buf0; 
wire alu__abc_42281_new_n299__bF_buf1; 
wire alu__abc_42281_new_n299__bF_buf2; 
wire alu__abc_42281_new_n299__bF_buf3; 
wire alu__abc_42281_new_n299__bF_buf4; 
wire alu__abc_42281_new_n299__bF_buf5; 
wire alu__abc_42281_new_n299__bF_buf6; 
wire alu__abc_42281_new_n300_; 
wire alu__abc_42281_new_n301_; 
wire alu__abc_42281_new_n302_; 
wire alu__abc_42281_new_n303_; 
wire alu__abc_42281_new_n304_; 
wire alu__abc_42281_new_n305_; 
wire alu__abc_42281_new_n306_; 
wire alu__abc_42281_new_n307_; 
wire alu__abc_42281_new_n308_; 
wire alu__abc_42281_new_n309_; 
wire alu__abc_42281_new_n310_; 
wire alu__abc_42281_new_n311_; 
wire alu__abc_42281_new_n312_; 
wire alu__abc_42281_new_n313_; 
wire alu__abc_42281_new_n314_; 
wire alu__abc_42281_new_n315_; 
wire alu__abc_42281_new_n316_; 
wire alu__abc_42281_new_n317_; 
wire alu__abc_42281_new_n318_; 
wire alu__abc_42281_new_n319_; 
wire alu__abc_42281_new_n320_; 
wire alu__abc_42281_new_n321_; 
wire alu__abc_42281_new_n322_; 
wire alu__abc_42281_new_n323_; 
wire alu__abc_42281_new_n324_; 
wire alu__abc_42281_new_n325_; 
wire alu__abc_42281_new_n326_; 
wire alu__abc_42281_new_n327_; 
wire alu__abc_42281_new_n328_; 
wire alu__abc_42281_new_n329_; 
wire alu__abc_42281_new_n330_; 
wire alu__abc_42281_new_n331_; 
wire alu__abc_42281_new_n332_; 
wire alu__abc_42281_new_n333_; 
wire alu__abc_42281_new_n334_; 
wire alu__abc_42281_new_n335_; 
wire alu__abc_42281_new_n336_; 
wire alu__abc_42281_new_n337_; 
wire alu__abc_42281_new_n338_; 
wire alu__abc_42281_new_n339_; 
wire alu__abc_42281_new_n340_; 
wire alu__abc_42281_new_n341_; 
wire alu__abc_42281_new_n342_; 
wire alu__abc_42281_new_n343_; 
wire alu__abc_42281_new_n344_; 
wire alu__abc_42281_new_n345_; 
wire alu__abc_42281_new_n346_; 
wire alu__abc_42281_new_n347_; 
wire alu__abc_42281_new_n348_; 
wire alu__abc_42281_new_n349_; 
wire alu__abc_42281_new_n350_; 
wire alu__abc_42281_new_n351_; 
wire alu__abc_42281_new_n352_; 
wire alu__abc_42281_new_n353_; 
wire alu__abc_42281_new_n354_; 
wire alu__abc_42281_new_n355_; 
wire alu__abc_42281_new_n356_; 
wire alu__abc_42281_new_n357_; 
wire alu__abc_42281_new_n358_; 
wire alu__abc_42281_new_n359_; 
wire alu__abc_42281_new_n360_; 
wire alu__abc_42281_new_n361_; 
wire alu__abc_42281_new_n362_; 
wire alu__abc_42281_new_n363_; 
wire alu__abc_42281_new_n364_; 
wire alu__abc_42281_new_n365_; 
wire alu__abc_42281_new_n366_; 
wire alu__abc_42281_new_n367_; 
wire alu__abc_42281_new_n368_; 
wire alu__abc_42281_new_n369_; 
wire alu__abc_42281_new_n370_; 
wire alu__abc_42281_new_n371_; 
wire alu__abc_42281_new_n372_; 
wire alu__abc_42281_new_n373_; 
wire alu__abc_42281_new_n374_; 
wire alu__abc_42281_new_n375_; 
wire alu__abc_42281_new_n376_; 
wire alu__abc_42281_new_n378_; 
wire alu__abc_42281_new_n379_; 
wire alu__abc_42281_new_n380_; 
wire alu__abc_42281_new_n382_; 
wire alu__abc_42281_new_n383_; 
wire alu__abc_42281_new_n384_; 
wire alu__abc_42281_new_n385_; 
wire alu__abc_42281_new_n387_; 
wire alu__abc_42281_new_n388_; 
wire alu__abc_42281_new_n389_; 
wire alu__abc_42281_new_n390_; 
wire alu__abc_42281_new_n391_; 
wire alu__abc_42281_new_n392_; 
wire alu__abc_42281_new_n393_; 
wire alu__abc_42281_new_n394_; 
wire alu__abc_42281_new_n395_; 
wire alu__abc_42281_new_n396_; 
wire alu__abc_42281_new_n397_; 
wire alu__abc_42281_new_n398_; 
wire alu__abc_42281_new_n399_; 
wire alu__abc_42281_new_n400_; 
wire alu__abc_42281_new_n401_; 
wire alu__abc_42281_new_n402_; 
wire alu__abc_42281_new_n403_; 
wire alu__abc_42281_new_n404_; 
wire alu__abc_42281_new_n405_; 
wire alu__abc_42281_new_n406_; 
wire alu__abc_42281_new_n407_; 
wire alu__abc_42281_new_n408_; 
wire alu__abc_42281_new_n409_; 
wire alu__abc_42281_new_n410_; 
wire alu__abc_42281_new_n411_; 
wire alu__abc_42281_new_n412_; 
wire alu__abc_42281_new_n413_; 
wire alu__abc_42281_new_n414_; 
wire alu__abc_42281_new_n415_; 
wire alu__abc_42281_new_n416_; 
wire alu__abc_42281_new_n417_; 
wire alu__abc_42281_new_n418_; 
wire alu__abc_42281_new_n419_; 
wire alu__abc_42281_new_n420_; 
wire alu__abc_42281_new_n421_; 
wire alu__abc_42281_new_n422_; 
wire alu__abc_42281_new_n423_; 
wire alu__abc_42281_new_n424_; 
wire alu__abc_42281_new_n425_; 
wire alu__abc_42281_new_n426_; 
wire alu__abc_42281_new_n427_; 
wire alu__abc_42281_new_n428_; 
wire alu__abc_42281_new_n429_; 
wire alu__abc_42281_new_n430_; 
wire alu__abc_42281_new_n431_; 
wire alu__abc_42281_new_n432_; 
wire alu__abc_42281_new_n433_; 
wire alu__abc_42281_new_n434_; 
wire alu__abc_42281_new_n435_; 
wire alu__abc_42281_new_n436_; 
wire alu__abc_42281_new_n437_; 
wire alu__abc_42281_new_n438_; 
wire alu__abc_42281_new_n439_; 
wire alu__abc_42281_new_n440_; 
wire alu__abc_42281_new_n441_; 
wire alu__abc_42281_new_n442_; 
wire alu__abc_42281_new_n443_; 
wire alu__abc_42281_new_n444_; 
wire alu__abc_42281_new_n445_; 
wire alu__abc_42281_new_n446_; 
wire alu__abc_42281_new_n447_; 
wire alu__abc_42281_new_n448_; 
wire alu__abc_42281_new_n449_; 
wire alu__abc_42281_new_n450_; 
wire alu__abc_42281_new_n451_; 
wire alu__abc_42281_new_n452_; 
wire alu__abc_42281_new_n453_; 
wire alu__abc_42281_new_n454_; 
wire alu__abc_42281_new_n455_; 
wire alu__abc_42281_new_n456_; 
wire alu__abc_42281_new_n457_; 
wire alu__abc_42281_new_n458_; 
wire alu__abc_42281_new_n459_; 
wire alu__abc_42281_new_n460_; 
wire alu__abc_42281_new_n461_; 
wire alu__abc_42281_new_n462_; 
wire alu__abc_42281_new_n463_; 
wire alu__abc_42281_new_n464_; 
wire alu__abc_42281_new_n465_; 
wire alu__abc_42281_new_n466_; 
wire alu__abc_42281_new_n467_; 
wire alu__abc_42281_new_n468_; 
wire alu__abc_42281_new_n469_; 
wire alu__abc_42281_new_n470_; 
wire alu__abc_42281_new_n471_; 
wire alu__abc_42281_new_n472_; 
wire alu__abc_42281_new_n473_; 
wire alu__abc_42281_new_n474_; 
wire alu__abc_42281_new_n475_; 
wire alu__abc_42281_new_n476_; 
wire alu__abc_42281_new_n477_; 
wire alu__abc_42281_new_n478_; 
wire alu__abc_42281_new_n479_; 
wire alu__abc_42281_new_n480_; 
wire alu__abc_42281_new_n481_; 
wire alu__abc_42281_new_n482_; 
wire alu__abc_42281_new_n483_; 
wire alu__abc_42281_new_n484_; 
wire alu__abc_42281_new_n485_; 
wire alu__abc_42281_new_n486_; 
wire alu__abc_42281_new_n487_; 
wire alu__abc_42281_new_n488_; 
wire alu__abc_42281_new_n489_; 
wire alu__abc_42281_new_n490_; 
wire alu__abc_42281_new_n491_; 
wire alu__abc_42281_new_n492_; 
wire alu__abc_42281_new_n493_; 
wire alu__abc_42281_new_n494_; 
wire alu__abc_42281_new_n495_; 
wire alu__abc_42281_new_n496_; 
wire alu__abc_42281_new_n497_; 
wire alu__abc_42281_new_n498_; 
wire alu__abc_42281_new_n499_; 
wire alu__abc_42281_new_n500_; 
wire alu__abc_42281_new_n501_; 
wire alu__abc_42281_new_n502_; 
wire alu__abc_42281_new_n503_; 
wire alu__abc_42281_new_n504_; 
wire alu__abc_42281_new_n505_; 
wire alu__abc_42281_new_n506_; 
wire alu__abc_42281_new_n507_; 
wire alu__abc_42281_new_n508_; 
wire alu__abc_42281_new_n509_; 
wire alu__abc_42281_new_n510_; 
wire alu__abc_42281_new_n512_; 
wire alu__abc_42281_new_n513_; 
wire alu__abc_42281_new_n514_; 
wire alu__abc_42281_new_n515_; 
wire alu__abc_42281_new_n516_; 
wire alu__abc_42281_new_n517_; 
wire alu__abc_42281_new_n518_; 
wire alu__abc_42281_new_n519_; 
wire alu__abc_42281_new_n520_; 
wire alu__abc_42281_new_n521_; 
wire alu__abc_42281_new_n522_; 
wire alu__abc_42281_new_n523_; 
wire alu__abc_42281_new_n524_; 
wire alu__abc_42281_new_n525_; 
wire alu__abc_42281_new_n526_; 
wire alu__abc_42281_new_n527_; 
wire alu__abc_42281_new_n528_; 
wire alu__abc_42281_new_n529_; 
wire alu__abc_42281_new_n530_; 
wire alu__abc_42281_new_n531_; 
wire alu__abc_42281_new_n532_; 
wire alu__abc_42281_new_n533_; 
wire alu__abc_42281_new_n534_; 
wire alu__abc_42281_new_n535_; 
wire alu__abc_42281_new_n536_; 
wire alu__abc_42281_new_n537_; 
wire alu__abc_42281_new_n538_; 
wire alu__abc_42281_new_n539_; 
wire alu__abc_42281_new_n540_; 
wire alu__abc_42281_new_n541_; 
wire alu__abc_42281_new_n542_; 
wire alu__abc_42281_new_n543_; 
wire alu__abc_42281_new_n544_; 
wire alu__abc_42281_new_n545_; 
wire alu__abc_42281_new_n546_; 
wire alu__abc_42281_new_n547_; 
wire alu__abc_42281_new_n548_; 
wire alu__abc_42281_new_n549_; 
wire alu__abc_42281_new_n550_; 
wire alu__abc_42281_new_n551_; 
wire alu__abc_42281_new_n552_; 
wire alu__abc_42281_new_n553_; 
wire alu__abc_42281_new_n554_; 
wire alu__abc_42281_new_n555_; 
wire alu__abc_42281_new_n556_; 
wire alu__abc_42281_new_n557_; 
wire alu__abc_42281_new_n558_; 
wire alu__abc_42281_new_n559_; 
wire alu__abc_42281_new_n560_; 
wire alu__abc_42281_new_n561_; 
wire alu__abc_42281_new_n562_; 
wire alu__abc_42281_new_n563_; 
wire alu__abc_42281_new_n564_; 
wire alu__abc_42281_new_n565_; 
wire alu__abc_42281_new_n566_; 
wire alu__abc_42281_new_n567_; 
wire alu__abc_42281_new_n568_; 
wire alu__abc_42281_new_n569_; 
wire alu__abc_42281_new_n570_; 
wire alu__abc_42281_new_n571_; 
wire alu__abc_42281_new_n572_; 
wire alu__abc_42281_new_n573_; 
wire alu__abc_42281_new_n574_; 
wire alu__abc_42281_new_n575_; 
wire alu__abc_42281_new_n576_; 
wire alu__abc_42281_new_n577_; 
wire alu__abc_42281_new_n578_; 
wire alu__abc_42281_new_n579_; 
wire alu__abc_42281_new_n580_; 
wire alu__abc_42281_new_n581_; 
wire alu__abc_42281_new_n582_; 
wire alu__abc_42281_new_n583_; 
wire alu__abc_42281_new_n584_; 
wire alu__abc_42281_new_n585_; 
wire alu__abc_42281_new_n586_; 
wire alu__abc_42281_new_n587_; 
wire alu__abc_42281_new_n588_; 
wire alu__abc_42281_new_n589_; 
wire alu__abc_42281_new_n590_; 
wire alu__abc_42281_new_n591_; 
wire alu__abc_42281_new_n592_; 
wire alu__abc_42281_new_n593_; 
wire alu__abc_42281_new_n594_; 
wire alu__abc_42281_new_n595_; 
wire alu__abc_42281_new_n596_; 
wire alu__abc_42281_new_n597_; 
wire alu__abc_42281_new_n598_; 
wire alu__abc_42281_new_n599_; 
wire alu__abc_42281_new_n600_; 
wire alu__abc_42281_new_n601_; 
wire alu__abc_42281_new_n602_; 
wire alu__abc_42281_new_n603_; 
wire alu__abc_42281_new_n604_; 
wire alu__abc_42281_new_n605_; 
wire alu__abc_42281_new_n606_; 
wire alu__abc_42281_new_n607_; 
wire alu__abc_42281_new_n608_; 
wire alu__abc_42281_new_n609_; 
wire alu__abc_42281_new_n610_; 
wire alu__abc_42281_new_n611_; 
wire alu__abc_42281_new_n612_; 
wire alu__abc_42281_new_n613_; 
wire alu__abc_42281_new_n614_; 
wire alu__abc_42281_new_n615_; 
wire alu__abc_42281_new_n616_; 
wire alu__abc_42281_new_n617_; 
wire alu__abc_42281_new_n618_; 
wire alu__abc_42281_new_n619_; 
wire alu__abc_42281_new_n620_; 
wire alu__abc_42281_new_n621_; 
wire alu__abc_42281_new_n622_; 
wire alu__abc_42281_new_n623_; 
wire alu__abc_42281_new_n624_; 
wire alu__abc_42281_new_n625_; 
wire alu__abc_42281_new_n626_; 
wire alu__abc_42281_new_n627_; 
wire alu__abc_42281_new_n628_; 
wire alu__abc_42281_new_n629_; 
wire alu__abc_42281_new_n630_; 
wire alu__abc_42281_new_n631_; 
wire alu__abc_42281_new_n632_; 
wire alu__abc_42281_new_n633_; 
wire alu__abc_42281_new_n634_; 
wire alu__abc_42281_new_n635_; 
wire alu__abc_42281_new_n636_; 
wire alu__abc_42281_new_n637_; 
wire alu__abc_42281_new_n638_; 
wire alu__abc_42281_new_n639_; 
wire alu__abc_42281_new_n640_; 
wire alu__abc_42281_new_n641_; 
wire alu__abc_42281_new_n642_; 
wire alu__abc_42281_new_n643_; 
wire alu__abc_42281_new_n644_; 
wire alu__abc_42281_new_n645_; 
wire alu__abc_42281_new_n646_; 
wire alu__abc_42281_new_n647_; 
wire alu__abc_42281_new_n648_; 
wire alu__abc_42281_new_n649_; 
wire alu__abc_42281_new_n650_; 
wire alu__abc_42281_new_n651_; 
wire alu__abc_42281_new_n652_; 
wire alu__abc_42281_new_n653_; 
wire alu__abc_42281_new_n654_; 
wire alu__abc_42281_new_n655_; 
wire alu__abc_42281_new_n656_; 
wire alu__abc_42281_new_n657_; 
wire alu__abc_42281_new_n658_; 
wire alu__abc_42281_new_n659_; 
wire alu__abc_42281_new_n660_; 
wire alu__abc_42281_new_n661_; 
wire alu__abc_42281_new_n662_; 
wire alu__abc_42281_new_n663_; 
wire alu__abc_42281_new_n664_; 
wire alu__abc_42281_new_n665_; 
wire alu__abc_42281_new_n666_; 
wire alu__abc_42281_new_n667_; 
wire alu__abc_42281_new_n668_; 
wire alu__abc_42281_new_n669_; 
wire alu__abc_42281_new_n670_; 
wire alu__abc_42281_new_n671_; 
wire alu__abc_42281_new_n672_; 
wire alu__abc_42281_new_n673_; 
wire alu__abc_42281_new_n674_; 
wire alu__abc_42281_new_n675_; 
wire alu__abc_42281_new_n676_; 
wire alu__abc_42281_new_n677_; 
wire alu__abc_42281_new_n678_; 
wire alu__abc_42281_new_n679_; 
wire alu__abc_42281_new_n680_; 
wire alu__abc_42281_new_n681_; 
wire alu__abc_42281_new_n682_; 
wire alu__abc_42281_new_n683_; 
wire alu__abc_42281_new_n684_; 
wire alu__abc_42281_new_n685_; 
wire alu__abc_42281_new_n686_; 
wire alu__abc_42281_new_n687_; 
wire alu__abc_42281_new_n688_; 
wire alu__abc_42281_new_n689_; 
wire alu__abc_42281_new_n690_; 
wire alu__abc_42281_new_n691_; 
wire alu__abc_42281_new_n692_; 
wire alu__abc_42281_new_n693_; 
wire alu__abc_42281_new_n694_; 
wire alu__abc_42281_new_n695_; 
wire alu__abc_42281_new_n696_; 
wire alu__abc_42281_new_n697_; 
wire alu__abc_42281_new_n698_; 
wire alu__abc_42281_new_n699_; 
wire alu__abc_42281_new_n700_; 
wire alu__abc_42281_new_n701_; 
wire alu__abc_42281_new_n702_; 
wire alu__abc_42281_new_n703_; 
wire alu__abc_42281_new_n704_; 
wire alu__abc_42281_new_n705_; 
wire alu__abc_42281_new_n706_; 
wire alu__abc_42281_new_n707_; 
wire alu__abc_42281_new_n708_; 
wire alu__abc_42281_new_n709_; 
wire alu__abc_42281_new_n710_; 
wire alu__abc_42281_new_n711_; 
wire alu__abc_42281_new_n712_; 
wire alu__abc_42281_new_n713_; 
wire alu__abc_42281_new_n714_; 
wire alu__abc_42281_new_n715_; 
wire alu__abc_42281_new_n716_; 
wire alu__abc_42281_new_n717_; 
wire alu__abc_42281_new_n718_; 
wire alu__abc_42281_new_n719_; 
wire alu__abc_42281_new_n720_; 
wire alu__abc_42281_new_n721_; 
wire alu__abc_42281_new_n722_; 
wire alu__abc_42281_new_n723_; 
wire alu__abc_42281_new_n724_; 
wire alu__abc_42281_new_n725_; 
wire alu__abc_42281_new_n726_; 
wire alu__abc_42281_new_n727_; 
wire alu__abc_42281_new_n728_; 
wire alu__abc_42281_new_n729_; 
wire alu__abc_42281_new_n730_; 
wire alu__abc_42281_new_n731_; 
wire alu__abc_42281_new_n732_; 
wire alu__abc_42281_new_n733_; 
wire alu__abc_42281_new_n734_; 
wire alu__abc_42281_new_n735_; 
wire alu__abc_42281_new_n736_; 
wire alu__abc_42281_new_n737_; 
wire alu__abc_42281_new_n738_; 
wire alu__abc_42281_new_n739_; 
wire alu__abc_42281_new_n740_; 
wire alu__abc_42281_new_n741_; 
wire alu__abc_42281_new_n742_; 
wire alu__abc_42281_new_n743_; 
wire alu__abc_42281_new_n744_; 
wire alu__abc_42281_new_n745_; 
wire alu__abc_42281_new_n746_; 
wire alu__abc_42281_new_n747_; 
wire alu__abc_42281_new_n748_; 
wire alu__abc_42281_new_n749_; 
wire alu__abc_42281_new_n750_; 
wire alu__abc_42281_new_n751_; 
wire alu__abc_42281_new_n752_; 
wire alu__abc_42281_new_n753_; 
wire alu__abc_42281_new_n754_; 
wire alu__abc_42281_new_n755_; 
wire alu__abc_42281_new_n756_; 
wire alu__abc_42281_new_n757_; 
wire alu__abc_42281_new_n758_; 
wire alu__abc_42281_new_n759_; 
wire alu__abc_42281_new_n760_; 
wire alu__abc_42281_new_n761_; 
wire alu__abc_42281_new_n762_; 
wire alu__abc_42281_new_n763_; 
wire alu__abc_42281_new_n764_; 
wire alu__abc_42281_new_n765_; 
wire alu__abc_42281_new_n766_; 
wire alu__abc_42281_new_n767_; 
wire alu__abc_42281_new_n768_; 
wire alu__abc_42281_new_n769_; 
wire alu__abc_42281_new_n770_; 
wire alu__abc_42281_new_n771_; 
wire alu__abc_42281_new_n772_; 
wire alu__abc_42281_new_n773_; 
wire alu__abc_42281_new_n774_; 
wire alu__abc_42281_new_n775_; 
wire alu__abc_42281_new_n776_; 
wire alu__abc_42281_new_n777_; 
wire alu__abc_42281_new_n778_; 
wire alu__abc_42281_new_n779_; 
wire alu__abc_42281_new_n780_; 
wire alu__abc_42281_new_n781_; 
wire alu__abc_42281_new_n782_; 
wire alu__abc_42281_new_n783_; 
wire alu__abc_42281_new_n784_; 
wire alu__abc_42281_new_n785_; 
wire alu__abc_42281_new_n786_; 
wire alu__abc_42281_new_n787_; 
wire alu__abc_42281_new_n788_; 
wire alu__abc_42281_new_n789_; 
wire alu__abc_42281_new_n790_; 
wire alu__abc_42281_new_n791_; 
wire alu__abc_42281_new_n792_; 
wire alu__abc_42281_new_n793_; 
wire alu__abc_42281_new_n794_; 
wire alu__abc_42281_new_n795_; 
wire alu__abc_42281_new_n796_; 
wire alu__abc_42281_new_n797_; 
wire alu__abc_42281_new_n798_; 
wire alu__abc_42281_new_n799_; 
wire alu__abc_42281_new_n800_; 
wire alu__abc_42281_new_n801_; 
wire alu__abc_42281_new_n802_; 
wire alu__abc_42281_new_n803_; 
wire alu__abc_42281_new_n804_; 
wire alu__abc_42281_new_n805_; 
wire alu__abc_42281_new_n806_; 
wire alu__abc_42281_new_n807_; 
wire alu__abc_42281_new_n808_; 
wire alu__abc_42281_new_n809_; 
wire alu__abc_42281_new_n810_; 
wire alu__abc_42281_new_n811_; 
wire alu__abc_42281_new_n812_; 
wire alu__abc_42281_new_n813_; 
wire alu__abc_42281_new_n814_; 
wire alu__abc_42281_new_n815_; 
wire alu__abc_42281_new_n816_; 
wire alu__abc_42281_new_n817_; 
wire alu__abc_42281_new_n818_; 
wire alu__abc_42281_new_n819_; 
wire alu__abc_42281_new_n820_; 
wire alu__abc_42281_new_n821_; 
wire alu__abc_42281_new_n822_; 
wire alu__abc_42281_new_n823_; 
wire alu__abc_42281_new_n824_; 
wire alu__abc_42281_new_n825_; 
wire alu__abc_42281_new_n826_; 
wire alu__abc_42281_new_n827_; 
wire alu__abc_42281_new_n828_; 
wire alu__abc_42281_new_n830_; 
wire alu__abc_42281_new_n831_; 
wire alu__abc_42281_new_n832_; 
wire alu__abc_42281_new_n833_; 
wire alu__abc_42281_new_n834_; 
wire alu__abc_42281_new_n835_; 
wire alu__abc_42281_new_n836_; 
wire alu__abc_42281_new_n837_; 
wire alu__abc_42281_new_n838_; 
wire alu__abc_42281_new_n839_; 
wire alu__abc_42281_new_n840_; 
wire alu__abc_42281_new_n841_; 
wire alu__abc_42281_new_n842_; 
wire alu__abc_42281_new_n843_; 
wire alu__abc_42281_new_n844_; 
wire alu__abc_42281_new_n845_; 
wire alu__abc_42281_new_n846_; 
wire alu__abc_42281_new_n847_; 
wire alu__abc_42281_new_n848_; 
wire alu__abc_42281_new_n849_; 
wire alu__abc_42281_new_n850_; 
wire alu__abc_42281_new_n851_; 
wire alu__abc_42281_new_n852_; 
wire alu__abc_42281_new_n853_; 
wire alu__abc_42281_new_n854_; 
wire alu__abc_42281_new_n855_; 
wire alu__abc_42281_new_n856_; 
wire alu__abc_42281_new_n857_; 
wire alu__abc_42281_new_n858_; 
wire alu__abc_42281_new_n859_; 
wire alu__abc_42281_new_n860_; 
wire alu__abc_42281_new_n861_; 
wire alu__abc_42281_new_n862_; 
wire alu__abc_42281_new_n863_; 
wire alu__abc_42281_new_n864_; 
wire alu__abc_42281_new_n865_; 
wire alu__abc_42281_new_n866_; 
wire alu__abc_42281_new_n867_; 
wire alu__abc_42281_new_n868_; 
wire alu__abc_42281_new_n869_; 
wire alu__abc_42281_new_n870_; 
wire alu__abc_42281_new_n871_; 
wire alu__abc_42281_new_n872_; 
wire alu__abc_42281_new_n873_; 
wire alu__abc_42281_new_n874_; 
wire alu__abc_42281_new_n875_; 
wire alu__abc_42281_new_n876_; 
wire alu__abc_42281_new_n876__bF_buf0; 
wire alu__abc_42281_new_n876__bF_buf1; 
wire alu__abc_42281_new_n876__bF_buf2; 
wire alu__abc_42281_new_n876__bF_buf3; 
wire alu__abc_42281_new_n877_; 
wire alu__abc_42281_new_n878_; 
wire alu__abc_42281_new_n879_; 
wire alu__abc_42281_new_n880_; 
wire alu__abc_42281_new_n881_; 
wire alu__abc_42281_new_n882_; 
wire alu__abc_42281_new_n883_; 
wire alu__abc_42281_new_n884_; 
wire alu__abc_42281_new_n885_; 
wire alu__abc_42281_new_n886_; 
wire alu__abc_42281_new_n887_; 
wire alu__abc_42281_new_n888_; 
wire alu__abc_42281_new_n889_; 
wire alu__abc_42281_new_n890_; 
wire alu__abc_42281_new_n891_; 
wire alu__abc_42281_new_n892_; 
wire alu__abc_42281_new_n893_; 
wire alu__abc_42281_new_n894_; 
wire alu__abc_42281_new_n895_; 
wire alu__abc_42281_new_n896_; 
wire alu__abc_42281_new_n897_; 
wire alu__abc_42281_new_n898_; 
wire alu__abc_42281_new_n899_; 
wire alu__abc_42281_new_n900_; 
wire alu__abc_42281_new_n901_; 
wire alu__abc_42281_new_n902_; 
wire alu__abc_42281_new_n903_; 
wire alu__abc_42281_new_n904_; 
wire alu__abc_42281_new_n905_; 
wire alu__abc_42281_new_n906_; 
wire alu__abc_42281_new_n907_; 
wire alu__abc_42281_new_n908_; 
wire alu__abc_42281_new_n909_; 
wire alu__abc_42281_new_n910_; 
wire alu__abc_42281_new_n911_; 
wire alu__abc_42281_new_n912_; 
wire alu__abc_42281_new_n913_; 
wire alu__abc_42281_new_n914_; 
wire alu__abc_42281_new_n915_; 
wire alu__abc_42281_new_n916_; 
wire alu__abc_42281_new_n917_; 
wire alu__abc_42281_new_n918_; 
wire alu__abc_42281_new_n919_; 
wire alu__abc_42281_new_n920_; 
wire alu__abc_42281_new_n921_; 
wire alu__abc_42281_new_n922_; 
wire alu__abc_42281_new_n923_; 
wire alu__abc_42281_new_n924_; 
wire alu__abc_42281_new_n925_; 
wire alu__abc_42281_new_n926_; 
wire alu__abc_42281_new_n926__bF_buf0; 
wire alu__abc_42281_new_n926__bF_buf1; 
wire alu__abc_42281_new_n926__bF_buf2; 
wire alu__abc_42281_new_n926__bF_buf3; 
wire alu__abc_42281_new_n926__bF_buf4; 
wire alu__abc_42281_new_n927_; 
wire alu__abc_42281_new_n928_; 
wire alu__abc_42281_new_n928__bF_buf0; 
wire alu__abc_42281_new_n928__bF_buf1; 
wire alu__abc_42281_new_n928__bF_buf2; 
wire alu__abc_42281_new_n928__bF_buf3; 
wire alu__abc_42281_new_n928__bF_buf4; 
wire alu__abc_42281_new_n929_; 
wire alu__abc_42281_new_n930_; 
wire alu__abc_42281_new_n931_; 
wire alu__abc_42281_new_n932_; 
wire alu__abc_42281_new_n933_; 
wire alu__abc_42281_new_n934_; 
wire alu__abc_42281_new_n935_; 
wire alu__abc_42281_new_n936_; 
wire alu__abc_42281_new_n936__bF_buf0; 
wire alu__abc_42281_new_n936__bF_buf1; 
wire alu__abc_42281_new_n936__bF_buf2; 
wire alu__abc_42281_new_n936__bF_buf3; 
wire alu__abc_42281_new_n936__bF_buf4; 
wire alu__abc_42281_new_n937_; 
wire alu__abc_42281_new_n938_; 
wire alu__abc_42281_new_n939_; 
wire alu__abc_42281_new_n939__bF_buf0; 
wire alu__abc_42281_new_n939__bF_buf1; 
wire alu__abc_42281_new_n939__bF_buf2; 
wire alu__abc_42281_new_n939__bF_buf3; 
wire alu__abc_42281_new_n939__bF_buf4; 
wire alu__abc_42281_new_n940_; 
wire alu__abc_42281_new_n941_; 
wire alu__abc_42281_new_n941__bF_buf0; 
wire alu__abc_42281_new_n941__bF_buf1; 
wire alu__abc_42281_new_n941__bF_buf2; 
wire alu__abc_42281_new_n941__bF_buf3; 
wire alu__abc_42281_new_n941__bF_buf4; 
wire alu__abc_42281_new_n942_; 
wire alu__abc_42281_new_n942__bF_buf0; 
wire alu__abc_42281_new_n942__bF_buf1; 
wire alu__abc_42281_new_n942__bF_buf2; 
wire alu__abc_42281_new_n942__bF_buf3; 
wire alu__abc_42281_new_n942__bF_buf4; 
wire alu__abc_42281_new_n943_; 
wire alu__abc_42281_new_n944_; 
wire alu__abc_42281_new_n945_; 
wire alu__abc_42281_new_n946_; 
wire alu__abc_42281_new_n947_; 
wire alu__abc_42281_new_n948_; 
wire alu__abc_42281_new_n949_; 
wire alu__abc_42281_new_n950_; 
wire alu__abc_42281_new_n950__bF_buf0; 
wire alu__abc_42281_new_n950__bF_buf1; 
wire alu__abc_42281_new_n950__bF_buf2; 
wire alu__abc_42281_new_n950__bF_buf3; 
wire alu__abc_42281_new_n950__bF_buf4; 
wire alu__abc_42281_new_n951_; 
wire alu__abc_42281_new_n952_; 
wire alu__abc_42281_new_n952__bF_buf0; 
wire alu__abc_42281_new_n952__bF_buf1; 
wire alu__abc_42281_new_n952__bF_buf2; 
wire alu__abc_42281_new_n952__bF_buf3; 
wire alu__abc_42281_new_n952__bF_buf4; 
wire alu__abc_42281_new_n953_; 
wire alu__abc_42281_new_n954_; 
wire alu__abc_42281_new_n955_; 
wire alu__abc_42281_new_n956_; 
wire alu__abc_42281_new_n957_; 
wire alu__abc_42281_new_n958_; 
wire alu__abc_42281_new_n959_; 
wire alu__abc_42281_new_n961_; 
wire alu__abc_42281_new_n962_; 
wire alu__abc_42281_new_n963_; 
wire alu__abc_42281_new_n964_; 
wire alu__abc_42281_new_n965_; 
wire alu__abc_42281_new_n966_; 
wire alu__abc_42281_new_n967_; 
wire alu__abc_42281_new_n968_; 
wire alu__abc_42281_new_n969_; 
wire alu__abc_42281_new_n970_; 
wire alu__abc_42281_new_n971_; 
wire alu__abc_42281_new_n972_; 
wire alu__abc_42281_new_n973_; 
wire alu__abc_42281_new_n974_; 
wire alu__abc_42281_new_n975_; 
wire alu__abc_42281_new_n976_; 
wire alu__abc_42281_new_n977_; 
wire alu__abc_42281_new_n978_; 
wire alu__abc_42281_new_n979_; 
wire alu__abc_42281_new_n980_; 
wire alu__abc_42281_new_n981_; 
wire alu__abc_42281_new_n982_; 
wire alu__abc_42281_new_n983_; 
wire alu__abc_42281_new_n984_; 
wire alu__abc_42281_new_n985_; 
wire alu__abc_42281_new_n986_; 
wire alu__abc_42281_new_n987_; 
wire alu__abc_42281_new_n988_; 
wire alu__abc_42281_new_n989_; 
wire alu__abc_42281_new_n990_; 
wire alu__abc_42281_new_n991_; 
wire alu__abc_42281_new_n992_; 
wire alu__abc_42281_new_n993_; 
wire alu__abc_42281_new_n994_; 
wire alu__abc_42281_new_n995_; 
wire alu__abc_42281_new_n996_; 
wire alu__abc_42281_new_n997_; 
wire alu__abc_42281_new_n998_; 
wire alu__abc_42281_new_n999_; 
wire alu_a_i_0_; 
wire alu_a_i_10_; 
wire alu_a_i_11_; 
wire alu_a_i_12_; 
wire alu_a_i_13_; 
wire alu_a_i_14_; 
wire alu_a_i_15_; 
wire alu_a_i_16_; 
wire alu_a_i_17_; 
wire alu_a_i_18_; 
wire alu_a_i_19_; 
wire alu_a_i_1_; 
wire alu_a_i_20_; 
wire alu_a_i_21_; 
wire alu_a_i_22_; 
wire alu_a_i_23_; 
wire alu_a_i_24_; 
wire alu_a_i_25_; 
wire alu_a_i_26_; 
wire alu_a_i_27_; 
wire alu_a_i_28_; 
wire alu_a_i_29_; 
wire alu_a_i_2_; 
wire alu_a_i_30_; 
wire alu_a_i_31_; 
wire alu_a_i_3_; 
wire alu_a_i_4_; 
wire alu_a_i_5_; 
wire alu_a_i_6_; 
wire alu_a_i_7_; 
wire alu_a_i_8_; 
wire alu_a_i_9_; 
wire alu_b_i_0_; 
wire alu_b_i_0_bF_buf0_; 
wire alu_b_i_0_bF_buf1_; 
wire alu_b_i_0_bF_buf2_; 
wire alu_b_i_0_bF_buf3_; 
wire alu_b_i_0_bF_buf4_; 
wire alu_b_i_10_; 
wire alu_b_i_11_; 
wire alu_b_i_12_; 
wire alu_b_i_13_; 
wire alu_b_i_14_; 
wire alu_b_i_15_; 
wire alu_b_i_16_; 
wire alu_b_i_17_; 
wire alu_b_i_18_; 
wire alu_b_i_19_; 
wire alu_b_i_1_; 
wire alu_b_i_1_bF_buf0_; 
wire alu_b_i_1_bF_buf1_; 
wire alu_b_i_1_bF_buf2_; 
wire alu_b_i_1_bF_buf3_; 
wire alu_b_i_1_bF_buf4_; 
wire alu_b_i_1_bF_buf5_; 
wire alu_b_i_1_bF_buf6_; 
wire alu_b_i_1_bF_buf7_; 
wire alu_b_i_20_; 
wire alu_b_i_21_; 
wire alu_b_i_22_; 
wire alu_b_i_23_; 
wire alu_b_i_24_; 
wire alu_b_i_25_; 
wire alu_b_i_26_; 
wire alu_b_i_27_; 
wire alu_b_i_28_; 
wire alu_b_i_29_; 
wire alu_b_i_2_; 
wire alu_b_i_2_bF_buf0_; 
wire alu_b_i_2_bF_buf1_; 
wire alu_b_i_2_bF_buf2_; 
wire alu_b_i_2_bF_buf3_; 
wire alu_b_i_2_bF_buf4_; 
wire alu_b_i_2_bF_buf5_; 
wire alu_b_i_2_bF_buf6_; 
wire alu_b_i_30_; 
wire alu_b_i_31_; 
wire alu_b_i_3_; 
wire alu_b_i_3_bF_buf0_; 
wire alu_b_i_3_bF_buf1_; 
wire alu_b_i_3_bF_buf2_; 
wire alu_b_i_3_bF_buf3_; 
wire alu_b_i_3_bF_buf4_; 
wire alu_b_i_3_bF_buf5_; 
wire alu_b_i_3_bF_buf6_; 
wire alu_b_i_4_; 
wire alu_b_i_4_bF_buf0_; 
wire alu_b_i_4_bF_buf1_; 
wire alu_b_i_4_bF_buf2_; 
wire alu_b_i_4_bF_buf3_; 
wire alu_b_i_4_bF_buf4_; 
wire alu_b_i_4_bF_buf5_; 
wire alu_b_i_5_; 
wire alu_b_i_6_; 
wire alu_b_i_7_; 
wire alu_b_i_8_; 
wire alu_b_i_9_; 
wire alu_c_i; 
wire alu_c_o; 
wire alu_c_update_o; 
wire alu_equal_o; 
wire alu_flag_update_o; 
wire alu_func_r_0_; 
wire alu_func_r_1_; 
wire alu_func_r_2_; 
wire alu_func_r_3_; 
wire alu_greater_than_o; 
wire alu_greater_than_signed_o; 
wire alu_input_a_r_0_; 
wire alu_input_a_r_10_; 
wire alu_input_a_r_11_; 
wire alu_input_a_r_12_; 
wire alu_input_a_r_13_; 
wire alu_input_a_r_14_; 
wire alu_input_a_r_15_; 
wire alu_input_a_r_16_; 
wire alu_input_a_r_17_; 
wire alu_input_a_r_18_; 
wire alu_input_a_r_19_; 
wire alu_input_a_r_1_; 
wire alu_input_a_r_20_; 
wire alu_input_a_r_21_; 
wire alu_input_a_r_22_; 
wire alu_input_a_r_23_; 
wire alu_input_a_r_24_; 
wire alu_input_a_r_25_; 
wire alu_input_a_r_26_; 
wire alu_input_a_r_27_; 
wire alu_input_a_r_28_; 
wire alu_input_a_r_29_; 
wire alu_input_a_r_2_; 
wire alu_input_a_r_30_; 
wire alu_input_a_r_31_; 
wire alu_input_a_r_3_; 
wire alu_input_a_r_4_; 
wire alu_input_a_r_5_; 
wire alu_input_a_r_6_; 
wire alu_input_a_r_7_; 
wire alu_input_a_r_8_; 
wire alu_input_a_r_9_; 
wire alu_input_b_r_0_; 
wire alu_input_b_r_10_; 
wire alu_input_b_r_11_; 
wire alu_input_b_r_12_; 
wire alu_input_b_r_13_; 
wire alu_input_b_r_14_; 
wire alu_input_b_r_15_; 
wire alu_input_b_r_16_; 
wire alu_input_b_r_17_; 
wire alu_input_b_r_18_; 
wire alu_input_b_r_19_; 
wire alu_input_b_r_1_; 
wire alu_input_b_r_20_; 
wire alu_input_b_r_21_; 
wire alu_input_b_r_22_; 
wire alu_input_b_r_23_; 
wire alu_input_b_r_24_; 
wire alu_input_b_r_25_; 
wire alu_input_b_r_26_; 
wire alu_input_b_r_27_; 
wire alu_input_b_r_28_; 
wire alu_input_b_r_29_; 
wire alu_input_b_r_2_; 
wire alu_input_b_r_30_; 
wire alu_input_b_r_31_; 
wire alu_input_b_r_3_; 
wire alu_input_b_r_4_; 
wire alu_input_b_r_5_; 
wire alu_input_b_r_6_; 
wire alu_input_b_r_7_; 
wire alu_input_b_r_8_; 
wire alu_input_b_r_9_; 
wire alu_less_than_o; 
wire alu_less_than_signed_o; 
wire alu_op_i_0_; 
wire alu_op_i_1_; 
wire alu_op_i_2_; 
wire alu_op_i_3_; 
wire alu_op_r_0_; 
wire alu_op_r_1_; 
wire alu_op_r_2_; 
wire alu_op_r_3_; 
wire alu_op_r_4_; 
wire alu_op_r_5_; 
wire alu_op_r_6_; 
wire alu_op_r_7_; 
wire alu_p_o_0_; 
wire alu_p_o_10_; 
wire alu_p_o_11_; 
wire alu_p_o_12_; 
wire alu_p_o_13_; 
wire alu_p_o_14_; 
wire alu_p_o_15_; 
wire alu_p_o_16_; 
wire alu_p_o_17_; 
wire alu_p_o_18_; 
wire alu_p_o_19_; 
wire alu_p_o_1_; 
wire alu_p_o_20_; 
wire alu_p_o_21_; 
wire alu_p_o_22_; 
wire alu_p_o_23_; 
wire alu_p_o_24_; 
wire alu_p_o_25_; 
wire alu_p_o_26_; 
wire alu_p_o_27_; 
wire alu_p_o_28_; 
wire alu_p_o_29_; 
wire alu_p_o_2_; 
wire alu_p_o_30_; 
wire alu_p_o_31_; 
wire alu_p_o_3_; 
wire alu_p_o_4_; 
wire alu_p_o_5_; 
wire alu_p_o_6_; 
wire alu_p_o_7_; 
wire alu_p_o_8_; 
wire alu_p_o_9_; 
output break_o;
input clk_i;
wire clk_i_bF_buf0; 
wire clk_i_bF_buf1; 
wire clk_i_bF_buf10; 
wire clk_i_bF_buf100; 
wire clk_i_bF_buf101; 
wire clk_i_bF_buf102; 
wire clk_i_bF_buf103; 
wire clk_i_bF_buf104; 
wire clk_i_bF_buf105; 
wire clk_i_bF_buf106; 
wire clk_i_bF_buf107; 
wire clk_i_bF_buf108; 
wire clk_i_bF_buf109; 
wire clk_i_bF_buf11; 
wire clk_i_bF_buf110; 
wire clk_i_bF_buf111; 
wire clk_i_bF_buf112; 
wire clk_i_bF_buf113; 
wire clk_i_bF_buf114; 
wire clk_i_bF_buf12; 
wire clk_i_bF_buf13; 
wire clk_i_bF_buf14; 
wire clk_i_bF_buf15; 
wire clk_i_bF_buf16; 
wire clk_i_bF_buf17; 
wire clk_i_bF_buf18; 
wire clk_i_bF_buf19; 
wire clk_i_bF_buf2; 
wire clk_i_bF_buf20; 
wire clk_i_bF_buf21; 
wire clk_i_bF_buf22; 
wire clk_i_bF_buf23; 
wire clk_i_bF_buf24; 
wire clk_i_bF_buf25; 
wire clk_i_bF_buf26; 
wire clk_i_bF_buf27; 
wire clk_i_bF_buf28; 
wire clk_i_bF_buf29; 
wire clk_i_bF_buf3; 
wire clk_i_bF_buf30; 
wire clk_i_bF_buf31; 
wire clk_i_bF_buf32; 
wire clk_i_bF_buf33; 
wire clk_i_bF_buf34; 
wire clk_i_bF_buf35; 
wire clk_i_bF_buf36; 
wire clk_i_bF_buf37; 
wire clk_i_bF_buf38; 
wire clk_i_bF_buf39; 
wire clk_i_bF_buf4; 
wire clk_i_bF_buf40; 
wire clk_i_bF_buf41; 
wire clk_i_bF_buf42; 
wire clk_i_bF_buf43; 
wire clk_i_bF_buf44; 
wire clk_i_bF_buf45; 
wire clk_i_bF_buf46; 
wire clk_i_bF_buf47; 
wire clk_i_bF_buf48; 
wire clk_i_bF_buf49; 
wire clk_i_bF_buf5; 
wire clk_i_bF_buf50; 
wire clk_i_bF_buf51; 
wire clk_i_bF_buf52; 
wire clk_i_bF_buf53; 
wire clk_i_bF_buf54; 
wire clk_i_bF_buf55; 
wire clk_i_bF_buf56; 
wire clk_i_bF_buf57; 
wire clk_i_bF_buf58; 
wire clk_i_bF_buf59; 
wire clk_i_bF_buf6; 
wire clk_i_bF_buf60; 
wire clk_i_bF_buf61; 
wire clk_i_bF_buf62; 
wire clk_i_bF_buf63; 
wire clk_i_bF_buf64; 
wire clk_i_bF_buf65; 
wire clk_i_bF_buf66; 
wire clk_i_bF_buf67; 
wire clk_i_bF_buf68; 
wire clk_i_bF_buf69; 
wire clk_i_bF_buf7; 
wire clk_i_bF_buf70; 
wire clk_i_bF_buf71; 
wire clk_i_bF_buf72; 
wire clk_i_bF_buf73; 
wire clk_i_bF_buf74; 
wire clk_i_bF_buf75; 
wire clk_i_bF_buf76; 
wire clk_i_bF_buf77; 
wire clk_i_bF_buf78; 
wire clk_i_bF_buf79; 
wire clk_i_bF_buf8; 
wire clk_i_bF_buf80; 
wire clk_i_bF_buf81; 
wire clk_i_bF_buf82; 
wire clk_i_bF_buf83; 
wire clk_i_bF_buf84; 
wire clk_i_bF_buf85; 
wire clk_i_bF_buf86; 
wire clk_i_bF_buf87; 
wire clk_i_bF_buf88; 
wire clk_i_bF_buf89; 
wire clk_i_bF_buf9; 
wire clk_i_bF_buf90; 
wire clk_i_bF_buf91; 
wire clk_i_bF_buf92; 
wire clk_i_bF_buf93; 
wire clk_i_bF_buf94; 
wire clk_i_bF_buf95; 
wire clk_i_bF_buf96; 
wire clk_i_bF_buf97; 
wire clk_i_bF_buf98; 
wire clk_i_bF_buf99; 
wire clk_i_hier0_bF_buf0; 
wire clk_i_hier0_bF_buf1; 
wire clk_i_hier0_bF_buf2; 
wire clk_i_hier0_bF_buf3; 
wire clk_i_hier0_bF_buf4; 
wire clk_i_hier0_bF_buf5; 
wire clk_i_hier0_bF_buf6; 
wire clk_i_hier0_bF_buf7; 
wire clk_i_hier0_bF_buf8; 
wire clk_i_hier0_bF_buf9; 
input enable_i;
wire enable_i_bF_buf0; 
wire enable_i_bF_buf1; 
wire enable_i_bF_buf2; 
wire enable_i_bF_buf3; 
wire enable_i_bF_buf4; 
wire enable_i_bF_buf5; 
wire enable_i_bF_buf6; 
wire enable_i_bF_buf7; 
wire epc_q_0_; 
wire epc_q_10_; 
wire epc_q_11_; 
wire epc_q_12_; 
wire epc_q_13_; 
wire epc_q_14_; 
wire epc_q_15_; 
wire epc_q_16_; 
wire epc_q_17_; 
wire epc_q_18_; 
wire epc_q_19_; 
wire epc_q_1_; 
wire epc_q_20_; 
wire epc_q_21_; 
wire epc_q_22_; 
wire epc_q_23_; 
wire epc_q_24_; 
wire epc_q_25_; 
wire epc_q_26_; 
wire epc_q_27_; 
wire epc_q_28_; 
wire epc_q_29_; 
wire epc_q_2_; 
wire epc_q_30_; 
wire epc_q_31_; 
wire epc_q_3_; 
wire epc_q_4_; 
wire epc_q_5_; 
wire epc_q_6_; 
wire epc_q_7_; 
wire epc_q_8_; 
wire epc_q_9_; 
wire esr_q_10_; 
wire esr_q_2_; 
wire esr_q_9_; 
output fault_o;
wire inst_r_0_; 
wire inst_r_1_; 
wire inst_r_2_; 
wire inst_r_3_; 
wire inst_r_4_; 
wire inst_r_5_; 
wire inst_trap_w; 
wire int32_r_10_; 
wire int32_r_4_; 
wire int32_r_5_; 
input intr_i;
input mem_ack_i;
output \mem_addr_o[0] ;
output \mem_addr_o[10] ;
output \mem_addr_o[11] ;
output \mem_addr_o[12] ;
output \mem_addr_o[13] ;
output \mem_addr_o[14] ;
output \mem_addr_o[15] ;
output \mem_addr_o[16] ;
output \mem_addr_o[17] ;
output \mem_addr_o[18] ;
output \mem_addr_o[19] ;
output \mem_addr_o[1] ;
output \mem_addr_o[20] ;
output \mem_addr_o[21] ;
output \mem_addr_o[22] ;
output \mem_addr_o[23] ;
output \mem_addr_o[24] ;
output \mem_addr_o[25] ;
output \mem_addr_o[26] ;
output \mem_addr_o[27] ;
output \mem_addr_o[28] ;
output \mem_addr_o[29] ;
output \mem_addr_o[2] ;
output \mem_addr_o[30] ;
output \mem_addr_o[31] ;
output \mem_addr_o[3] ;
output \mem_addr_o[4] ;
output \mem_addr_o[5] ;
output \mem_addr_o[6] ;
output \mem_addr_o[7] ;
output \mem_addr_o[8] ;
output \mem_addr_o[9] ;
output \mem_cti_o[0] ;
output \mem_cti_o[1] ;
output \mem_cti_o[2] ;
output mem_cyc_o;
input \mem_dat_i[0] ;
input \mem_dat_i[10] ;
input \mem_dat_i[11] ;
input \mem_dat_i[12] ;
input \mem_dat_i[13] ;
input \mem_dat_i[14] ;
input \mem_dat_i[15] ;
input \mem_dat_i[16] ;
input \mem_dat_i[17] ;
input \mem_dat_i[18] ;
input \mem_dat_i[19] ;
input \mem_dat_i[1] ;
input \mem_dat_i[20] ;
input \mem_dat_i[21] ;
input \mem_dat_i[22] ;
input \mem_dat_i[23] ;
input \mem_dat_i[24] ;
input \mem_dat_i[25] ;
input \mem_dat_i[26] ;
input \mem_dat_i[27] ;
input \mem_dat_i[28] ;
input \mem_dat_i[29] ;
input \mem_dat_i[2] ;
input \mem_dat_i[30] ;
input \mem_dat_i[31] ;
input \mem_dat_i[3] ;
input \mem_dat_i[4] ;
input \mem_dat_i[5] ;
input \mem_dat_i[6] ;
input \mem_dat_i[7] ;
input \mem_dat_i[8] ;
input \mem_dat_i[9] ;
output \mem_dat_o[0] ;
output \mem_dat_o[10] ;
output \mem_dat_o[11] ;
output \mem_dat_o[12] ;
output \mem_dat_o[13] ;
output \mem_dat_o[14] ;
output \mem_dat_o[15] ;
output \mem_dat_o[16] ;
output \mem_dat_o[17] ;
output \mem_dat_o[18] ;
output \mem_dat_o[19] ;
output \mem_dat_o[1] ;
output \mem_dat_o[20] ;
output \mem_dat_o[21] ;
output \mem_dat_o[22] ;
output \mem_dat_o[23] ;
output \mem_dat_o[24] ;
output \mem_dat_o[25] ;
output \mem_dat_o[26] ;
output \mem_dat_o[27] ;
output \mem_dat_o[28] ;
output \mem_dat_o[29] ;
output \mem_dat_o[2] ;
output \mem_dat_o[30] ;
output \mem_dat_o[31] ;
output \mem_dat_o[3] ;
output \mem_dat_o[4] ;
output \mem_dat_o[5] ;
output \mem_dat_o[6] ;
output \mem_dat_o[7] ;
output \mem_dat_o[8] ;
output \mem_dat_o[9] ;
wire mem_offset_q_0_; 
wire mem_offset_q_1_; 
output \mem_sel_o[0] ;
output \mem_sel_o[1] ;
output \mem_sel_o[2] ;
output \mem_sel_o[3] ;
input mem_stall_i;
output mem_stb_o;
output mem_we_o;
wire next_pc_r_0_; 
wire next_pc_r_1_; 
input nmi_i;
wire nmi_q; 
wire opcode_q_21_; 
wire opcode_q_22_; 
wire opcode_q_23_; 
wire opcode_q_24_; 
wire opcode_q_25_; 
wire pc_q_10_; 
wire pc_q_11_; 
wire pc_q_12_; 
wire pc_q_13_; 
wire pc_q_14_; 
wire pc_q_15_; 
wire pc_q_16_; 
wire pc_q_17_; 
wire pc_q_18_; 
wire pc_q_19_; 
wire pc_q_20_; 
wire pc_q_21_; 
wire pc_q_22_; 
wire pc_q_23_; 
wire pc_q_24_; 
wire pc_q_25_; 
wire pc_q_26_; 
wire pc_q_27_; 
wire pc_q_28_; 
wire pc_q_29_; 
wire pc_q_2_; 
wire pc_q_30_; 
wire pc_q_31_; 
wire pc_q_3_; 
wire pc_q_4_; 
wire pc_q_5_; 
wire pc_q_6_; 
wire pc_q_7_; 
wire pc_q_8_; 
wire pc_q_9_; 
input rst_i;
wire sr_q_2_; 
wire sr_q_9_; 
wire state_q_0_; 
wire state_q_1_; 
wire state_q_1_bF_buf0_; 
wire state_q_1_bF_buf1_; 
wire state_q_1_bF_buf2_; 
wire state_q_1_bF_buf3_; 
wire state_q_1_bF_buf4_; 
wire state_q_2_; 
wire state_q_3_; 
wire state_q_3_bF_buf0_; 
wire state_q_3_bF_buf1_; 
wire state_q_3_bF_buf2_; 
wire state_q_3_bF_buf3_; 
wire state_q_3_bF_buf4_; 
wire state_q_3_bF_buf5_; 
wire state_q_4_; 
wire state_q_5_; 
wire state_q_5_bF_buf0_; 
wire state_q_5_bF_buf1_; 
wire state_q_5_bF_buf2_; 
wire state_q_5_bF_buf3_; 
AND2X2 AND2X2_1 ( .A(_abc_44694_new_n617_), .B(_abc_44694_new_n618_), .Y(_abc_44694_new_n619_));
AND2X2 AND2X2_10 ( .A(_abc_44694_new_n632_), .B(_abc_44694_new_n633_), .Y(_abc_44694_new_n634_));
AND2X2 AND2X2_100 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[30] ), .Y(_abc_44694_new_n787_));
AND2X2 AND2X2_1000 ( .A(_abc_44694_new_n1522__bF_buf4), .B(epc_q_30_), .Y(_abc_44694_new_n2501_));
AND2X2 AND2X2_1001 ( .A(_abc_44694_new_n1348__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_44694_new_n2502_));
AND2X2 AND2X2_1002 ( .A(_abc_44694_new_n1207__bF_buf1), .B(_abc_44694_new_n2504_), .Y(_abc_44694_new_n2505_));
AND2X2 AND2X2_1003 ( .A(_abc_44694_new_n2500_), .B(_abc_44694_new_n2505_), .Y(_abc_44694_new_n2506_));
AND2X2 AND2X2_1004 ( .A(_abc_44694_new_n2508_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n2509_));
AND2X2 AND2X2_1005 ( .A(_abc_44694_new_n2507_), .B(_abc_44694_new_n2509_), .Y(_0epc_q_31_0__30_));
AND2X2 AND2X2_1006 ( .A(_abc_44694_new_n2471_), .B(pc_q_31_), .Y(_abc_44694_new_n2512_));
AND2X2 AND2X2_1007 ( .A(_abc_44694_new_n2513_), .B(_abc_44694_new_n2511_), .Y(_abc_44694_new_n2514_));
AND2X2 AND2X2_1008 ( .A(_abc_44694_new_n2514_), .B(_abc_44694_new_n1382__bF_buf2), .Y(_abc_44694_new_n2515_));
AND2X2 AND2X2_1009 ( .A(_abc_44694_new_n2479_), .B(_abc_44694_new_n2485_), .Y(_abc_44694_new_n2518_));
AND2X2 AND2X2_101 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[22] ), .Y(_abc_44694_new_n788_));
AND2X2 AND2X2_1010 ( .A(_abc_44694_new_n2519_), .B(_abc_44694_new_n2520_), .Y(_abc_44694_new_n2521_));
AND2X2 AND2X2_1011 ( .A(_abc_44694_new_n2524_), .B(_abc_44694_new_n1194__bF_buf3), .Y(_abc_44694_new_n2525_));
AND2X2 AND2X2_1012 ( .A(_abc_44694_new_n2525_), .B(_abc_44694_new_n2523_), .Y(_abc_44694_new_n2526_));
AND2X2 AND2X2_1013 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_31_), .Y(_abc_44694_new_n2527_));
AND2X2 AND2X2_1014 ( .A(_abc_44694_new_n2529_), .B(_abc_44694_new_n2530_), .Y(_abc_44694_new_n2531_));
AND2X2 AND2X2_1015 ( .A(_abc_44694_new_n2533_), .B(_abc_44694_new_n2532_), .Y(_abc_44694_new_n2534_));
AND2X2 AND2X2_1016 ( .A(_abc_44694_new_n1522__bF_buf3), .B(epc_q_31_), .Y(_abc_44694_new_n2536_));
AND2X2 AND2X2_1017 ( .A(_abc_44694_new_n1348__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_44694_new_n2537_));
AND2X2 AND2X2_1018 ( .A(_abc_44694_new_n1207__bF_buf0), .B(_abc_44694_new_n2539_), .Y(_abc_44694_new_n2540_));
AND2X2 AND2X2_1019 ( .A(_abc_44694_new_n2535_), .B(_abc_44694_new_n2540_), .Y(_abc_44694_new_n2541_));
AND2X2 AND2X2_102 ( .A(_abc_44694_new_n791_), .B(state_q_1_bF_buf0_), .Y(_abc_44694_new_n792_));
AND2X2 AND2X2_1020 ( .A(_abc_44694_new_n2543_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n2544_));
AND2X2 AND2X2_1021 ( .A(_abc_44694_new_n2542_), .B(_abc_44694_new_n2544_), .Y(_0epc_q_31_0__31_));
AND2X2 AND2X2_1022 ( .A(_abc_44694_new_n1206_), .B(_abc_44694_new_n1278__bF_buf0), .Y(_abc_44694_new_n2546_));
AND2X2 AND2X2_1023 ( .A(_abc_44694_new_n2546__bF_buf4), .B(_abc_44694_new_n1342_), .Y(_abc_44694_new_n2547_));
AND2X2 AND2X2_1024 ( .A(_abc_44694_new_n2549_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n2550_));
AND2X2 AND2X2_1025 ( .A(_abc_44694_new_n2548_), .B(_abc_44694_new_n2550_), .Y(_0pc_q_31_0__0_));
AND2X2 AND2X2_1026 ( .A(_abc_44694_new_n2546__bF_buf3), .B(_abc_44694_new_n1367_), .Y(_abc_44694_new_n2552_));
AND2X2 AND2X2_1027 ( .A(_abc_44694_new_n2554_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n2555_));
AND2X2 AND2X2_1028 ( .A(_abc_44694_new_n2553_), .B(_abc_44694_new_n2555_), .Y(_0pc_q_31_0__1_));
AND2X2 AND2X2_1029 ( .A(_abc_44694_new_n2546__bF_buf2), .B(_abc_44694_new_n1414_), .Y(_abc_44694_new_n2557_));
AND2X2 AND2X2_103 ( .A(_abc_44694_new_n783_), .B(_abc_44694_new_n792_), .Y(_abc_44694_new_n793_));
AND2X2 AND2X2_1030 ( .A(_abc_44694_new_n2559_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n2560_));
AND2X2 AND2X2_1031 ( .A(_abc_44694_new_n2558_), .B(_abc_44694_new_n2560_), .Y(_0pc_q_31_0__2_));
AND2X2 AND2X2_1032 ( .A(_abc_44694_new_n2546__bF_buf1), .B(_abc_44694_new_n1450_), .Y(_abc_44694_new_n2562_));
AND2X2 AND2X2_1033 ( .A(_abc_44694_new_n2564_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n2565_));
AND2X2 AND2X2_1034 ( .A(_abc_44694_new_n2563_), .B(_abc_44694_new_n2565_), .Y(_0pc_q_31_0__3_));
AND2X2 AND2X2_1035 ( .A(_abc_44694_new_n2546__bF_buf0), .B(_abc_44694_new_n1488_), .Y(_abc_44694_new_n2567_));
AND2X2 AND2X2_1036 ( .A(_abc_44694_new_n2569_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n2570_));
AND2X2 AND2X2_1037 ( .A(_abc_44694_new_n2568_), .B(_abc_44694_new_n2570_), .Y(_0pc_q_31_0__4_));
AND2X2 AND2X2_1038 ( .A(_abc_44694_new_n2546__bF_buf4), .B(_abc_44694_new_n1520_), .Y(_abc_44694_new_n2572_));
AND2X2 AND2X2_1039 ( .A(_abc_44694_new_n2574_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n2575_));
AND2X2 AND2X2_104 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[31] ), .Y(_abc_44694_new_n795_));
AND2X2 AND2X2_1040 ( .A(_abc_44694_new_n2573_), .B(_abc_44694_new_n2575_), .Y(_0pc_q_31_0__5_));
AND2X2 AND2X2_1041 ( .A(_abc_44694_new_n2546__bF_buf3), .B(_abc_44694_new_n1563_), .Y(_abc_44694_new_n2577_));
AND2X2 AND2X2_1042 ( .A(_abc_44694_new_n2579_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n2580_));
AND2X2 AND2X2_1043 ( .A(_abc_44694_new_n2578_), .B(_abc_44694_new_n2580_), .Y(_0pc_q_31_0__6_));
AND2X2 AND2X2_1044 ( .A(_abc_44694_new_n2546__bF_buf2), .B(_abc_44694_new_n1602_), .Y(_abc_44694_new_n2582_));
AND2X2 AND2X2_1045 ( .A(_abc_44694_new_n2584_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n2585_));
AND2X2 AND2X2_1046 ( .A(_abc_44694_new_n2583_), .B(_abc_44694_new_n2585_), .Y(_0pc_q_31_0__7_));
AND2X2 AND2X2_1047 ( .A(_abc_44694_new_n2587_), .B(_abc_44694_new_n1330_), .Y(_abc_44694_new_n2588_));
AND2X2 AND2X2_1048 ( .A(_abc_44694_new_n1210__bF_buf1), .B(pc_q_8_), .Y(_abc_44694_new_n2589_));
AND2X2 AND2X2_1049 ( .A(_abc_44694_new_n2592_), .B(_abc_44694_new_n1659_), .Y(_abc_44694_new_n2593_));
AND2X2 AND2X2_105 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[15] ), .Y(_abc_44694_new_n796_));
AND2X2 AND2X2_1050 ( .A(_abc_44694_new_n2593_), .B(_abc_44694_new_n1206_), .Y(_abc_44694_new_n2594_));
AND2X2 AND2X2_1051 ( .A(_abc_44694_new_n2597_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n2598_));
AND2X2 AND2X2_1052 ( .A(_abc_44694_new_n2596_), .B(_abc_44694_new_n2598_), .Y(_0pc_q_31_0__9_));
AND2X2 AND2X2_1053 ( .A(_abc_44694_new_n1719_), .B(_abc_44694_new_n1277_), .Y(_abc_44694_new_n2601_));
AND2X2 AND2X2_1054 ( .A(_abc_44694_new_n2603_), .B(_abc_44694_new_n1206_), .Y(_abc_44694_new_n2604_));
AND2X2 AND2X2_1055 ( .A(_abc_44694_new_n2605_), .B(_abc_44694_new_n2600_), .Y(_abc_44694_new_n2606_));
AND2X2 AND2X2_1056 ( .A(_abc_44694_new_n2606_), .B(enable_i_bF_buf6), .Y(_0pc_q_31_0__10_));
AND2X2 AND2X2_1057 ( .A(_abc_44694_new_n1755_), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n2609_));
AND2X2 AND2X2_1058 ( .A(_abc_44694_new_n2610_), .B(_abc_44694_new_n2608_), .Y(_abc_44694_new_n2611_));
AND2X2 AND2X2_1059 ( .A(_abc_44694_new_n2613_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n2614_));
AND2X2 AND2X2_106 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[23] ), .Y(_abc_44694_new_n798_));
AND2X2 AND2X2_1060 ( .A(_abc_44694_new_n2612_), .B(_abc_44694_new_n2614_), .Y(_0pc_q_31_0__11_));
AND2X2 AND2X2_1061 ( .A(_abc_44694_new_n1797_), .B(_abc_44694_new_n2546__bF_buf1), .Y(_abc_44694_new_n2616_));
AND2X2 AND2X2_1062 ( .A(_abc_44694_new_n2618_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n2619_));
AND2X2 AND2X2_1063 ( .A(_abc_44694_new_n2617_), .B(_abc_44694_new_n2619_), .Y(_0pc_q_31_0__12_));
AND2X2 AND2X2_1064 ( .A(_abc_44694_new_n1836_), .B(_abc_44694_new_n2546__bF_buf0), .Y(_abc_44694_new_n2621_));
AND2X2 AND2X2_1065 ( .A(_abc_44694_new_n2623_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n2624_));
AND2X2 AND2X2_1066 ( .A(_abc_44694_new_n2622_), .B(_abc_44694_new_n2624_), .Y(_0pc_q_31_0__13_));
AND2X2 AND2X2_1067 ( .A(_abc_44694_new_n1873_), .B(_abc_44694_new_n2546__bF_buf4), .Y(_abc_44694_new_n2626_));
AND2X2 AND2X2_1068 ( .A(_abc_44694_new_n2628_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n2629_));
AND2X2 AND2X2_1069 ( .A(_abc_44694_new_n2627_), .B(_abc_44694_new_n2629_), .Y(_0pc_q_31_0__14_));
AND2X2 AND2X2_107 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[7] ), .Y(_abc_44694_new_n799_));
AND2X2 AND2X2_1070 ( .A(_abc_44694_new_n1909_), .B(_abc_44694_new_n2546__bF_buf3), .Y(_abc_44694_new_n2631_));
AND2X2 AND2X2_1071 ( .A(_abc_44694_new_n2633_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n2634_));
AND2X2 AND2X2_1072 ( .A(_abc_44694_new_n2632_), .B(_abc_44694_new_n2634_), .Y(_0pc_q_31_0__15_));
AND2X2 AND2X2_1073 ( .A(_abc_44694_new_n1955_), .B(_abc_44694_new_n2546__bF_buf2), .Y(_abc_44694_new_n2636_));
AND2X2 AND2X2_1074 ( .A(_abc_44694_new_n2638_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n2639_));
AND2X2 AND2X2_1075 ( .A(_abc_44694_new_n2637_), .B(_abc_44694_new_n2639_), .Y(_0pc_q_31_0__16_));
AND2X2 AND2X2_1076 ( .A(_abc_44694_new_n1991_), .B(_abc_44694_new_n2546__bF_buf1), .Y(_abc_44694_new_n2641_));
AND2X2 AND2X2_1077 ( .A(_abc_44694_new_n2643_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n2644_));
AND2X2 AND2X2_1078 ( .A(_abc_44694_new_n2642_), .B(_abc_44694_new_n2644_), .Y(_0pc_q_31_0__17_));
AND2X2 AND2X2_1079 ( .A(_abc_44694_new_n2027_), .B(_abc_44694_new_n2546__bF_buf0), .Y(_abc_44694_new_n2646_));
AND2X2 AND2X2_108 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[23] ), .Y(_abc_44694_new_n803_));
AND2X2 AND2X2_1080 ( .A(_abc_44694_new_n2648_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n2649_));
AND2X2 AND2X2_1081 ( .A(_abc_44694_new_n2647_), .B(_abc_44694_new_n2649_), .Y(_0pc_q_31_0__18_));
AND2X2 AND2X2_1082 ( .A(_abc_44694_new_n2063_), .B(_abc_44694_new_n2546__bF_buf4), .Y(_abc_44694_new_n2651_));
AND2X2 AND2X2_1083 ( .A(_abc_44694_new_n2653_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n2654_));
AND2X2 AND2X2_1084 ( .A(_abc_44694_new_n2652_), .B(_abc_44694_new_n2654_), .Y(_0pc_q_31_0__19_));
AND2X2 AND2X2_1085 ( .A(_abc_44694_new_n2112_), .B(_abc_44694_new_n2546__bF_buf3), .Y(_abc_44694_new_n2656_));
AND2X2 AND2X2_1086 ( .A(_abc_44694_new_n2658_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n2659_));
AND2X2 AND2X2_1087 ( .A(_abc_44694_new_n2657_), .B(_abc_44694_new_n2659_), .Y(_0pc_q_31_0__20_));
AND2X2 AND2X2_1088 ( .A(_abc_44694_new_n2151_), .B(_abc_44694_new_n2546__bF_buf2), .Y(_abc_44694_new_n2661_));
AND2X2 AND2X2_1089 ( .A(_abc_44694_new_n2663_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n2664_));
AND2X2 AND2X2_109 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[7] ), .Y(_abc_44694_new_n804_));
AND2X2 AND2X2_1090 ( .A(_abc_44694_new_n2662_), .B(_abc_44694_new_n2664_), .Y(_0pc_q_31_0__21_));
AND2X2 AND2X2_1091 ( .A(_abc_44694_new_n2188_), .B(_abc_44694_new_n2546__bF_buf1), .Y(_abc_44694_new_n2666_));
AND2X2 AND2X2_1092 ( .A(_abc_44694_new_n2668_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n2669_));
AND2X2 AND2X2_1093 ( .A(_abc_44694_new_n2667_), .B(_abc_44694_new_n2669_), .Y(_0pc_q_31_0__22_));
AND2X2 AND2X2_1094 ( .A(_abc_44694_new_n2224_), .B(_abc_44694_new_n2546__bF_buf0), .Y(_abc_44694_new_n2671_));
AND2X2 AND2X2_1095 ( .A(_abc_44694_new_n2673_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n2674_));
AND2X2 AND2X2_1096 ( .A(_abc_44694_new_n2672_), .B(_abc_44694_new_n2674_), .Y(_0pc_q_31_0__23_));
AND2X2 AND2X2_1097 ( .A(_abc_44694_new_n2270_), .B(_abc_44694_new_n2546__bF_buf4), .Y(_abc_44694_new_n2676_));
AND2X2 AND2X2_1098 ( .A(_abc_44694_new_n2678_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n2679_));
AND2X2 AND2X2_1099 ( .A(_abc_44694_new_n2677_), .B(_abc_44694_new_n2679_), .Y(_0pc_q_31_0__24_));
AND2X2 AND2X2_11 ( .A(_abc_44694_new_n634_), .B(_abc_44694_new_n630_), .Y(_abc_44694_new_n635_));
AND2X2 AND2X2_110 ( .A(_abc_44694_new_n806_), .B(_abc_44694_new_n802_), .Y(_abc_44694_new_n807_));
AND2X2 AND2X2_1100 ( .A(_abc_44694_new_n2309_), .B(_abc_44694_new_n2546__bF_buf3), .Y(_abc_44694_new_n2681_));
AND2X2 AND2X2_1101 ( .A(_abc_44694_new_n2683_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n2684_));
AND2X2 AND2X2_1102 ( .A(_abc_44694_new_n2682_), .B(_abc_44694_new_n2684_), .Y(_0pc_q_31_0__25_));
AND2X2 AND2X2_1103 ( .A(_abc_44694_new_n2346_), .B(_abc_44694_new_n2546__bF_buf2), .Y(_abc_44694_new_n2686_));
AND2X2 AND2X2_1104 ( .A(_abc_44694_new_n2688_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n2689_));
AND2X2 AND2X2_1105 ( .A(_abc_44694_new_n2687_), .B(_abc_44694_new_n2689_), .Y(_0pc_q_31_0__26_));
AND2X2 AND2X2_1106 ( .A(_abc_44694_new_n2385_), .B(_abc_44694_new_n2546__bF_buf1), .Y(_abc_44694_new_n2691_));
AND2X2 AND2X2_1107 ( .A(_abc_44694_new_n2693_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n2694_));
AND2X2 AND2X2_1108 ( .A(_abc_44694_new_n2692_), .B(_abc_44694_new_n2694_), .Y(_0pc_q_31_0__27_));
AND2X2 AND2X2_1109 ( .A(_abc_44694_new_n2422_), .B(_abc_44694_new_n2546__bF_buf0), .Y(_abc_44694_new_n2696_));
AND2X2 AND2X2_111 ( .A(_abc_44694_new_n808_), .B(_abc_44694_new_n809_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_));
AND2X2 AND2X2_1110 ( .A(_abc_44694_new_n2698_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n2699_));
AND2X2 AND2X2_1111 ( .A(_abc_44694_new_n2697_), .B(_abc_44694_new_n2699_), .Y(_0pc_q_31_0__28_));
AND2X2 AND2X2_1112 ( .A(_abc_44694_new_n2458_), .B(_abc_44694_new_n2546__bF_buf4), .Y(_abc_44694_new_n2701_));
AND2X2 AND2X2_1113 ( .A(_abc_44694_new_n2703_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n2704_));
AND2X2 AND2X2_1114 ( .A(_abc_44694_new_n2702_), .B(_abc_44694_new_n2704_), .Y(_0pc_q_31_0__29_));
AND2X2 AND2X2_1115 ( .A(_abc_44694_new_n2499_), .B(_abc_44694_new_n2546__bF_buf3), .Y(_abc_44694_new_n2706_));
AND2X2 AND2X2_1116 ( .A(_abc_44694_new_n2708_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n2709_));
AND2X2 AND2X2_1117 ( .A(_abc_44694_new_n2707_), .B(_abc_44694_new_n2709_), .Y(_0pc_q_31_0__30_));
AND2X2 AND2X2_1118 ( .A(_abc_44694_new_n2534_), .B(_abc_44694_new_n2546__bF_buf2), .Y(_abc_44694_new_n2711_));
AND2X2 AND2X2_1119 ( .A(_abc_44694_new_n2713_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n2714_));
AND2X2 AND2X2_112 ( .A(_abc_44694_new_n813_), .B(_abc_44694_new_n812_), .Y(_abc_44694_new_n814_));
AND2X2 AND2X2_1120 ( .A(_abc_44694_new_n2712_), .B(_abc_44694_new_n2714_), .Y(_0pc_q_31_0__31_));
AND2X2 AND2X2_1121 ( .A(_abc_44694_new_n1073_), .B(_abc_44694_new_n1156_), .Y(_abc_44694_new_n2717_));
AND2X2 AND2X2_1122 ( .A(_abc_44694_new_n1100_), .B(_abc_44694_new_n1076_), .Y(_abc_44694_new_n2718_));
AND2X2 AND2X2_1123 ( .A(alu_op_r_6_), .B(alu_op_r_7_), .Y(_abc_44694_new_n2720_));
AND2X2 AND2X2_1124 ( .A(_abc_44694_new_n1058_), .B(_abc_44694_new_n2720_), .Y(_abc_44694_new_n2721_));
AND2X2 AND2X2_1125 ( .A(_abc_44694_new_n1052_), .B(_abc_44694_new_n2721_), .Y(_abc_44694_new_n2722_));
AND2X2 AND2X2_1126 ( .A(_abc_44694_new_n2722_), .B(_abc_44694_new_n2719_), .Y(_abc_44694_new_n2723_));
AND2X2 AND2X2_1127 ( .A(_abc_44694_new_n2729_), .B(_abc_44694_new_n1114__bF_buf3), .Y(_abc_44694_new_n2730_));
AND2X2 AND2X2_1128 ( .A(_abc_44694_new_n2732_), .B(opcode_q_21_), .Y(_abc_44694_new_n2733_));
AND2X2 AND2X2_1129 ( .A(_abc_44694_new_n1179__bF_buf2), .B(opcode_q_22_), .Y(_abc_44694_new_n2735_));
AND2X2 AND2X2_113 ( .A(_abc_44694_new_n814_), .B(_abc_44694_new_n673__bF_buf1), .Y(_abc_44694_new_n815_));
AND2X2 AND2X2_1130 ( .A(_abc_44694_new_n2732_), .B(_abc_44694_new_n2735_), .Y(_0ex_rd_q_4_0__1_));
AND2X2 AND2X2_1131 ( .A(_abc_44694_new_n1179__bF_buf1), .B(opcode_q_23_), .Y(_abc_44694_new_n2737_));
AND2X2 AND2X2_1132 ( .A(_abc_44694_new_n2732_), .B(_abc_44694_new_n2737_), .Y(_0ex_rd_q_4_0__2_));
AND2X2 AND2X2_1133 ( .A(_abc_44694_new_n2732_), .B(opcode_q_24_), .Y(_abc_44694_new_n2739_));
AND2X2 AND2X2_1134 ( .A(_abc_44694_new_n1179__bF_buf0), .B(opcode_q_25_), .Y(_abc_44694_new_n2741_));
AND2X2 AND2X2_1135 ( .A(_abc_44694_new_n2732_), .B(_abc_44694_new_n2741_), .Y(_0ex_rd_q_4_0__4_));
AND2X2 AND2X2_1136 ( .A(_abc_44694_new_n1184_), .B(_abc_44694_new_n1085_), .Y(_abc_44694_new_n2743_));
AND2X2 AND2X2_1137 ( .A(_abc_44694_new_n1147_), .B(_abc_44694_new_n1057_), .Y(_abc_44694_new_n2745_));
AND2X2 AND2X2_1138 ( .A(_abc_44694_new_n1056_), .B(alu_op_r_5_), .Y(_abc_44694_new_n2747_));
AND2X2 AND2X2_1139 ( .A(_abc_44694_new_n1142_), .B(_abc_44694_new_n2747_), .Y(_abc_44694_new_n2748_));
AND2X2 AND2X2_114 ( .A(_abc_44694_new_n801_), .B(_abc_44694_new_n643_), .Y(_abc_44694_new_n816_));
AND2X2 AND2X2_1140 ( .A(_abc_44694_new_n2752_), .B(alu_op_r_0_), .Y(_abc_44694_new_n2753_));
AND2X2 AND2X2_1141 ( .A(_abc_44694_new_n2755_), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n2756_));
AND2X2 AND2X2_1142 ( .A(_abc_44694_new_n2752_), .B(alu_op_r_1_), .Y(_abc_44694_new_n2758_));
AND2X2 AND2X2_1143 ( .A(_abc_44694_new_n2755_), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n2759_));
AND2X2 AND2X2_1144 ( .A(_abc_44694_new_n2752_), .B(alu_op_r_2_), .Y(_abc_44694_new_n2761_));
AND2X2 AND2X2_1145 ( .A(_abc_44694_new_n2755_), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n2762_));
AND2X2 AND2X2_1146 ( .A(_abc_44694_new_n2752_), .B(alu_op_r_3_), .Y(_abc_44694_new_n2764_));
AND2X2 AND2X2_1147 ( .A(_abc_44694_new_n2755_), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n2765_));
AND2X2 AND2X2_1148 ( .A(_abc_44694_new_n2752_), .B(int32_r_4_), .Y(_abc_44694_new_n2767_));
AND2X2 AND2X2_1149 ( .A(_abc_44694_new_n2755_), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n2768_));
AND2X2 AND2X2_115 ( .A(_abc_44694_new_n818_), .B(_abc_44694_new_n811_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_));
AND2X2 AND2X2_1150 ( .A(_abc_44694_new_n2752_), .B(int32_r_5_), .Y(_abc_44694_new_n2770_));
AND2X2 AND2X2_1151 ( .A(_abc_44694_new_n2755_), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n2771_));
AND2X2 AND2X2_1152 ( .A(_abc_44694_new_n2743_), .B(_abc_44694_new_n1188_), .Y(_abc_44694_new_n2773_));
AND2X2 AND2X2_1153 ( .A(_abc_44694_new_n2775_), .B(alu_op_r_4_), .Y(_abc_44694_new_n2776_));
AND2X2 AND2X2_1154 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n2777_));
AND2X2 AND2X2_1155 ( .A(_abc_44694_new_n2779__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n2780_));
AND2X2 AND2X2_1156 ( .A(_abc_44694_new_n2775_), .B(alu_op_r_5_), .Y(_abc_44694_new_n2782_));
AND2X2 AND2X2_1157 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n2783_));
AND2X2 AND2X2_1158 ( .A(_abc_44694_new_n2779__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n2785_));
AND2X2 AND2X2_1159 ( .A(_abc_44694_new_n2775_), .B(alu_op_r_6_), .Y(_abc_44694_new_n2787_));
AND2X2 AND2X2_116 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[9] ), .Y(_abc_44694_new_n820_));
AND2X2 AND2X2_1160 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n2788_));
AND2X2 AND2X2_1161 ( .A(_abc_44694_new_n2779__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n2790_));
AND2X2 AND2X2_1162 ( .A(_abc_44694_new_n2775_), .B(alu_op_r_7_), .Y(_abc_44694_new_n2792_));
AND2X2 AND2X2_1163 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n2793_));
AND2X2 AND2X2_1164 ( .A(_abc_44694_new_n2779__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n2795_));
AND2X2 AND2X2_1165 ( .A(_abc_44694_new_n2775_), .B(int32_r_10_), .Y(_abc_44694_new_n2797_));
AND2X2 AND2X2_1166 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n2798_));
AND2X2 AND2X2_1167 ( .A(_abc_44694_new_n2779__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n2800_));
AND2X2 AND2X2_1168 ( .A(_abc_44694_new_n2775_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_44694_new_n2802_));
AND2X2 AND2X2_1169 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n2803_));
AND2X2 AND2X2_117 ( .A(_abc_44694_new_n676_), .B(_abc_44694_new_n707_), .Y(_abc_44694_new_n821_));
AND2X2 AND2X2_1170 ( .A(_abc_44694_new_n2779__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n2805_));
AND2X2 AND2X2_1171 ( .A(_abc_44694_new_n2775_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_44694_new_n2807_));
AND2X2 AND2X2_1172 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n2808_));
AND2X2 AND2X2_1173 ( .A(_abc_44694_new_n2779__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n2810_));
AND2X2 AND2X2_1174 ( .A(_abc_44694_new_n2775_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_44694_new_n2812_));
AND2X2 AND2X2_1175 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n2813_));
AND2X2 AND2X2_1176 ( .A(_abc_44694_new_n2779__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n2815_));
AND2X2 AND2X2_1177 ( .A(_abc_44694_new_n2775_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_44694_new_n2817_));
AND2X2 AND2X2_1178 ( .A(_abc_44694_new_n1086_), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n2818_));
AND2X2 AND2X2_1179 ( .A(_abc_44694_new_n2779__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n2820_));
AND2X2 AND2X2_118 ( .A(_abc_44694_new_n822_), .B(_abc_44694_new_n673__bF_buf0), .Y(_abc_44694_new_n823_));
AND2X2 AND2X2_1180 ( .A(_abc_44694_new_n2779__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n2823_));
AND2X2 AND2X2_1181 ( .A(_abc_44694_new_n1146_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2_), .Y(_abc_44694_new_n2825_));
AND2X2 AND2X2_1182 ( .A(_abc_44694_new_n2827_), .B(_abc_44694_new_n2824_), .Y(_abc_44694_new_n2828_));
AND2X2 AND2X2_1183 ( .A(_abc_44694_new_n2829_), .B(_abc_44694_new_n2822_), .Y(alu_input_b_r_15_));
AND2X2 AND2X2_1184 ( .A(_abc_44694_new_n1084__bF_buf2), .B(_abc_44694_new_n2833_), .Y(_abc_44694_new_n2834_));
AND2X2 AND2X2_1185 ( .A(_abc_44694_new_n2826__bF_buf2), .B(_abc_44694_new_n2836_), .Y(_abc_44694_new_n2837_));
AND2X2 AND2X2_1186 ( .A(_abc_44694_new_n2838_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2839_));
AND2X2 AND2X2_1187 ( .A(_abc_44694_new_n2840_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2841_));
AND2X2 AND2X2_1188 ( .A(_abc_44694_new_n2779__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_44694_new_n2842_));
AND2X2 AND2X2_1189 ( .A(_abc_44694_new_n2826__bF_buf1), .B(_abc_44694_new_n2844_), .Y(_abc_44694_new_n2845_));
AND2X2 AND2X2_119 ( .A(_abc_44694_new_n824_), .B(_abc_44694_new_n825_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_));
AND2X2 AND2X2_1190 ( .A(_abc_44694_new_n2846_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2847_));
AND2X2 AND2X2_1191 ( .A(_abc_44694_new_n2848_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2849_));
AND2X2 AND2X2_1192 ( .A(_abc_44694_new_n2779__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_44694_new_n2850_));
AND2X2 AND2X2_1193 ( .A(_abc_44694_new_n2826__bF_buf0), .B(_abc_44694_new_n2852_), .Y(_abc_44694_new_n2853_));
AND2X2 AND2X2_1194 ( .A(_abc_44694_new_n2854_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2855_));
AND2X2 AND2X2_1195 ( .A(_abc_44694_new_n2856_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2857_));
AND2X2 AND2X2_1196 ( .A(_abc_44694_new_n2779__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_44694_new_n2858_));
AND2X2 AND2X2_1197 ( .A(_abc_44694_new_n2826__bF_buf3), .B(_abc_44694_new_n2860_), .Y(_abc_44694_new_n2861_));
AND2X2 AND2X2_1198 ( .A(_abc_44694_new_n2862_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2863_));
AND2X2 AND2X2_1199 ( .A(_abc_44694_new_n2864_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2865_));
AND2X2 AND2X2_12 ( .A(_abc_44694_new_n617_), .B(inst_r_5_), .Y(_abc_44694_new_n637_));
AND2X2 AND2X2_120 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[10] ), .Y(_abc_44694_new_n827_));
AND2X2 AND2X2_1200 ( .A(_abc_44694_new_n2779__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_44694_new_n2866_));
AND2X2 AND2X2_1201 ( .A(_abc_44694_new_n2826__bF_buf2), .B(_abc_44694_new_n2868_), .Y(_abc_44694_new_n2869_));
AND2X2 AND2X2_1202 ( .A(_abc_44694_new_n2870_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2871_));
AND2X2 AND2X2_1203 ( .A(_abc_44694_new_n2872_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2873_));
AND2X2 AND2X2_1204 ( .A(_abc_44694_new_n2779__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_44694_new_n2874_));
AND2X2 AND2X2_1205 ( .A(_abc_44694_new_n2826__bF_buf1), .B(_abc_44694_new_n2876_), .Y(_abc_44694_new_n2877_));
AND2X2 AND2X2_1206 ( .A(_abc_44694_new_n2878_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2879_));
AND2X2 AND2X2_1207 ( .A(_abc_44694_new_n2880_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2881_));
AND2X2 AND2X2_1208 ( .A(_abc_44694_new_n2779__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_44694_new_n2882_));
AND2X2 AND2X2_1209 ( .A(_abc_44694_new_n2826__bF_buf0), .B(_abc_44694_new_n2884_), .Y(_abc_44694_new_n2885_));
AND2X2 AND2X2_121 ( .A(_abc_44694_new_n676_), .B(_abc_44694_new_n723_), .Y(_abc_44694_new_n828_));
AND2X2 AND2X2_1210 ( .A(_abc_44694_new_n2886_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2887_));
AND2X2 AND2X2_1211 ( .A(_abc_44694_new_n2888_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2889_));
AND2X2 AND2X2_1212 ( .A(_abc_44694_new_n2779__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_44694_new_n2890_));
AND2X2 AND2X2_1213 ( .A(_abc_44694_new_n2826__bF_buf3), .B(_abc_44694_new_n2892_), .Y(_abc_44694_new_n2893_));
AND2X2 AND2X2_1214 ( .A(_abc_44694_new_n2894_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2895_));
AND2X2 AND2X2_1215 ( .A(_abc_44694_new_n2896_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2897_));
AND2X2 AND2X2_1216 ( .A(_abc_44694_new_n2779__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_44694_new_n2898_));
AND2X2 AND2X2_1217 ( .A(_abc_44694_new_n2826__bF_buf2), .B(_abc_44694_new_n2900_), .Y(_abc_44694_new_n2901_));
AND2X2 AND2X2_1218 ( .A(_abc_44694_new_n2902_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2903_));
AND2X2 AND2X2_1219 ( .A(_abc_44694_new_n2904_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2905_));
AND2X2 AND2X2_122 ( .A(_abc_44694_new_n829_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n830_));
AND2X2 AND2X2_1220 ( .A(_abc_44694_new_n2779__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_44694_new_n2906_));
AND2X2 AND2X2_1221 ( .A(_abc_44694_new_n2826__bF_buf1), .B(_abc_44694_new_n2908_), .Y(_abc_44694_new_n2909_));
AND2X2 AND2X2_1222 ( .A(_abc_44694_new_n2910_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2911_));
AND2X2 AND2X2_1223 ( .A(_abc_44694_new_n2912_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2913_));
AND2X2 AND2X2_1224 ( .A(_abc_44694_new_n2779__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_44694_new_n2914_));
AND2X2 AND2X2_1225 ( .A(_abc_44694_new_n2826__bF_buf0), .B(_abc_44694_new_n2916_), .Y(_abc_44694_new_n2917_));
AND2X2 AND2X2_1226 ( .A(_abc_44694_new_n2918_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2919_));
AND2X2 AND2X2_1227 ( .A(_abc_44694_new_n2920_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2921_));
AND2X2 AND2X2_1228 ( .A(_abc_44694_new_n2779__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_44694_new_n2922_));
AND2X2 AND2X2_1229 ( .A(_abc_44694_new_n2826__bF_buf3), .B(_abc_44694_new_n2924_), .Y(_abc_44694_new_n2925_));
AND2X2 AND2X2_123 ( .A(_abc_44694_new_n831_), .B(_abc_44694_new_n832_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_));
AND2X2 AND2X2_1230 ( .A(_abc_44694_new_n2926_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2927_));
AND2X2 AND2X2_1231 ( .A(_abc_44694_new_n2928_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2929_));
AND2X2 AND2X2_1232 ( .A(_abc_44694_new_n2779__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_44694_new_n2930_));
AND2X2 AND2X2_1233 ( .A(_abc_44694_new_n2826__bF_buf2), .B(_abc_44694_new_n2932_), .Y(_abc_44694_new_n2933_));
AND2X2 AND2X2_1234 ( .A(_abc_44694_new_n2934_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2935_));
AND2X2 AND2X2_1235 ( .A(_abc_44694_new_n2936_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2937_));
AND2X2 AND2X2_1236 ( .A(_abc_44694_new_n2779__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_44694_new_n2938_));
AND2X2 AND2X2_1237 ( .A(_abc_44694_new_n2826__bF_buf1), .B(_abc_44694_new_n2940_), .Y(_abc_44694_new_n2941_));
AND2X2 AND2X2_1238 ( .A(_abc_44694_new_n2942_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2943_));
AND2X2 AND2X2_1239 ( .A(_abc_44694_new_n2944_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2945_));
AND2X2 AND2X2_124 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[11] ), .Y(_abc_44694_new_n834_));
AND2X2 AND2X2_1240 ( .A(_abc_44694_new_n2779__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_44694_new_n2946_));
AND2X2 AND2X2_1241 ( .A(_abc_44694_new_n2826__bF_buf0), .B(_abc_44694_new_n2948_), .Y(_abc_44694_new_n2949_));
AND2X2 AND2X2_1242 ( .A(_abc_44694_new_n2950_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2951_));
AND2X2 AND2X2_1243 ( .A(_abc_44694_new_n2952_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2953_));
AND2X2 AND2X2_1244 ( .A(_abc_44694_new_n2779__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_44694_new_n2954_));
AND2X2 AND2X2_1245 ( .A(_abc_44694_new_n2826__bF_buf3), .B(_abc_44694_new_n2956_), .Y(_abc_44694_new_n2957_));
AND2X2 AND2X2_1246 ( .A(_abc_44694_new_n2958_), .B(_abc_44694_new_n2835_), .Y(_abc_44694_new_n2959_));
AND2X2 AND2X2_1247 ( .A(_abc_44694_new_n2960_), .B(_abc_44694_new_n2832_), .Y(_abc_44694_new_n2961_));
AND2X2 AND2X2_1248 ( .A(_abc_44694_new_n2779__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_44694_new_n2962_));
AND2X2 AND2X2_1249 ( .A(_abc_44694_new_n2965__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_0_), .Y(_abc_44694_new_n2966_));
AND2X2 AND2X2_125 ( .A(_abc_44694_new_n676_), .B(_abc_44694_new_n739_), .Y(_abc_44694_new_n835_));
AND2X2 AND2X2_1250 ( .A(_abc_44694_new_n1114__bF_buf2), .B(epc_q_0_), .Y(_abc_44694_new_n2967_));
AND2X2 AND2X2_1251 ( .A(_abc_44694_new_n1347__bF_buf2), .B(_abc_44694_new_n2967_), .Y(_abc_44694_new_n2968_));
AND2X2 AND2X2_1252 ( .A(_abc_44694_new_n1178__bF_buf1), .B(next_pc_r_0_), .Y(_abc_44694_new_n2970_));
AND2X2 AND2X2_1253 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_0_), .Y(_abc_44694_new_n2973_));
AND2X2 AND2X2_1254 ( .A(_abc_44694_new_n2965__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_1_), .Y(_abc_44694_new_n2975_));
AND2X2 AND2X2_1255 ( .A(_abc_44694_new_n1114__bF_buf1), .B(epc_q_1_), .Y(_abc_44694_new_n2976_));
AND2X2 AND2X2_1256 ( .A(_abc_44694_new_n1347__bF_buf1), .B(_abc_44694_new_n2976_), .Y(_abc_44694_new_n2977_));
AND2X2 AND2X2_1257 ( .A(_abc_44694_new_n1178__bF_buf0), .B(next_pc_r_1_), .Y(_abc_44694_new_n2979_));
AND2X2 AND2X2_1258 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_1_), .Y(_abc_44694_new_n2981_));
AND2X2 AND2X2_1259 ( .A(_abc_44694_new_n1027_), .B(_abc_44694_new_n1011_), .Y(_abc_44694_new_n2983_));
AND2X2 AND2X2_126 ( .A(_abc_44694_new_n836_), .B(_abc_44694_new_n673__bF_buf3), .Y(_abc_44694_new_n837_));
AND2X2 AND2X2_1260 ( .A(_abc_44694_new_n1347__bF_buf0), .B(epc_q_2_), .Y(_abc_44694_new_n2984_));
AND2X2 AND2X2_1261 ( .A(_abc_44694_new_n1037_), .B(esr_q_2_), .Y(_abc_44694_new_n2985_));
AND2X2 AND2X2_1262 ( .A(_abc_44694_new_n2987_), .B(_abc_44694_new_n1114__bF_buf0), .Y(_abc_44694_new_n2988_));
AND2X2 AND2X2_1263 ( .A(_abc_44694_new_n2965__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_44694_new_n2989_));
AND2X2 AND2X2_1264 ( .A(_abc_44694_new_n2991_), .B(_abc_44694_new_n2992_), .Y(_abc_44694_new_n2993_));
AND2X2 AND2X2_1265 ( .A(_abc_44694_new_n2972__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_2_), .Y(_abc_44694_new_n2994_));
AND2X2 AND2X2_1266 ( .A(_abc_44694_new_n2965__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_44694_new_n2996_));
AND2X2 AND2X2_1267 ( .A(_abc_44694_new_n1114__bF_buf4), .B(epc_q_3_), .Y(_abc_44694_new_n2997_));
AND2X2 AND2X2_1268 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n2997_), .Y(_abc_44694_new_n2998_));
AND2X2 AND2X2_1269 ( .A(_abc_44694_new_n1178__bF_buf3), .B(_abc_44694_new_n1448_), .Y(_abc_44694_new_n3000_));
AND2X2 AND2X2_127 ( .A(_abc_44694_new_n838_), .B(_abc_44694_new_n839_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_));
AND2X2 AND2X2_1270 ( .A(_abc_44694_new_n2972__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_3_), .Y(_abc_44694_new_n3002_));
AND2X2 AND2X2_1271 ( .A(_abc_44694_new_n1115_), .B(REGFILE_SIM_reg_bank_reg_ra_o_4_), .Y(_abc_44694_new_n3004_));
AND2X2 AND2X2_1272 ( .A(_abc_44694_new_n2965__bF_buf0), .B(_abc_44694_new_n3004_), .Y(_abc_44694_new_n3005_));
AND2X2 AND2X2_1273 ( .A(_abc_44694_new_n1114__bF_buf3), .B(epc_q_4_), .Y(_abc_44694_new_n3006_));
AND2X2 AND2X2_1274 ( .A(_abc_44694_new_n1347__bF_buf3), .B(_abc_44694_new_n3006_), .Y(_abc_44694_new_n3007_));
AND2X2 AND2X2_1275 ( .A(_abc_44694_new_n1178__bF_buf2), .B(_abc_44694_new_n1486_), .Y(_abc_44694_new_n3009_));
AND2X2 AND2X2_1276 ( .A(_abc_44694_new_n2972__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_4_), .Y(_abc_44694_new_n3011_));
AND2X2 AND2X2_1277 ( .A(_abc_44694_new_n2965__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_5_), .Y(_abc_44694_new_n3013_));
AND2X2 AND2X2_1278 ( .A(_abc_44694_new_n1114__bF_buf2), .B(epc_q_5_), .Y(_abc_44694_new_n3014_));
AND2X2 AND2X2_1279 ( .A(_abc_44694_new_n1347__bF_buf2), .B(_abc_44694_new_n3014_), .Y(_abc_44694_new_n3015_));
AND2X2 AND2X2_128 ( .A(_abc_44694_new_n843_), .B(_abc_44694_new_n842_), .Y(_abc_44694_new_n844_));
AND2X2 AND2X2_1280 ( .A(_abc_44694_new_n1178__bF_buf1), .B(_abc_44694_new_n1501_), .Y(_abc_44694_new_n3017_));
AND2X2 AND2X2_1281 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_5_), .Y(_abc_44694_new_n3019_));
AND2X2 AND2X2_1282 ( .A(_abc_44694_new_n1115_), .B(REGFILE_SIM_reg_bank_reg_ra_o_6_), .Y(_abc_44694_new_n3021_));
AND2X2 AND2X2_1283 ( .A(_abc_44694_new_n2965__bF_buf3), .B(_abc_44694_new_n3021_), .Y(_abc_44694_new_n3022_));
AND2X2 AND2X2_1284 ( .A(_abc_44694_new_n1114__bF_buf1), .B(epc_q_6_), .Y(_abc_44694_new_n3023_));
AND2X2 AND2X2_1285 ( .A(_abc_44694_new_n1347__bF_buf1), .B(_abc_44694_new_n3023_), .Y(_abc_44694_new_n3024_));
AND2X2 AND2X2_1286 ( .A(_abc_44694_new_n1539_), .B(_abc_44694_new_n1178__bF_buf0), .Y(_abc_44694_new_n3026_));
AND2X2 AND2X2_1287 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_6_), .Y(_abc_44694_new_n3028_));
AND2X2 AND2X2_1288 ( .A(_abc_44694_new_n2965__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_7_), .Y(_abc_44694_new_n3030_));
AND2X2 AND2X2_1289 ( .A(_abc_44694_new_n1114__bF_buf0), .B(epc_q_7_), .Y(_abc_44694_new_n3031_));
AND2X2 AND2X2_129 ( .A(_abc_44694_new_n844_), .B(_abc_44694_new_n673__bF_buf2), .Y(_abc_44694_new_n845_));
AND2X2 AND2X2_1290 ( .A(_abc_44694_new_n1347__bF_buf0), .B(_abc_44694_new_n3031_), .Y(_abc_44694_new_n3032_));
AND2X2 AND2X2_1291 ( .A(_abc_44694_new_n1578_), .B(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n3034_));
AND2X2 AND2X2_1292 ( .A(_abc_44694_new_n2972__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_7_), .Y(_abc_44694_new_n3036_));
AND2X2 AND2X2_1293 ( .A(_abc_44694_new_n1115_), .B(REGFILE_SIM_reg_bank_reg_ra_o_8_), .Y(_abc_44694_new_n3038_));
AND2X2 AND2X2_1294 ( .A(_abc_44694_new_n2965__bF_buf1), .B(_abc_44694_new_n3038_), .Y(_abc_44694_new_n3039_));
AND2X2 AND2X2_1295 ( .A(_abc_44694_new_n1114__bF_buf4), .B(epc_q_8_), .Y(_abc_44694_new_n3040_));
AND2X2 AND2X2_1296 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n3040_), .Y(_abc_44694_new_n3041_));
AND2X2 AND2X2_1297 ( .A(_abc_44694_new_n1617_), .B(_abc_44694_new_n1178__bF_buf3), .Y(_abc_44694_new_n3043_));
AND2X2 AND2X2_1298 ( .A(_abc_44694_new_n2972__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_8_), .Y(_abc_44694_new_n3045_));
AND2X2 AND2X2_1299 ( .A(_abc_44694_new_n1347__bF_buf3), .B(epc_q_9_), .Y(_abc_44694_new_n3047_));
AND2X2 AND2X2_13 ( .A(inst_r_1_), .B(inst_r_0_), .Y(_abc_44694_new_n638_));
AND2X2 AND2X2_130 ( .A(_abc_44694_new_n846_), .B(_abc_44694_new_n841_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_));
AND2X2 AND2X2_1300 ( .A(_abc_44694_new_n1037_), .B(esr_q_9_), .Y(_abc_44694_new_n3048_));
AND2X2 AND2X2_1301 ( .A(_abc_44694_new_n1276_), .B(_abc_44694_new_n1011_), .Y(_abc_44694_new_n3051_));
AND2X2 AND2X2_1302 ( .A(_abc_44694_new_n2965__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_9_), .Y(_abc_44694_new_n3053_));
AND2X2 AND2X2_1303 ( .A(_abc_44694_new_n3052_), .B(_abc_44694_new_n3054_), .Y(_abc_44694_new_n3055_));
AND2X2 AND2X2_1304 ( .A(_abc_44694_new_n1654_), .B(_abc_44694_new_n1178__bF_buf2), .Y(_abc_44694_new_n3056_));
AND2X2 AND2X2_1305 ( .A(_abc_44694_new_n2972__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_9_), .Y(_abc_44694_new_n3058_));
AND2X2 AND2X2_1306 ( .A(_abc_44694_new_n2965__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_10_), .Y(_abc_44694_new_n3060_));
AND2X2 AND2X2_1307 ( .A(_abc_44694_new_n1347__bF_buf2), .B(epc_q_10_), .Y(_abc_44694_new_n3061_));
AND2X2 AND2X2_1308 ( .A(_abc_44694_new_n1037_), .B(esr_q_10_), .Y(_abc_44694_new_n3062_));
AND2X2 AND2X2_1309 ( .A(_abc_44694_new_n1309_), .B(_abc_44694_new_n1011_), .Y(_abc_44694_new_n3064_));
AND2X2 AND2X2_131 ( .A(_abc_44694_new_n850_), .B(_abc_44694_new_n849_), .Y(_abc_44694_new_n851_));
AND2X2 AND2X2_1310 ( .A(_abc_44694_new_n3065_), .B(_abc_44694_new_n1114__bF_buf2), .Y(_abc_44694_new_n3066_));
AND2X2 AND2X2_1311 ( .A(_abc_44694_new_n1696_), .B(_abc_44694_new_n1178__bF_buf1), .Y(_abc_44694_new_n3068_));
AND2X2 AND2X2_1312 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_10_), .Y(_abc_44694_new_n3070_));
AND2X2 AND2X2_1313 ( .A(_abc_44694_new_n1347__bF_buf1), .B(epc_q_11_), .Y(_abc_44694_new_n3072_));
AND2X2 AND2X2_1314 ( .A(_abc_44694_new_n2965__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_44694_new_n3074_));
AND2X2 AND2X2_1315 ( .A(_abc_44694_new_n3075_), .B(_abc_44694_new_n3073_), .Y(_abc_44694_new_n3076_));
AND2X2 AND2X2_1316 ( .A(_abc_44694_new_n3077_), .B(_abc_44694_new_n3078_), .Y(_abc_44694_new_n3079_));
AND2X2 AND2X2_1317 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_44694_new_n3080_));
AND2X2 AND2X2_1318 ( .A(_abc_44694_new_n2965__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_44694_new_n3082_));
AND2X2 AND2X2_1319 ( .A(_abc_44694_new_n1114__bF_buf0), .B(epc_q_12_), .Y(_abc_44694_new_n3083_));
AND2X2 AND2X2_132 ( .A(_abc_44694_new_n851_), .B(_abc_44694_new_n673__bF_buf1), .Y(_abc_44694_new_n852_));
AND2X2 AND2X2_1320 ( .A(_abc_44694_new_n1347__bF_buf0), .B(_abc_44694_new_n3083_), .Y(_abc_44694_new_n3084_));
AND2X2 AND2X2_1321 ( .A(_abc_44694_new_n1770_), .B(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n3086_));
AND2X2 AND2X2_1322 ( .A(_abc_44694_new_n2972__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_44694_new_n3088_));
AND2X2 AND2X2_1323 ( .A(_abc_44694_new_n2965__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_44694_new_n3090_));
AND2X2 AND2X2_1324 ( .A(_abc_44694_new_n1114__bF_buf4), .B(epc_q_13_), .Y(_abc_44694_new_n3091_));
AND2X2 AND2X2_1325 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n3091_), .Y(_abc_44694_new_n3092_));
AND2X2 AND2X2_1326 ( .A(_abc_44694_new_n1812_), .B(_abc_44694_new_n1178__bF_buf3), .Y(_abc_44694_new_n3094_));
AND2X2 AND2X2_1327 ( .A(_abc_44694_new_n2972__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_44694_new_n3096_));
AND2X2 AND2X2_1328 ( .A(_abc_44694_new_n2965__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_44694_new_n3098_));
AND2X2 AND2X2_1329 ( .A(_abc_44694_new_n1114__bF_buf3), .B(epc_q_14_), .Y(_abc_44694_new_n3099_));
AND2X2 AND2X2_133 ( .A(_abc_44694_new_n853_), .B(_abc_44694_new_n848_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_));
AND2X2 AND2X2_1330 ( .A(_abc_44694_new_n1347__bF_buf3), .B(_abc_44694_new_n3099_), .Y(_abc_44694_new_n3100_));
AND2X2 AND2X2_1331 ( .A(_abc_44694_new_n1851_), .B(_abc_44694_new_n1178__bF_buf2), .Y(_abc_44694_new_n3102_));
AND2X2 AND2X2_1332 ( .A(_abc_44694_new_n2972__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_44694_new_n3104_));
AND2X2 AND2X2_1333 ( .A(_abc_44694_new_n2965__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_44694_new_n3106_));
AND2X2 AND2X2_1334 ( .A(_abc_44694_new_n1114__bF_buf2), .B(epc_q_15_), .Y(_abc_44694_new_n3107_));
AND2X2 AND2X2_1335 ( .A(_abc_44694_new_n1347__bF_buf2), .B(_abc_44694_new_n3107_), .Y(_abc_44694_new_n3108_));
AND2X2 AND2X2_1336 ( .A(_abc_44694_new_n1888_), .B(_abc_44694_new_n1178__bF_buf1), .Y(_abc_44694_new_n3110_));
AND2X2 AND2X2_1337 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_44694_new_n3112_));
AND2X2 AND2X2_1338 ( .A(_abc_44694_new_n1186__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_44694_new_n3115_));
AND2X2 AND2X2_1339 ( .A(_abc_44694_new_n2965__bF_buf3), .B(_abc_44694_new_n3115_), .Y(_abc_44694_new_n3116_));
AND2X2 AND2X2_134 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[14] ), .Y(_abc_44694_new_n855_));
AND2X2 AND2X2_1340 ( .A(_abc_44694_new_n1185__bF_buf2), .B(alu_op_r_0_), .Y(_abc_44694_new_n3117_));
AND2X2 AND2X2_1341 ( .A(_abc_44694_new_n1114__bF_buf1), .B(epc_q_16_), .Y(_abc_44694_new_n3119_));
AND2X2 AND2X2_1342 ( .A(_abc_44694_new_n1347__bF_buf1), .B(_abc_44694_new_n3119_), .Y(_abc_44694_new_n3120_));
AND2X2 AND2X2_1343 ( .A(_abc_44694_new_n3114_), .B(_abc_44694_new_n3122_), .Y(_abc_44694_new_n3123_));
AND2X2 AND2X2_1344 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_44694_new_n3124_));
AND2X2 AND2X2_1345 ( .A(_abc_44694_new_n1186__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_44694_new_n3127_));
AND2X2 AND2X2_1346 ( .A(_abc_44694_new_n2965__bF_buf2), .B(_abc_44694_new_n3127_), .Y(_abc_44694_new_n3128_));
AND2X2 AND2X2_1347 ( .A(_abc_44694_new_n1185__bF_buf1), .B(alu_op_r_1_), .Y(_abc_44694_new_n3129_));
AND2X2 AND2X2_1348 ( .A(_abc_44694_new_n1114__bF_buf0), .B(epc_q_17_), .Y(_abc_44694_new_n3131_));
AND2X2 AND2X2_1349 ( .A(_abc_44694_new_n1347__bF_buf0), .B(_abc_44694_new_n3131_), .Y(_abc_44694_new_n3132_));
AND2X2 AND2X2_135 ( .A(_abc_44694_new_n676_), .B(_abc_44694_new_n787_), .Y(_abc_44694_new_n856_));
AND2X2 AND2X2_1350 ( .A(_abc_44694_new_n3126_), .B(_abc_44694_new_n3134_), .Y(_abc_44694_new_n3135_));
AND2X2 AND2X2_1351 ( .A(_abc_44694_new_n2972__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_44694_new_n3136_));
AND2X2 AND2X2_1352 ( .A(_abc_44694_new_n1186__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_44694_new_n3139_));
AND2X2 AND2X2_1353 ( .A(_abc_44694_new_n2965__bF_buf1), .B(_abc_44694_new_n3139_), .Y(_abc_44694_new_n3140_));
AND2X2 AND2X2_1354 ( .A(_abc_44694_new_n1185__bF_buf0), .B(alu_op_r_2_), .Y(_abc_44694_new_n3141_));
AND2X2 AND2X2_1355 ( .A(_abc_44694_new_n1114__bF_buf4), .B(epc_q_18_), .Y(_abc_44694_new_n3143_));
AND2X2 AND2X2_1356 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n3143_), .Y(_abc_44694_new_n3144_));
AND2X2 AND2X2_1357 ( .A(_abc_44694_new_n3138_), .B(_abc_44694_new_n3146_), .Y(_abc_44694_new_n3147_));
AND2X2 AND2X2_1358 ( .A(_abc_44694_new_n2972__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_44694_new_n3148_));
AND2X2 AND2X2_1359 ( .A(_abc_44694_new_n1186__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_44694_new_n3151_));
AND2X2 AND2X2_136 ( .A(_abc_44694_new_n857_), .B(_abc_44694_new_n673__bF_buf0), .Y(_abc_44694_new_n858_));
AND2X2 AND2X2_1360 ( .A(_abc_44694_new_n2965__bF_buf0), .B(_abc_44694_new_n3151_), .Y(_abc_44694_new_n3152_));
AND2X2 AND2X2_1361 ( .A(_abc_44694_new_n1185__bF_buf3), .B(alu_op_r_3_), .Y(_abc_44694_new_n3153_));
AND2X2 AND2X2_1362 ( .A(_abc_44694_new_n1114__bF_buf3), .B(epc_q_19_), .Y(_abc_44694_new_n3155_));
AND2X2 AND2X2_1363 ( .A(_abc_44694_new_n1347__bF_buf3), .B(_abc_44694_new_n3155_), .Y(_abc_44694_new_n3156_));
AND2X2 AND2X2_1364 ( .A(_abc_44694_new_n3150_), .B(_abc_44694_new_n3158_), .Y(_abc_44694_new_n3159_));
AND2X2 AND2X2_1365 ( .A(_abc_44694_new_n2972__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_44694_new_n3160_));
AND2X2 AND2X2_1366 ( .A(_abc_44694_new_n1186__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_44694_new_n3163_));
AND2X2 AND2X2_1367 ( .A(_abc_44694_new_n2965__bF_buf4), .B(_abc_44694_new_n3163_), .Y(_abc_44694_new_n3164_));
AND2X2 AND2X2_1368 ( .A(_abc_44694_new_n1185__bF_buf2), .B(int32_r_4_), .Y(_abc_44694_new_n3165_));
AND2X2 AND2X2_1369 ( .A(_abc_44694_new_n1114__bF_buf2), .B(epc_q_20_), .Y(_abc_44694_new_n3167_));
AND2X2 AND2X2_137 ( .A(_abc_44694_new_n859_), .B(_abc_44694_new_n860_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_));
AND2X2 AND2X2_1370 ( .A(_abc_44694_new_n1347__bF_buf2), .B(_abc_44694_new_n3167_), .Y(_abc_44694_new_n3168_));
AND2X2 AND2X2_1371 ( .A(_abc_44694_new_n3162_), .B(_abc_44694_new_n3170_), .Y(_abc_44694_new_n3171_));
AND2X2 AND2X2_1372 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_44694_new_n3172_));
AND2X2 AND2X2_1373 ( .A(_abc_44694_new_n1186__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_44694_new_n3175_));
AND2X2 AND2X2_1374 ( .A(_abc_44694_new_n2965__bF_buf3), .B(_abc_44694_new_n3175_), .Y(_abc_44694_new_n3176_));
AND2X2 AND2X2_1375 ( .A(_abc_44694_new_n1185__bF_buf1), .B(int32_r_5_), .Y(_abc_44694_new_n3177_));
AND2X2 AND2X2_1376 ( .A(_abc_44694_new_n1114__bF_buf1), .B(epc_q_21_), .Y(_abc_44694_new_n3179_));
AND2X2 AND2X2_1377 ( .A(_abc_44694_new_n1347__bF_buf1), .B(_abc_44694_new_n3179_), .Y(_abc_44694_new_n3180_));
AND2X2 AND2X2_1378 ( .A(_abc_44694_new_n3174_), .B(_abc_44694_new_n3182_), .Y(_abc_44694_new_n3183_));
AND2X2 AND2X2_1379 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_44694_new_n3184_));
AND2X2 AND2X2_138 ( .A(_abc_44694_new_n864_), .B(_abc_44694_new_n863_), .Y(_abc_44694_new_n865_));
AND2X2 AND2X2_1380 ( .A(_abc_44694_new_n1186__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_44694_new_n3187_));
AND2X2 AND2X2_1381 ( .A(_abc_44694_new_n2965__bF_buf2), .B(_abc_44694_new_n3187_), .Y(_abc_44694_new_n3188_));
AND2X2 AND2X2_1382 ( .A(_abc_44694_new_n1185__bF_buf0), .B(alu_op_r_4_), .Y(_abc_44694_new_n3189_));
AND2X2 AND2X2_1383 ( .A(_abc_44694_new_n1114__bF_buf0), .B(epc_q_22_), .Y(_abc_44694_new_n3191_));
AND2X2 AND2X2_1384 ( .A(_abc_44694_new_n1347__bF_buf0), .B(_abc_44694_new_n3191_), .Y(_abc_44694_new_n3192_));
AND2X2 AND2X2_1385 ( .A(_abc_44694_new_n3186_), .B(_abc_44694_new_n3194_), .Y(_abc_44694_new_n3195_));
AND2X2 AND2X2_1386 ( .A(_abc_44694_new_n2972__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_44694_new_n3196_));
AND2X2 AND2X2_1387 ( .A(_abc_44694_new_n1186__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_44694_new_n3199_));
AND2X2 AND2X2_1388 ( .A(_abc_44694_new_n2965__bF_buf1), .B(_abc_44694_new_n3199_), .Y(_abc_44694_new_n3200_));
AND2X2 AND2X2_1389 ( .A(_abc_44694_new_n1185__bF_buf3), .B(alu_op_r_5_), .Y(_abc_44694_new_n3201_));
AND2X2 AND2X2_139 ( .A(_abc_44694_new_n865_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n866_));
AND2X2 AND2X2_1390 ( .A(_abc_44694_new_n1114__bF_buf4), .B(epc_q_23_), .Y(_abc_44694_new_n3203_));
AND2X2 AND2X2_1391 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n3203_), .Y(_abc_44694_new_n3204_));
AND2X2 AND2X2_1392 ( .A(_abc_44694_new_n3198_), .B(_abc_44694_new_n3206_), .Y(_abc_44694_new_n3207_));
AND2X2 AND2X2_1393 ( .A(_abc_44694_new_n2972__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_44694_new_n3208_));
AND2X2 AND2X2_1394 ( .A(_abc_44694_new_n1186__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_44694_new_n3211_));
AND2X2 AND2X2_1395 ( .A(_abc_44694_new_n2965__bF_buf0), .B(_abc_44694_new_n3211_), .Y(_abc_44694_new_n3212_));
AND2X2 AND2X2_1396 ( .A(_abc_44694_new_n1185__bF_buf2), .B(alu_op_r_6_), .Y(_abc_44694_new_n3213_));
AND2X2 AND2X2_1397 ( .A(_abc_44694_new_n1114__bF_buf3), .B(epc_q_24_), .Y(_abc_44694_new_n3215_));
AND2X2 AND2X2_1398 ( .A(_abc_44694_new_n1347__bF_buf3), .B(_abc_44694_new_n3215_), .Y(_abc_44694_new_n3216_));
AND2X2 AND2X2_1399 ( .A(_abc_44694_new_n3210_), .B(_abc_44694_new_n3218_), .Y(_abc_44694_new_n3219_));
AND2X2 AND2X2_14 ( .A(_abc_44694_new_n620_), .B(_abc_44694_new_n631_), .Y(_abc_44694_new_n639_));
AND2X2 AND2X2_140 ( .A(_abc_44694_new_n867_), .B(_abc_44694_new_n862_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_));
AND2X2 AND2X2_1400 ( .A(_abc_44694_new_n2972__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_44694_new_n3220_));
AND2X2 AND2X2_1401 ( .A(_abc_44694_new_n1186__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_44694_new_n3223_));
AND2X2 AND2X2_1402 ( .A(_abc_44694_new_n2965__bF_buf4), .B(_abc_44694_new_n3223_), .Y(_abc_44694_new_n3224_));
AND2X2 AND2X2_1403 ( .A(_abc_44694_new_n1185__bF_buf1), .B(alu_op_r_7_), .Y(_abc_44694_new_n3225_));
AND2X2 AND2X2_1404 ( .A(_abc_44694_new_n1114__bF_buf2), .B(epc_q_25_), .Y(_abc_44694_new_n3227_));
AND2X2 AND2X2_1405 ( .A(_abc_44694_new_n1347__bF_buf2), .B(_abc_44694_new_n3227_), .Y(_abc_44694_new_n3228_));
AND2X2 AND2X2_1406 ( .A(_abc_44694_new_n3222_), .B(_abc_44694_new_n3230_), .Y(_abc_44694_new_n3231_));
AND2X2 AND2X2_1407 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_44694_new_n3232_));
AND2X2 AND2X2_1408 ( .A(_abc_44694_new_n1186__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_44694_new_n3235_));
AND2X2 AND2X2_1409 ( .A(_abc_44694_new_n2965__bF_buf3), .B(_abc_44694_new_n3235_), .Y(_abc_44694_new_n3236_));
AND2X2 AND2X2_141 ( .A(_abc_44694_new_n632_), .B(_abc_44694_new_n645_), .Y(_abc_44694_new_n869_));
AND2X2 AND2X2_1410 ( .A(_abc_44694_new_n1185__bF_buf0), .B(int32_r_10_), .Y(_abc_44694_new_n3237_));
AND2X2 AND2X2_1411 ( .A(_abc_44694_new_n1114__bF_buf1), .B(epc_q_26_), .Y(_abc_44694_new_n3239_));
AND2X2 AND2X2_1412 ( .A(_abc_44694_new_n1347__bF_buf1), .B(_abc_44694_new_n3239_), .Y(_abc_44694_new_n3240_));
AND2X2 AND2X2_1413 ( .A(_abc_44694_new_n3234_), .B(_abc_44694_new_n3242_), .Y(_abc_44694_new_n3243_));
AND2X2 AND2X2_1414 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_44694_new_n3244_));
AND2X2 AND2X2_1415 ( .A(_abc_44694_new_n1186__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_44694_new_n3247_));
AND2X2 AND2X2_1416 ( .A(_abc_44694_new_n2965__bF_buf2), .B(_abc_44694_new_n3247_), .Y(_abc_44694_new_n3248_));
AND2X2 AND2X2_1417 ( .A(_abc_44694_new_n1185__bF_buf3), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_44694_new_n3249_));
AND2X2 AND2X2_1418 ( .A(_abc_44694_new_n1114__bF_buf0), .B(epc_q_27_), .Y(_abc_44694_new_n3251_));
AND2X2 AND2X2_1419 ( .A(_abc_44694_new_n1347__bF_buf0), .B(_abc_44694_new_n3251_), .Y(_abc_44694_new_n3252_));
AND2X2 AND2X2_142 ( .A(_abc_44694_new_n869_), .B(_abc_44694_new_n637_), .Y(_abc_44694_new_n870_));
AND2X2 AND2X2_1420 ( .A(_abc_44694_new_n3246_), .B(_abc_44694_new_n3254_), .Y(_abc_44694_new_n3255_));
AND2X2 AND2X2_1421 ( .A(_abc_44694_new_n2972__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_44694_new_n3256_));
AND2X2 AND2X2_1422 ( .A(_abc_44694_new_n1186__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_44694_new_n3259_));
AND2X2 AND2X2_1423 ( .A(_abc_44694_new_n2965__bF_buf1), .B(_abc_44694_new_n3259_), .Y(_abc_44694_new_n3260_));
AND2X2 AND2X2_1424 ( .A(_abc_44694_new_n1185__bF_buf2), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_44694_new_n3261_));
AND2X2 AND2X2_1425 ( .A(_abc_44694_new_n1114__bF_buf4), .B(epc_q_28_), .Y(_abc_44694_new_n3263_));
AND2X2 AND2X2_1426 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n3263_), .Y(_abc_44694_new_n3264_));
AND2X2 AND2X2_1427 ( .A(_abc_44694_new_n3258_), .B(_abc_44694_new_n3266_), .Y(_abc_44694_new_n3267_));
AND2X2 AND2X2_1428 ( .A(_abc_44694_new_n2972__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_44694_new_n3268_));
AND2X2 AND2X2_1429 ( .A(_abc_44694_new_n1186__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_44694_new_n3271_));
AND2X2 AND2X2_143 ( .A(_abc_44694_new_n797_), .B(_abc_44694_new_n870_), .Y(_abc_44694_new_n871_));
AND2X2 AND2X2_1430 ( .A(_abc_44694_new_n2965__bF_buf0), .B(_abc_44694_new_n3271_), .Y(_abc_44694_new_n3272_));
AND2X2 AND2X2_1431 ( .A(_abc_44694_new_n1185__bF_buf1), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_44694_new_n3273_));
AND2X2 AND2X2_1432 ( .A(_abc_44694_new_n1114__bF_buf3), .B(epc_q_29_), .Y(_abc_44694_new_n3275_));
AND2X2 AND2X2_1433 ( .A(_abc_44694_new_n1347__bF_buf3), .B(_abc_44694_new_n3275_), .Y(_abc_44694_new_n3276_));
AND2X2 AND2X2_1434 ( .A(_abc_44694_new_n3270_), .B(_abc_44694_new_n3278_), .Y(_abc_44694_new_n3279_));
AND2X2 AND2X2_1435 ( .A(_abc_44694_new_n2972__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_44694_new_n3280_));
AND2X2 AND2X2_1436 ( .A(_abc_44694_new_n1186__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_44694_new_n3283_));
AND2X2 AND2X2_1437 ( .A(_abc_44694_new_n2965__bF_buf4), .B(_abc_44694_new_n3283_), .Y(_abc_44694_new_n3284_));
AND2X2 AND2X2_1438 ( .A(_abc_44694_new_n1185__bF_buf0), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_44694_new_n3285_));
AND2X2 AND2X2_1439 ( .A(_abc_44694_new_n1114__bF_buf2), .B(epc_q_30_), .Y(_abc_44694_new_n3287_));
AND2X2 AND2X2_144 ( .A(_abc_44694_new_n677__bF_buf2), .B(\mem_dat_i[16] ), .Y(_abc_44694_new_n872_));
AND2X2 AND2X2_1440 ( .A(_abc_44694_new_n1347__bF_buf2), .B(_abc_44694_new_n3287_), .Y(_abc_44694_new_n3288_));
AND2X2 AND2X2_1441 ( .A(_abc_44694_new_n3282_), .B(_abc_44694_new_n3290_), .Y(_abc_44694_new_n3291_));
AND2X2 AND2X2_1442 ( .A(_abc_44694_new_n2972__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_44694_new_n3292_));
AND2X2 AND2X2_1443 ( .A(_abc_44694_new_n1186__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_44694_new_n3295_));
AND2X2 AND2X2_1444 ( .A(_abc_44694_new_n2965__bF_buf3), .B(_abc_44694_new_n3295_), .Y(_abc_44694_new_n3296_));
AND2X2 AND2X2_1445 ( .A(_abc_44694_new_n1185__bF_buf3), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf5_), .Y(_abc_44694_new_n3297_));
AND2X2 AND2X2_1446 ( .A(_abc_44694_new_n1114__bF_buf1), .B(epc_q_31_), .Y(_abc_44694_new_n3299_));
AND2X2 AND2X2_1447 ( .A(_abc_44694_new_n1347__bF_buf1), .B(_abc_44694_new_n3299_), .Y(_abc_44694_new_n3300_));
AND2X2 AND2X2_1448 ( .A(_abc_44694_new_n3294_), .B(_abc_44694_new_n3302_), .Y(_abc_44694_new_n3303_));
AND2X2 AND2X2_1449 ( .A(_abc_44694_new_n2972__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_44694_new_n3304_));
AND2X2 AND2X2_145 ( .A(_abc_44694_new_n873_), .B(_abc_44694_new_n673__bF_buf3), .Y(_abc_44694_new_n874_));
AND2X2 AND2X2_1450 ( .A(_abc_44694_new_n1070_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n3308_));
AND2X2 AND2X2_1451 ( .A(_abc_44694_new_n1055_), .B(_abc_44694_new_n1076_), .Y(_abc_44694_new_n3312_));
AND2X2 AND2X2_1452 ( .A(_abc_44694_new_n1062_), .B(_abc_44694_new_n3312_), .Y(_abc_44694_new_n3313_));
AND2X2 AND2X2_1453 ( .A(_abc_44694_new_n3313_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n3314_));
AND2X2 AND2X2_1454 ( .A(_abc_44694_new_n1061_), .B(_abc_44694_new_n2747_), .Y(_abc_44694_new_n3315_));
AND2X2 AND2X2_1455 ( .A(_abc_44694_new_n1101_), .B(_abc_44694_new_n3315_), .Y(_abc_44694_new_n3316_));
AND2X2 AND2X2_1456 ( .A(_abc_44694_new_n3316_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n3317_));
AND2X2 AND2X2_1457 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .B(alu_op_r_0_), .Y(_abc_44694_new_n3332_));
AND2X2 AND2X2_1458 ( .A(_abc_44694_new_n3333_), .B(_abc_44694_new_n992_), .Y(_abc_44694_new_n3334_));
AND2X2 AND2X2_1459 ( .A(_abc_44694_new_n3335_), .B(_abc_44694_new_n3336_), .Y(_0mem_offset_q_1_0__0_));
AND2X2 AND2X2_146 ( .A(_abc_44694_new_n875_), .B(_abc_44694_new_n876_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_));
AND2X2 AND2X2_1460 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .B(alu_op_r_1_), .Y(_abc_44694_new_n3339_));
AND2X2 AND2X2_1461 ( .A(_abc_44694_new_n3340_), .B(_abc_44694_new_n995_), .Y(_abc_44694_new_n3341_));
AND2X2 AND2X2_1462 ( .A(_abc_44694_new_n3341_), .B(_abc_44694_new_n3332_), .Y(_abc_44694_new_n3342_));
AND2X2 AND2X2_1463 ( .A(_abc_44694_new_n3343_), .B(_abc_44694_new_n3333_), .Y(_abc_44694_new_n3344_));
AND2X2 AND2X2_1464 ( .A(_abc_44694_new_n3347_), .B(_abc_44694_new_n3338_), .Y(_0mem_offset_q_1_0__1_));
AND2X2 AND2X2_1465 ( .A(mem_ack_i), .B(state_q_2_), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424));
AND2X2 AND2X2_1466 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3351_), .Y(_abc_44694_new_n3352_));
AND2X2 AND2X2_1467 ( .A(_abc_44694_new_n3353_), .B(_abc_44694_new_n3350_), .Y(_0opcode_q_31_0__0_));
AND2X2 AND2X2_1468 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3356_), .Y(_abc_44694_new_n3357_));
AND2X2 AND2X2_1469 ( .A(_abc_44694_new_n3358_), .B(_abc_44694_new_n3355_), .Y(_0opcode_q_31_0__1_));
AND2X2 AND2X2_147 ( .A(_abc_44694_new_n677__bF_buf1), .B(\mem_dat_i[17] ), .Y(_abc_44694_new_n878_));
AND2X2 AND2X2_1470 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3361_), .Y(_abc_44694_new_n3362_));
AND2X2 AND2X2_1471 ( .A(_abc_44694_new_n3363_), .B(_abc_44694_new_n3360_), .Y(_0opcode_q_31_0__2_));
AND2X2 AND2X2_1472 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3366_), .Y(_abc_44694_new_n3367_));
AND2X2 AND2X2_1473 ( .A(_abc_44694_new_n3368_), .B(_abc_44694_new_n3365_), .Y(_0opcode_q_31_0__3_));
AND2X2 AND2X2_1474 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3371_), .Y(_abc_44694_new_n3372_));
AND2X2 AND2X2_1475 ( .A(_abc_44694_new_n3373_), .B(_abc_44694_new_n3370_), .Y(_0opcode_q_31_0__4_));
AND2X2 AND2X2_1476 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3376_), .Y(_abc_44694_new_n3377_));
AND2X2 AND2X2_1477 ( .A(_abc_44694_new_n3378_), .B(_abc_44694_new_n3375_), .Y(_0opcode_q_31_0__5_));
AND2X2 AND2X2_1478 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3381_), .Y(_abc_44694_new_n3382_));
AND2X2 AND2X2_1479 ( .A(_abc_44694_new_n3383_), .B(_abc_44694_new_n3380_), .Y(_0opcode_q_31_0__6_));
AND2X2 AND2X2_148 ( .A(_abc_44694_new_n879_), .B(_abc_44694_new_n673__bF_buf2), .Y(_abc_44694_new_n880_));
AND2X2 AND2X2_1480 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3386_), .Y(_abc_44694_new_n3387_));
AND2X2 AND2X2_1481 ( .A(_abc_44694_new_n3388_), .B(_abc_44694_new_n3385_), .Y(_0opcode_q_31_0__7_));
AND2X2 AND2X2_1482 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3391_), .Y(_abc_44694_new_n3392_));
AND2X2 AND2X2_1483 ( .A(_abc_44694_new_n3393_), .B(_abc_44694_new_n3390_), .Y(_0opcode_q_31_0__8_));
AND2X2 AND2X2_1484 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3396_), .Y(_abc_44694_new_n3397_));
AND2X2 AND2X2_1485 ( .A(_abc_44694_new_n3398_), .B(_abc_44694_new_n3395_), .Y(_0opcode_q_31_0__9_));
AND2X2 AND2X2_1486 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3401_), .Y(_abc_44694_new_n3402_));
AND2X2 AND2X2_1487 ( .A(_abc_44694_new_n3403_), .B(_abc_44694_new_n3400_), .Y(_0opcode_q_31_0__10_));
AND2X2 AND2X2_1488 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3406_), .Y(_abc_44694_new_n3407_));
AND2X2 AND2X2_1489 ( .A(_abc_44694_new_n3408_), .B(_abc_44694_new_n3405_), .Y(_0opcode_q_31_0__11_));
AND2X2 AND2X2_149 ( .A(_abc_44694_new_n881_), .B(_abc_44694_new_n882_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_));
AND2X2 AND2X2_1490 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3411_), .Y(_abc_44694_new_n3412_));
AND2X2 AND2X2_1491 ( .A(_abc_44694_new_n3413_), .B(_abc_44694_new_n3410_), .Y(_0opcode_q_31_0__12_));
AND2X2 AND2X2_1492 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3416_), .Y(_abc_44694_new_n3417_));
AND2X2 AND2X2_1493 ( .A(_abc_44694_new_n3418_), .B(_abc_44694_new_n3415_), .Y(_0opcode_q_31_0__13_));
AND2X2 AND2X2_1494 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3421_), .Y(_abc_44694_new_n3422_));
AND2X2 AND2X2_1495 ( .A(_abc_44694_new_n3423_), .B(_abc_44694_new_n3420_), .Y(_0opcode_q_31_0__14_));
AND2X2 AND2X2_1496 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3426_), .Y(_abc_44694_new_n3427_));
AND2X2 AND2X2_1497 ( .A(_abc_44694_new_n3428_), .B(_abc_44694_new_n3425_), .Y(_0opcode_q_31_0__15_));
AND2X2 AND2X2_1498 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3431_), .Y(_abc_44694_new_n3432_));
AND2X2 AND2X2_1499 ( .A(_abc_44694_new_n3433_), .B(_abc_44694_new_n3430_), .Y(_0opcode_q_31_0__16_));
AND2X2 AND2X2_15 ( .A(_abc_44694_new_n639_), .B(_abc_44694_new_n638_), .Y(_abc_44694_new_n640_));
AND2X2 AND2X2_150 ( .A(_abc_44694_new_n677__bF_buf0), .B(\mem_dat_i[18] ), .Y(_abc_44694_new_n884_));
AND2X2 AND2X2_1500 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3436_), .Y(_abc_44694_new_n3437_));
AND2X2 AND2X2_1501 ( .A(_abc_44694_new_n3438_), .B(_abc_44694_new_n3435_), .Y(_0opcode_q_31_0__17_));
AND2X2 AND2X2_1502 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3441_), .Y(_abc_44694_new_n3442_));
AND2X2 AND2X2_1503 ( .A(_abc_44694_new_n3443_), .B(_abc_44694_new_n3440_), .Y(_0opcode_q_31_0__18_));
AND2X2 AND2X2_1504 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3446_), .Y(_abc_44694_new_n3447_));
AND2X2 AND2X2_1505 ( .A(_abc_44694_new_n3448_), .B(_abc_44694_new_n3445_), .Y(_0opcode_q_31_0__19_));
AND2X2 AND2X2_1506 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3451_), .Y(_abc_44694_new_n3452_));
AND2X2 AND2X2_1507 ( .A(_abc_44694_new_n3453_), .B(_abc_44694_new_n3450_), .Y(_0opcode_q_31_0__20_));
AND2X2 AND2X2_1508 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3456_), .Y(_abc_44694_new_n3457_));
AND2X2 AND2X2_1509 ( .A(_abc_44694_new_n3458_), .B(_abc_44694_new_n3455_), .Y(_0opcode_q_31_0__21_));
AND2X2 AND2X2_151 ( .A(_abc_44694_new_n885_), .B(_abc_44694_new_n673__bF_buf1), .Y(_abc_44694_new_n886_));
AND2X2 AND2X2_1510 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3461_), .Y(_abc_44694_new_n3462_));
AND2X2 AND2X2_1511 ( .A(_abc_44694_new_n3463_), .B(_abc_44694_new_n3460_), .Y(_0opcode_q_31_0__22_));
AND2X2 AND2X2_1512 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3466_), .Y(_abc_44694_new_n3467_));
AND2X2 AND2X2_1513 ( .A(_abc_44694_new_n3468_), .B(_abc_44694_new_n3465_), .Y(_0opcode_q_31_0__23_));
AND2X2 AND2X2_1514 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3471_), .Y(_abc_44694_new_n3472_));
AND2X2 AND2X2_1515 ( .A(_abc_44694_new_n3473_), .B(_abc_44694_new_n3470_), .Y(_0opcode_q_31_0__24_));
AND2X2 AND2X2_1516 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3476_), .Y(_abc_44694_new_n3477_));
AND2X2 AND2X2_1517 ( .A(_abc_44694_new_n3478_), .B(_abc_44694_new_n3475_), .Y(_0opcode_q_31_0__25_));
AND2X2 AND2X2_1518 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3481_), .Y(_abc_44694_new_n3482_));
AND2X2 AND2X2_1519 ( .A(_abc_44694_new_n3483_), .B(_abc_44694_new_n3480_), .Y(_0opcode_q_31_0__26_));
AND2X2 AND2X2_152 ( .A(_abc_44694_new_n887_), .B(_abc_44694_new_n888_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_));
AND2X2 AND2X2_1520 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3486_), .Y(_abc_44694_new_n3487_));
AND2X2 AND2X2_1521 ( .A(_abc_44694_new_n3488_), .B(_abc_44694_new_n3485_), .Y(_0opcode_q_31_0__27_));
AND2X2 AND2X2_1522 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6), .B(_abc_44694_new_n3491_), .Y(_abc_44694_new_n3492_));
AND2X2 AND2X2_1523 ( .A(_abc_44694_new_n3493_), .B(_abc_44694_new_n3490_), .Y(_0opcode_q_31_0__28_));
AND2X2 AND2X2_1524 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4), .B(_abc_44694_new_n3496_), .Y(_abc_44694_new_n3497_));
AND2X2 AND2X2_1525 ( .A(_abc_44694_new_n3498_), .B(_abc_44694_new_n3495_), .Y(_0opcode_q_31_0__29_));
AND2X2 AND2X2_1526 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2), .B(_abc_44694_new_n3501_), .Y(_abc_44694_new_n3502_));
AND2X2 AND2X2_1527 ( .A(_abc_44694_new_n3503_), .B(_abc_44694_new_n3500_), .Y(_0opcode_q_31_0__30_));
AND2X2 AND2X2_1528 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0), .B(_abc_44694_new_n3506_), .Y(_abc_44694_new_n3507_));
AND2X2 AND2X2_1529 ( .A(_abc_44694_new_n3508_), .B(_abc_44694_new_n3505_), .Y(_0opcode_q_31_0__31_));
AND2X2 AND2X2_153 ( .A(_abc_44694_new_n677__bF_buf3), .B(\mem_dat_i[19] ), .Y(_abc_44694_new_n890_));
AND2X2 AND2X2_1530 ( .A(_abc_44694_new_n3334__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48783_0_), .Y(_abc_44694_new_n3511_));
AND2X2 AND2X2_1531 ( .A(_abc_44694_new_n634_), .B(_abc_44694_new_n638_), .Y(_abc_44694_new_n3512_));
AND2X2 AND2X2_1532 ( .A(_abc_44694_new_n3346_), .B(_abc_44694_new_n3514_), .Y(_abc_44694_new_n3515_));
AND2X2 AND2X2_1533 ( .A(_abc_44694_new_n634_), .B(_abc_44694_new_n645_), .Y(_abc_44694_new_n3518_));
AND2X2 AND2X2_1534 ( .A(_abc_44694_new_n634_), .B(_abc_44694_new_n647_), .Y(_abc_44694_new_n3520_));
AND2X2 AND2X2_1535 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_abc_44694_new_n3513__bF_buf3), .Y(_abc_44694_new_n3522_));
AND2X2 AND2X2_1536 ( .A(_abc_44694_new_n3524_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3525_));
AND2X2 AND2X2_1537 ( .A(_abc_44694_new_n3517_), .B(_abc_44694_new_n3525_), .Y(_abc_44694_new_n3526_));
AND2X2 AND2X2_1538 ( .A(_abc_44694_new_n654_), .B(state_q_5_bF_buf0_), .Y(_abc_44694_new_n3527_));
AND2X2 AND2X2_1539 ( .A(_abc_44694_new_n3518__bF_buf2), .B(_abc_44694_new_n3334__bF_buf2), .Y(_abc_44694_new_n3529_));
AND2X2 AND2X2_154 ( .A(_abc_44694_new_n891_), .B(_abc_44694_new_n673__bF_buf0), .Y(_abc_44694_new_n892_));
AND2X2 AND2X2_1540 ( .A(_abc_44694_new_n3529_), .B(_abc_44694_new_n3341_), .Y(_abc_44694_new_n3530_));
AND2X2 AND2X2_1541 ( .A(_abc_44694_new_n3532_), .B(_abc_44694_new_n3510_), .Y(_0mem_sel_o_3_0__0_));
AND2X2 AND2X2_1542 ( .A(_abc_44694_new_n3516_), .B(_abc_44694_new_n635_), .Y(_abc_44694_new_n3534_));
AND2X2 AND2X2_1543 ( .A(_abc_44694_new_n3512__bF_buf3), .B(_abc_44694_new_n3514_), .Y(_abc_44694_new_n3536_));
AND2X2 AND2X2_1544 ( .A(_abc_44694_new_n3535_), .B(_abc_44694_new_n3539_), .Y(_abc_44694_new_n3540_));
AND2X2 AND2X2_1545 ( .A(_abc_44694_new_n3541_), .B(_abc_44694_new_n3542_), .Y(_0mem_sel_o_3_0__1_));
AND2X2 AND2X2_1546 ( .A(_abc_44694_new_n3334__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48783_2_), .Y(_abc_44694_new_n3545_));
AND2X2 AND2X2_1547 ( .A(_abc_44694_new_n3345_), .B(_abc_44694_new_n3514_), .Y(_abc_44694_new_n3546_));
AND2X2 AND2X2_1548 ( .A(_abc_44694_new_n3549_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n3550_));
AND2X2 AND2X2_1549 ( .A(_abc_44694_new_n3548_), .B(_abc_44694_new_n3550_), .Y(_abc_44694_new_n3551_));
AND2X2 AND2X2_155 ( .A(_abc_44694_new_n893_), .B(_abc_44694_new_n894_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_));
AND2X2 AND2X2_1550 ( .A(_abc_44694_new_n3529_), .B(_abc_44694_new_n3343_), .Y(_abc_44694_new_n3552_));
AND2X2 AND2X2_1551 ( .A(_abc_44694_new_n3554_), .B(_abc_44694_new_n3544_), .Y(_0mem_sel_o_3_0__2_));
AND2X2 AND2X2_1552 ( .A(_abc_44694_new_n3547_), .B(_abc_44694_new_n635_), .Y(_abc_44694_new_n3556_));
AND2X2 AND2X2_1553 ( .A(_abc_44694_new_n3557_), .B(_abc_44694_new_n3558_), .Y(_abc_44694_new_n3559_));
AND2X2 AND2X2_1554 ( .A(_abc_44694_new_n3560_), .B(_abc_44694_new_n3561_), .Y(_0mem_sel_o_3_0__3_));
AND2X2 AND2X2_1555 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_0_), .Y(_abc_44694_new_n3564_));
AND2X2 AND2X2_1556 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n3565_));
AND2X2 AND2X2_1557 ( .A(_abc_44694_new_n3515__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n3566_));
AND2X2 AND2X2_1558 ( .A(_abc_44694_new_n3334__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_0_), .Y(_abc_44694_new_n3567_));
AND2X2 AND2X2_1559 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_0_), .Y(_abc_44694_new_n3570_));
AND2X2 AND2X2_156 ( .A(_abc_44694_new_n677__bF_buf2), .B(\mem_dat_i[20] ), .Y(_abc_44694_new_n896_));
AND2X2 AND2X2_1560 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n3571_));
AND2X2 AND2X2_1561 ( .A(_abc_44694_new_n3573_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n3574_));
AND2X2 AND2X2_1562 ( .A(_abc_44694_new_n3569_), .B(_abc_44694_new_n3574_), .Y(_abc_44694_new_n3575_));
AND2X2 AND2X2_1563 ( .A(_abc_44694_new_n3576_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n3577_));
AND2X2 AND2X2_1564 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_1_), .Y(_abc_44694_new_n3579_));
AND2X2 AND2X2_1565 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n3580_));
AND2X2 AND2X2_1566 ( .A(_abc_44694_new_n3515__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n3581_));
AND2X2 AND2X2_1567 ( .A(_abc_44694_new_n3334__bF_buf5), .B(_auto_iopadmap_cc_368_execute_48750_1_), .Y(_abc_44694_new_n3582_));
AND2X2 AND2X2_1568 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_1_), .Y(_abc_44694_new_n3585_));
AND2X2 AND2X2_1569 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n3586_));
AND2X2 AND2X2_157 ( .A(_abc_44694_new_n897_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n898_));
AND2X2 AND2X2_1570 ( .A(_abc_44694_new_n3588_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n3589_));
AND2X2 AND2X2_1571 ( .A(_abc_44694_new_n3584_), .B(_abc_44694_new_n3589_), .Y(_abc_44694_new_n3590_));
AND2X2 AND2X2_1572 ( .A(_abc_44694_new_n3591_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n3592_));
AND2X2 AND2X2_1573 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_2_), .Y(_abc_44694_new_n3594_));
AND2X2 AND2X2_1574 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n3595_));
AND2X2 AND2X2_1575 ( .A(_abc_44694_new_n3515__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n3596_));
AND2X2 AND2X2_1576 ( .A(_abc_44694_new_n3334__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_2_), .Y(_abc_44694_new_n3597_));
AND2X2 AND2X2_1577 ( .A(_abc_44694_new_n3521__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_2_), .Y(_abc_44694_new_n3600_));
AND2X2 AND2X2_1578 ( .A(_abc_44694_new_n3520__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n3601_));
AND2X2 AND2X2_1579 ( .A(_abc_44694_new_n3603_), .B(_abc_44694_new_n3519__bF_buf0), .Y(_abc_44694_new_n3604_));
AND2X2 AND2X2_158 ( .A(_abc_44694_new_n899_), .B(_abc_44694_new_n900_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_));
AND2X2 AND2X2_1580 ( .A(_abc_44694_new_n3599_), .B(_abc_44694_new_n3604_), .Y(_abc_44694_new_n3605_));
AND2X2 AND2X2_1581 ( .A(_abc_44694_new_n3606_), .B(_abc_44694_new_n3527__bF_buf1), .Y(_abc_44694_new_n3607_));
AND2X2 AND2X2_1582 ( .A(_abc_44694_new_n3563__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_3_), .Y(_abc_44694_new_n3609_));
AND2X2 AND2X2_1583 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n3610_));
AND2X2 AND2X2_1584 ( .A(_abc_44694_new_n3515__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n3611_));
AND2X2 AND2X2_1585 ( .A(_abc_44694_new_n3334__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_3_), .Y(_abc_44694_new_n3612_));
AND2X2 AND2X2_1586 ( .A(_abc_44694_new_n3521__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_3_), .Y(_abc_44694_new_n3615_));
AND2X2 AND2X2_1587 ( .A(_abc_44694_new_n3520__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n3616_));
AND2X2 AND2X2_1588 ( .A(_abc_44694_new_n3618_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3619_));
AND2X2 AND2X2_1589 ( .A(_abc_44694_new_n3614_), .B(_abc_44694_new_n3619_), .Y(_abc_44694_new_n3620_));
AND2X2 AND2X2_159 ( .A(_abc_44694_new_n677__bF_buf1), .B(\mem_dat_i[21] ), .Y(_abc_44694_new_n902_));
AND2X2 AND2X2_1590 ( .A(_abc_44694_new_n3621_), .B(_abc_44694_new_n3527__bF_buf0), .Y(_abc_44694_new_n3622_));
AND2X2 AND2X2_1591 ( .A(_abc_44694_new_n3563__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_4_), .Y(_abc_44694_new_n3624_));
AND2X2 AND2X2_1592 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n3625_));
AND2X2 AND2X2_1593 ( .A(_abc_44694_new_n3515__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n3626_));
AND2X2 AND2X2_1594 ( .A(_abc_44694_new_n3334__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_4_), .Y(_abc_44694_new_n3627_));
AND2X2 AND2X2_1595 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_4_), .Y(_abc_44694_new_n3630_));
AND2X2 AND2X2_1596 ( .A(_abc_44694_new_n3520__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n3631_));
AND2X2 AND2X2_1597 ( .A(_abc_44694_new_n3633_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n3634_));
AND2X2 AND2X2_1598 ( .A(_abc_44694_new_n3629_), .B(_abc_44694_new_n3634_), .Y(_abc_44694_new_n3635_));
AND2X2 AND2X2_1599 ( .A(_abc_44694_new_n3636_), .B(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n3637_));
AND2X2 AND2X2_16 ( .A(_abc_44694_new_n640_), .B(_abc_44694_new_n637_), .Y(_abc_44694_new_n641_));
AND2X2 AND2X2_160 ( .A(_abc_44694_new_n903_), .B(_abc_44694_new_n673__bF_buf3), .Y(_abc_44694_new_n904_));
AND2X2 AND2X2_1600 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_5_), .Y(_abc_44694_new_n3639_));
AND2X2 AND2X2_1601 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n3640_));
AND2X2 AND2X2_1602 ( .A(_abc_44694_new_n3515__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n3641_));
AND2X2 AND2X2_1603 ( .A(_abc_44694_new_n3334__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_5_), .Y(_abc_44694_new_n3642_));
AND2X2 AND2X2_1604 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_5_), .Y(_abc_44694_new_n3645_));
AND2X2 AND2X2_1605 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n3646_));
AND2X2 AND2X2_1606 ( .A(_abc_44694_new_n3648_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n3649_));
AND2X2 AND2X2_1607 ( .A(_abc_44694_new_n3644_), .B(_abc_44694_new_n3649_), .Y(_abc_44694_new_n3650_));
AND2X2 AND2X2_1608 ( .A(_abc_44694_new_n3651_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n3652_));
AND2X2 AND2X2_1609 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_6_), .Y(_abc_44694_new_n3654_));
AND2X2 AND2X2_161 ( .A(_abc_44694_new_n905_), .B(_abc_44694_new_n906_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_));
AND2X2 AND2X2_1610 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n3655_));
AND2X2 AND2X2_1611 ( .A(_abc_44694_new_n3515__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n3656_));
AND2X2 AND2X2_1612 ( .A(_abc_44694_new_n3334__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_6_), .Y(_abc_44694_new_n3657_));
AND2X2 AND2X2_1613 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_6_), .Y(_abc_44694_new_n3660_));
AND2X2 AND2X2_1614 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n3661_));
AND2X2 AND2X2_1615 ( .A(_abc_44694_new_n3663_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n3664_));
AND2X2 AND2X2_1616 ( .A(_abc_44694_new_n3659_), .B(_abc_44694_new_n3664_), .Y(_abc_44694_new_n3665_));
AND2X2 AND2X2_1617 ( .A(_abc_44694_new_n3666_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n3667_));
AND2X2 AND2X2_1618 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_7_), .Y(_abc_44694_new_n3669_));
AND2X2 AND2X2_1619 ( .A(_abc_44694_new_n3530_), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n3670_));
AND2X2 AND2X2_162 ( .A(_abc_44694_new_n677__bF_buf0), .B(\mem_dat_i[22] ), .Y(_abc_44694_new_n908_));
AND2X2 AND2X2_1620 ( .A(_abc_44694_new_n3515__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n3671_));
AND2X2 AND2X2_1621 ( .A(_abc_44694_new_n3334__bF_buf5), .B(_auto_iopadmap_cc_368_execute_48750_7_), .Y(_abc_44694_new_n3672_));
AND2X2 AND2X2_1622 ( .A(_abc_44694_new_n3521__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_7_), .Y(_abc_44694_new_n3675_));
AND2X2 AND2X2_1623 ( .A(_abc_44694_new_n3520__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n3676_));
AND2X2 AND2X2_1624 ( .A(_abc_44694_new_n3678_), .B(_abc_44694_new_n3519__bF_buf0), .Y(_abc_44694_new_n3679_));
AND2X2 AND2X2_1625 ( .A(_abc_44694_new_n3674_), .B(_abc_44694_new_n3679_), .Y(_abc_44694_new_n3680_));
AND2X2 AND2X2_1626 ( .A(_abc_44694_new_n3681_), .B(_abc_44694_new_n3527__bF_buf1), .Y(_abc_44694_new_n3682_));
AND2X2 AND2X2_1627 ( .A(_abc_44694_new_n3563__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_8_), .Y(_abc_44694_new_n3684_));
AND2X2 AND2X2_1628 ( .A(_abc_44694_new_n3521__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_8_), .Y(_abc_44694_new_n3685_));
AND2X2 AND2X2_1629 ( .A(_abc_44694_new_n3520__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n3686_));
AND2X2 AND2X2_163 ( .A(_abc_44694_new_n909_), .B(_abc_44694_new_n673__bF_buf2), .Y(_abc_44694_new_n910_));
AND2X2 AND2X2_1630 ( .A(_abc_44694_new_n3515__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n3689_));
AND2X2 AND2X2_1631 ( .A(_abc_44694_new_n3334__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_8_), .Y(_abc_44694_new_n3690_));
AND2X2 AND2X2_1632 ( .A(_abc_44694_new_n3692_), .B(_abc_44694_new_n3688_), .Y(_abc_44694_new_n3693_));
AND2X2 AND2X2_1633 ( .A(_abc_44694_new_n3695_), .B(_abc_44694_new_n3527__bF_buf0), .Y(_abc_44694_new_n3696_));
AND2X2 AND2X2_1634 ( .A(_abc_44694_new_n3694_), .B(_abc_44694_new_n3696_), .Y(_abc_44694_new_n3697_));
AND2X2 AND2X2_1635 ( .A(_abc_44694_new_n3563__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_9_), .Y(_abc_44694_new_n3699_));
AND2X2 AND2X2_1636 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_9_), .Y(_abc_44694_new_n3700_));
AND2X2 AND2X2_1637 ( .A(_abc_44694_new_n3520__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n3701_));
AND2X2 AND2X2_1638 ( .A(_abc_44694_new_n3515__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n3704_));
AND2X2 AND2X2_1639 ( .A(_abc_44694_new_n3334__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_9_), .Y(_abc_44694_new_n3705_));
AND2X2 AND2X2_164 ( .A(_abc_44694_new_n911_), .B(_abc_44694_new_n912_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_));
AND2X2 AND2X2_1640 ( .A(_abc_44694_new_n3707_), .B(_abc_44694_new_n3703_), .Y(_abc_44694_new_n3708_));
AND2X2 AND2X2_1641 ( .A(_abc_44694_new_n3710_), .B(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n3711_));
AND2X2 AND2X2_1642 ( .A(_abc_44694_new_n3709_), .B(_abc_44694_new_n3711_), .Y(_abc_44694_new_n3712_));
AND2X2 AND2X2_1643 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_10_), .Y(_abc_44694_new_n3714_));
AND2X2 AND2X2_1644 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_10_), .Y(_abc_44694_new_n3715_));
AND2X2 AND2X2_1645 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n3716_));
AND2X2 AND2X2_1646 ( .A(_abc_44694_new_n3515__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n3719_));
AND2X2 AND2X2_1647 ( .A(_abc_44694_new_n3334__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_10_), .Y(_abc_44694_new_n3720_));
AND2X2 AND2X2_1648 ( .A(_abc_44694_new_n3722_), .B(_abc_44694_new_n3718_), .Y(_abc_44694_new_n3723_));
AND2X2 AND2X2_1649 ( .A(_abc_44694_new_n3725_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n3726_));
AND2X2 AND2X2_165 ( .A(_abc_44694_new_n677__bF_buf3), .B(\mem_dat_i[23] ), .Y(_abc_44694_new_n914_));
AND2X2 AND2X2_1650 ( .A(_abc_44694_new_n3724_), .B(_abc_44694_new_n3726_), .Y(_abc_44694_new_n3727_));
AND2X2 AND2X2_1651 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_11_), .Y(_abc_44694_new_n3729_));
AND2X2 AND2X2_1652 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_11_), .Y(_abc_44694_new_n3730_));
AND2X2 AND2X2_1653 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n3731_));
AND2X2 AND2X2_1654 ( .A(_abc_44694_new_n3515__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n3734_));
AND2X2 AND2X2_1655 ( .A(_abc_44694_new_n3334__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_11_), .Y(_abc_44694_new_n3735_));
AND2X2 AND2X2_1656 ( .A(_abc_44694_new_n3737_), .B(_abc_44694_new_n3733_), .Y(_abc_44694_new_n3738_));
AND2X2 AND2X2_1657 ( .A(_abc_44694_new_n3740_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n3741_));
AND2X2 AND2X2_1658 ( .A(_abc_44694_new_n3739_), .B(_abc_44694_new_n3741_), .Y(_abc_44694_new_n3742_));
AND2X2 AND2X2_1659 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_12_), .Y(_abc_44694_new_n3744_));
AND2X2 AND2X2_166 ( .A(_abc_44694_new_n915_), .B(_abc_44694_new_n673__bF_buf1), .Y(_abc_44694_new_n916_));
AND2X2 AND2X2_1660 ( .A(_abc_44694_new_n3521__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_12_), .Y(_abc_44694_new_n3745_));
AND2X2 AND2X2_1661 ( .A(_abc_44694_new_n3520__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n3746_));
AND2X2 AND2X2_1662 ( .A(_abc_44694_new_n3515__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n3749_));
AND2X2 AND2X2_1663 ( .A(_abc_44694_new_n3334__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_12_), .Y(_abc_44694_new_n3750_));
AND2X2 AND2X2_1664 ( .A(_abc_44694_new_n3752_), .B(_abc_44694_new_n3748_), .Y(_abc_44694_new_n3753_));
AND2X2 AND2X2_1665 ( .A(_abc_44694_new_n3755_), .B(_abc_44694_new_n3527__bF_buf1), .Y(_abc_44694_new_n3756_));
AND2X2 AND2X2_1666 ( .A(_abc_44694_new_n3754_), .B(_abc_44694_new_n3756_), .Y(_abc_44694_new_n3757_));
AND2X2 AND2X2_1667 ( .A(_abc_44694_new_n3563__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_13_), .Y(_abc_44694_new_n3759_));
AND2X2 AND2X2_1668 ( .A(_abc_44694_new_n3521__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_13_), .Y(_abc_44694_new_n3760_));
AND2X2 AND2X2_1669 ( .A(_abc_44694_new_n3520__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n3761_));
AND2X2 AND2X2_167 ( .A(_abc_44694_new_n917_), .B(_abc_44694_new_n918_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_));
AND2X2 AND2X2_1670 ( .A(_abc_44694_new_n3515__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n3764_));
AND2X2 AND2X2_1671 ( .A(_abc_44694_new_n3334__bF_buf5), .B(_auto_iopadmap_cc_368_execute_48750_13_), .Y(_abc_44694_new_n3765_));
AND2X2 AND2X2_1672 ( .A(_abc_44694_new_n3767_), .B(_abc_44694_new_n3763_), .Y(_abc_44694_new_n3768_));
AND2X2 AND2X2_1673 ( .A(_abc_44694_new_n3770_), .B(_abc_44694_new_n3527__bF_buf0), .Y(_abc_44694_new_n3771_));
AND2X2 AND2X2_1674 ( .A(_abc_44694_new_n3769_), .B(_abc_44694_new_n3771_), .Y(_abc_44694_new_n3772_));
AND2X2 AND2X2_1675 ( .A(_abc_44694_new_n3563__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_14_), .Y(_abc_44694_new_n3774_));
AND2X2 AND2X2_1676 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_14_), .Y(_abc_44694_new_n3775_));
AND2X2 AND2X2_1677 ( .A(_abc_44694_new_n3520__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n3776_));
AND2X2 AND2X2_1678 ( .A(_abc_44694_new_n3515__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n3779_));
AND2X2 AND2X2_1679 ( .A(_abc_44694_new_n3334__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_14_), .Y(_abc_44694_new_n3780_));
AND2X2 AND2X2_168 ( .A(_abc_44694_new_n677__bF_buf2), .B(\mem_dat_i[24] ), .Y(_abc_44694_new_n920_));
AND2X2 AND2X2_1680 ( .A(_abc_44694_new_n3782_), .B(_abc_44694_new_n3778_), .Y(_abc_44694_new_n3783_));
AND2X2 AND2X2_1681 ( .A(_abc_44694_new_n3785_), .B(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n3786_));
AND2X2 AND2X2_1682 ( .A(_abc_44694_new_n3784_), .B(_abc_44694_new_n3786_), .Y(_abc_44694_new_n3787_));
AND2X2 AND2X2_1683 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_15_), .Y(_abc_44694_new_n3789_));
AND2X2 AND2X2_1684 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_15_), .Y(_abc_44694_new_n3790_));
AND2X2 AND2X2_1685 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n3791_));
AND2X2 AND2X2_1686 ( .A(_abc_44694_new_n3515__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n3794_));
AND2X2 AND2X2_1687 ( .A(_abc_44694_new_n3334__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_15_), .Y(_abc_44694_new_n3795_));
AND2X2 AND2X2_1688 ( .A(_abc_44694_new_n3797_), .B(_abc_44694_new_n3793_), .Y(_abc_44694_new_n3798_));
AND2X2 AND2X2_1689 ( .A(_abc_44694_new_n3800_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n3801_));
AND2X2 AND2X2_169 ( .A(_abc_44694_new_n921_), .B(_abc_44694_new_n673__bF_buf0), .Y(_abc_44694_new_n922_));
AND2X2 AND2X2_1690 ( .A(_abc_44694_new_n3799_), .B(_abc_44694_new_n3801_), .Y(_abc_44694_new_n3802_));
AND2X2 AND2X2_1691 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_16_), .Y(_abc_44694_new_n3804_));
AND2X2 AND2X2_1692 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n3805_));
AND2X2 AND2X2_1693 ( .A(_abc_44694_new_n3546__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n3806_));
AND2X2 AND2X2_1694 ( .A(_abc_44694_new_n3334__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_16_), .Y(_abc_44694_new_n3807_));
AND2X2 AND2X2_1695 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_16_), .Y(_abc_44694_new_n3810_));
AND2X2 AND2X2_1696 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_44694_new_n3811_));
AND2X2 AND2X2_1697 ( .A(_abc_44694_new_n3813_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n3814_));
AND2X2 AND2X2_1698 ( .A(_abc_44694_new_n3809_), .B(_abc_44694_new_n3814_), .Y(_abc_44694_new_n3815_));
AND2X2 AND2X2_1699 ( .A(_abc_44694_new_n3816_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n3817_));
AND2X2 AND2X2_17 ( .A(_abc_44694_new_n626_), .B(_abc_44694_new_n632_), .Y(_abc_44694_new_n642_));
AND2X2 AND2X2_170 ( .A(_abc_44694_new_n923_), .B(_abc_44694_new_n924_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_));
AND2X2 AND2X2_1700 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_17_), .Y(_abc_44694_new_n3819_));
AND2X2 AND2X2_1701 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n3820_));
AND2X2 AND2X2_1702 ( .A(_abc_44694_new_n3546__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n3821_));
AND2X2 AND2X2_1703 ( .A(_abc_44694_new_n3334__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_17_), .Y(_abc_44694_new_n3822_));
AND2X2 AND2X2_1704 ( .A(_abc_44694_new_n3521__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_17_), .Y(_abc_44694_new_n3825_));
AND2X2 AND2X2_1705 ( .A(_abc_44694_new_n3520__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_44694_new_n3826_));
AND2X2 AND2X2_1706 ( .A(_abc_44694_new_n3828_), .B(_abc_44694_new_n3519__bF_buf0), .Y(_abc_44694_new_n3829_));
AND2X2 AND2X2_1707 ( .A(_abc_44694_new_n3824_), .B(_abc_44694_new_n3829_), .Y(_abc_44694_new_n3830_));
AND2X2 AND2X2_1708 ( .A(_abc_44694_new_n3831_), .B(_abc_44694_new_n3527__bF_buf1), .Y(_abc_44694_new_n3832_));
AND2X2 AND2X2_1709 ( .A(_abc_44694_new_n3563__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_18_), .Y(_abc_44694_new_n3834_));
AND2X2 AND2X2_171 ( .A(_abc_44694_new_n677__bF_buf1), .B(\mem_dat_i[25] ), .Y(_abc_44694_new_n926_));
AND2X2 AND2X2_1710 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n3835_));
AND2X2 AND2X2_1711 ( .A(_abc_44694_new_n3546__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n3836_));
AND2X2 AND2X2_1712 ( .A(_abc_44694_new_n3334__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_18_), .Y(_abc_44694_new_n3837_));
AND2X2 AND2X2_1713 ( .A(_abc_44694_new_n3521__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_18_), .Y(_abc_44694_new_n3840_));
AND2X2 AND2X2_1714 ( .A(_abc_44694_new_n3520__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_44694_new_n3841_));
AND2X2 AND2X2_1715 ( .A(_abc_44694_new_n3843_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3844_));
AND2X2 AND2X2_1716 ( .A(_abc_44694_new_n3839_), .B(_abc_44694_new_n3844_), .Y(_abc_44694_new_n3845_));
AND2X2 AND2X2_1717 ( .A(_abc_44694_new_n3846_), .B(_abc_44694_new_n3527__bF_buf0), .Y(_abc_44694_new_n3847_));
AND2X2 AND2X2_1718 ( .A(_abc_44694_new_n3563__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_19_), .Y(_abc_44694_new_n3849_));
AND2X2 AND2X2_1719 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n3850_));
AND2X2 AND2X2_172 ( .A(_abc_44694_new_n927_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n928_));
AND2X2 AND2X2_1720 ( .A(_abc_44694_new_n3546__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n3851_));
AND2X2 AND2X2_1721 ( .A(_abc_44694_new_n3334__bF_buf5), .B(_auto_iopadmap_cc_368_execute_48750_19_), .Y(_abc_44694_new_n3852_));
AND2X2 AND2X2_1722 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_19_), .Y(_abc_44694_new_n3855_));
AND2X2 AND2X2_1723 ( .A(_abc_44694_new_n3520__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_44694_new_n3856_));
AND2X2 AND2X2_1724 ( .A(_abc_44694_new_n3858_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n3859_));
AND2X2 AND2X2_1725 ( .A(_abc_44694_new_n3854_), .B(_abc_44694_new_n3859_), .Y(_abc_44694_new_n3860_));
AND2X2 AND2X2_1726 ( .A(_abc_44694_new_n3861_), .B(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n3862_));
AND2X2 AND2X2_1727 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_20_), .Y(_abc_44694_new_n3864_));
AND2X2 AND2X2_1728 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n3865_));
AND2X2 AND2X2_1729 ( .A(_abc_44694_new_n3546__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n3866_));
AND2X2 AND2X2_173 ( .A(_abc_44694_new_n929_), .B(_abc_44694_new_n930_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_));
AND2X2 AND2X2_1730 ( .A(_abc_44694_new_n3334__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_20_), .Y(_abc_44694_new_n3867_));
AND2X2 AND2X2_1731 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_20_), .Y(_abc_44694_new_n3870_));
AND2X2 AND2X2_1732 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_44694_new_n3871_));
AND2X2 AND2X2_1733 ( .A(_abc_44694_new_n3873_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n3874_));
AND2X2 AND2X2_1734 ( .A(_abc_44694_new_n3869_), .B(_abc_44694_new_n3874_), .Y(_abc_44694_new_n3875_));
AND2X2 AND2X2_1735 ( .A(_abc_44694_new_n3876_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n3877_));
AND2X2 AND2X2_1736 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_21_), .Y(_abc_44694_new_n3879_));
AND2X2 AND2X2_1737 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n3880_));
AND2X2 AND2X2_1738 ( .A(_abc_44694_new_n3546__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n3881_));
AND2X2 AND2X2_1739 ( .A(_abc_44694_new_n3334__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_21_), .Y(_abc_44694_new_n3882_));
AND2X2 AND2X2_174 ( .A(_abc_44694_new_n677__bF_buf0), .B(\mem_dat_i[26] ), .Y(_abc_44694_new_n932_));
AND2X2 AND2X2_1740 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_21_), .Y(_abc_44694_new_n3885_));
AND2X2 AND2X2_1741 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_44694_new_n3886_));
AND2X2 AND2X2_1742 ( .A(_abc_44694_new_n3888_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n3889_));
AND2X2 AND2X2_1743 ( .A(_abc_44694_new_n3884_), .B(_abc_44694_new_n3889_), .Y(_abc_44694_new_n3890_));
AND2X2 AND2X2_1744 ( .A(_abc_44694_new_n3891_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n3892_));
AND2X2 AND2X2_1745 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_22_), .Y(_abc_44694_new_n3894_));
AND2X2 AND2X2_1746 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n3895_));
AND2X2 AND2X2_1747 ( .A(_abc_44694_new_n3546__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n3896_));
AND2X2 AND2X2_1748 ( .A(_abc_44694_new_n3334__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_22_), .Y(_abc_44694_new_n3897_));
AND2X2 AND2X2_1749 ( .A(_abc_44694_new_n3521__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_22_), .Y(_abc_44694_new_n3900_));
AND2X2 AND2X2_175 ( .A(_abc_44694_new_n933_), .B(_abc_44694_new_n673__bF_buf3), .Y(_abc_44694_new_n934_));
AND2X2 AND2X2_1750 ( .A(_abc_44694_new_n3520__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_44694_new_n3901_));
AND2X2 AND2X2_1751 ( .A(_abc_44694_new_n3903_), .B(_abc_44694_new_n3519__bF_buf0), .Y(_abc_44694_new_n3904_));
AND2X2 AND2X2_1752 ( .A(_abc_44694_new_n3899_), .B(_abc_44694_new_n3904_), .Y(_abc_44694_new_n3905_));
AND2X2 AND2X2_1753 ( .A(_abc_44694_new_n3906_), .B(_abc_44694_new_n3527__bF_buf1), .Y(_abc_44694_new_n3907_));
AND2X2 AND2X2_1754 ( .A(_abc_44694_new_n3563__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_23_), .Y(_abc_44694_new_n3909_));
AND2X2 AND2X2_1755 ( .A(_abc_44694_new_n3552_), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n3910_));
AND2X2 AND2X2_1756 ( .A(_abc_44694_new_n3546__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n3911_));
AND2X2 AND2X2_1757 ( .A(_abc_44694_new_n3334__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_23_), .Y(_abc_44694_new_n3912_));
AND2X2 AND2X2_1758 ( .A(_abc_44694_new_n3521__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_23_), .Y(_abc_44694_new_n3915_));
AND2X2 AND2X2_1759 ( .A(_abc_44694_new_n3520__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_44694_new_n3916_));
AND2X2 AND2X2_176 ( .A(_abc_44694_new_n935_), .B(_abc_44694_new_n936_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_));
AND2X2 AND2X2_1760 ( .A(_abc_44694_new_n3918_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3919_));
AND2X2 AND2X2_1761 ( .A(_abc_44694_new_n3914_), .B(_abc_44694_new_n3919_), .Y(_abc_44694_new_n3920_));
AND2X2 AND2X2_1762 ( .A(_abc_44694_new_n3921_), .B(_abc_44694_new_n3527__bF_buf0), .Y(_abc_44694_new_n3922_));
AND2X2 AND2X2_1763 ( .A(_abc_44694_new_n3563__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_24_), .Y(_abc_44694_new_n3924_));
AND2X2 AND2X2_1764 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_24_), .Y(_abc_44694_new_n3925_));
AND2X2 AND2X2_1765 ( .A(_abc_44694_new_n3520__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_44694_new_n3926_));
AND2X2 AND2X2_1766 ( .A(_abc_44694_new_n3546__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n3929_));
AND2X2 AND2X2_1767 ( .A(_abc_44694_new_n3334__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_24_), .Y(_abc_44694_new_n3930_));
AND2X2 AND2X2_1768 ( .A(_abc_44694_new_n3932_), .B(_abc_44694_new_n3928_), .Y(_abc_44694_new_n3933_));
AND2X2 AND2X2_1769 ( .A(_abc_44694_new_n3935_), .B(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n3936_));
AND2X2 AND2X2_177 ( .A(_abc_44694_new_n677__bF_buf3), .B(\mem_dat_i[27] ), .Y(_abc_44694_new_n938_));
AND2X2 AND2X2_1770 ( .A(_abc_44694_new_n3934_), .B(_abc_44694_new_n3936_), .Y(_abc_44694_new_n3937_));
AND2X2 AND2X2_1771 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_25_), .Y(_abc_44694_new_n3939_));
AND2X2 AND2X2_1772 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_25_), .Y(_abc_44694_new_n3940_));
AND2X2 AND2X2_1773 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_44694_new_n3941_));
AND2X2 AND2X2_1774 ( .A(_abc_44694_new_n3546__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n3944_));
AND2X2 AND2X2_1775 ( .A(_abc_44694_new_n3334__bF_buf5), .B(_auto_iopadmap_cc_368_execute_48750_25_), .Y(_abc_44694_new_n3945_));
AND2X2 AND2X2_1776 ( .A(_abc_44694_new_n3947_), .B(_abc_44694_new_n3943_), .Y(_abc_44694_new_n3948_));
AND2X2 AND2X2_1777 ( .A(_abc_44694_new_n3950_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n3951_));
AND2X2 AND2X2_1778 ( .A(_abc_44694_new_n3949_), .B(_abc_44694_new_n3951_), .Y(_abc_44694_new_n3952_));
AND2X2 AND2X2_1779 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_26_), .Y(_abc_44694_new_n3954_));
AND2X2 AND2X2_178 ( .A(_abc_44694_new_n939_), .B(_abc_44694_new_n673__bF_buf2), .Y(_abc_44694_new_n940_));
AND2X2 AND2X2_1780 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_26_), .Y(_abc_44694_new_n3955_));
AND2X2 AND2X2_1781 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_44694_new_n3956_));
AND2X2 AND2X2_1782 ( .A(_abc_44694_new_n3546__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n3959_));
AND2X2 AND2X2_1783 ( .A(_abc_44694_new_n3334__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_26_), .Y(_abc_44694_new_n3960_));
AND2X2 AND2X2_1784 ( .A(_abc_44694_new_n3962_), .B(_abc_44694_new_n3958_), .Y(_abc_44694_new_n3963_));
AND2X2 AND2X2_1785 ( .A(_abc_44694_new_n3965_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n3966_));
AND2X2 AND2X2_1786 ( .A(_abc_44694_new_n3964_), .B(_abc_44694_new_n3966_), .Y(_abc_44694_new_n3967_));
AND2X2 AND2X2_1787 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_27_), .Y(_abc_44694_new_n3969_));
AND2X2 AND2X2_1788 ( .A(_abc_44694_new_n3521__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_27_), .Y(_abc_44694_new_n3970_));
AND2X2 AND2X2_1789 ( .A(_abc_44694_new_n3520__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_44694_new_n3971_));
AND2X2 AND2X2_179 ( .A(_abc_44694_new_n941_), .B(_abc_44694_new_n942_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_));
AND2X2 AND2X2_1790 ( .A(_abc_44694_new_n3546__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n3974_));
AND2X2 AND2X2_1791 ( .A(_abc_44694_new_n3334__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_27_), .Y(_abc_44694_new_n3975_));
AND2X2 AND2X2_1792 ( .A(_abc_44694_new_n3977_), .B(_abc_44694_new_n3973_), .Y(_abc_44694_new_n3978_));
AND2X2 AND2X2_1793 ( .A(_abc_44694_new_n3980_), .B(_abc_44694_new_n3527__bF_buf1), .Y(_abc_44694_new_n3981_));
AND2X2 AND2X2_1794 ( .A(_abc_44694_new_n3979_), .B(_abc_44694_new_n3981_), .Y(_abc_44694_new_n3982_));
AND2X2 AND2X2_1795 ( .A(_abc_44694_new_n3563__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_28_), .Y(_abc_44694_new_n3984_));
AND2X2 AND2X2_1796 ( .A(_abc_44694_new_n3521__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_28_), .Y(_abc_44694_new_n3985_));
AND2X2 AND2X2_1797 ( .A(_abc_44694_new_n3520__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_44694_new_n3986_));
AND2X2 AND2X2_1798 ( .A(_abc_44694_new_n3546__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n3989_));
AND2X2 AND2X2_1799 ( .A(_abc_44694_new_n3334__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_28_), .Y(_abc_44694_new_n3990_));
AND2X2 AND2X2_18 ( .A(_abc_44694_new_n642_), .B(_abc_44694_new_n637_), .Y(_abc_44694_new_n643_));
AND2X2 AND2X2_180 ( .A(_abc_44694_new_n677__bF_buf2), .B(\mem_dat_i[28] ), .Y(_abc_44694_new_n944_));
AND2X2 AND2X2_1800 ( .A(_abc_44694_new_n3992_), .B(_abc_44694_new_n3988_), .Y(_abc_44694_new_n3993_));
AND2X2 AND2X2_1801 ( .A(_abc_44694_new_n3995_), .B(_abc_44694_new_n3527__bF_buf0), .Y(_abc_44694_new_n3996_));
AND2X2 AND2X2_1802 ( .A(_abc_44694_new_n3994_), .B(_abc_44694_new_n3996_), .Y(_abc_44694_new_n3997_));
AND2X2 AND2X2_1803 ( .A(_abc_44694_new_n3563__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_29_), .Y(_abc_44694_new_n3999_));
AND2X2 AND2X2_1804 ( .A(_abc_44694_new_n3521__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_29_), .Y(_abc_44694_new_n4000_));
AND2X2 AND2X2_1805 ( .A(_abc_44694_new_n3520__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_44694_new_n4001_));
AND2X2 AND2X2_1806 ( .A(_abc_44694_new_n3546__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n4004_));
AND2X2 AND2X2_1807 ( .A(_abc_44694_new_n3334__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48750_29_), .Y(_abc_44694_new_n4005_));
AND2X2 AND2X2_1808 ( .A(_abc_44694_new_n4007_), .B(_abc_44694_new_n4003_), .Y(_abc_44694_new_n4008_));
AND2X2 AND2X2_1809 ( .A(_abc_44694_new_n4010_), .B(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n4011_));
AND2X2 AND2X2_181 ( .A(_abc_44694_new_n945_), .B(_abc_44694_new_n673__bF_buf1), .Y(_abc_44694_new_n946_));
AND2X2 AND2X2_1810 ( .A(_abc_44694_new_n4009_), .B(_abc_44694_new_n4011_), .Y(_abc_44694_new_n4012_));
AND2X2 AND2X2_1811 ( .A(_abc_44694_new_n3563__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48750_30_), .Y(_abc_44694_new_n4014_));
AND2X2 AND2X2_1812 ( .A(_abc_44694_new_n3521__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_30_), .Y(_abc_44694_new_n4015_));
AND2X2 AND2X2_1813 ( .A(_abc_44694_new_n3520__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_44694_new_n4016_));
AND2X2 AND2X2_1814 ( .A(_abc_44694_new_n3546__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n4019_));
AND2X2 AND2X2_1815 ( .A(_abc_44694_new_n3334__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48750_30_), .Y(_abc_44694_new_n4020_));
AND2X2 AND2X2_1816 ( .A(_abc_44694_new_n4022_), .B(_abc_44694_new_n4018_), .Y(_abc_44694_new_n4023_));
AND2X2 AND2X2_1817 ( .A(_abc_44694_new_n4025_), .B(_abc_44694_new_n3527__bF_buf3), .Y(_abc_44694_new_n4026_));
AND2X2 AND2X2_1818 ( .A(_abc_44694_new_n4024_), .B(_abc_44694_new_n4026_), .Y(_abc_44694_new_n4027_));
AND2X2 AND2X2_1819 ( .A(_abc_44694_new_n3563__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48750_31_), .Y(_abc_44694_new_n4029_));
AND2X2 AND2X2_182 ( .A(_abc_44694_new_n947_), .B(_abc_44694_new_n948_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_));
AND2X2 AND2X2_1820 ( .A(_abc_44694_new_n3521__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48750_31_), .Y(_abc_44694_new_n4030_));
AND2X2 AND2X2_1821 ( .A(_abc_44694_new_n3520__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_44694_new_n4031_));
AND2X2 AND2X2_1822 ( .A(_abc_44694_new_n3546__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n4034_));
AND2X2 AND2X2_1823 ( .A(_abc_44694_new_n3334__bF_buf5), .B(_auto_iopadmap_cc_368_execute_48750_31_), .Y(_abc_44694_new_n4035_));
AND2X2 AND2X2_1824 ( .A(_abc_44694_new_n4037_), .B(_abc_44694_new_n4033_), .Y(_abc_44694_new_n4038_));
AND2X2 AND2X2_1825 ( .A(_abc_44694_new_n4040_), .B(_abc_44694_new_n3527__bF_buf2), .Y(_abc_44694_new_n4041_));
AND2X2 AND2X2_1826 ( .A(_abc_44694_new_n4039_), .B(_abc_44694_new_n4041_), .Y(_abc_44694_new_n4042_));
AND2X2 AND2X2_1827 ( .A(_abc_44694_new_n3563__bF_buf2), .B(_abc_44694_new_n4046_), .Y(_abc_44694_new_n4047_));
AND2X2 AND2X2_1828 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48790), .Y(_abc_44694_new_n4048_));
AND2X2 AND2X2_1829 ( .A(_abc_44694_new_n4049_), .B(_abc_44694_new_n4045_), .Y(_0mem_we_o_0_0_));
AND2X2 AND2X2_183 ( .A(_abc_44694_new_n677__bF_buf1), .B(\mem_dat_i[29] ), .Y(_abc_44694_new_n950_));
AND2X2 AND2X2_1830 ( .A(_abc_44694_new_n4051_), .B(state_q_5_bF_buf3_), .Y(_abc_44694_new_n4052_));
AND2X2 AND2X2_1831 ( .A(_auto_iopadmap_cc_368_execute_48788), .B(mem_stall_i), .Y(_abc_44694_new_n4053_));
AND2X2 AND2X2_1832 ( .A(_abc_44694_new_n671_), .B(_abc_44694_new_n4056_), .Y(_abc_44694_new_n4057_));
AND2X2 AND2X2_1833 ( .A(_abc_44694_new_n4059_), .B(_auto_iopadmap_cc_368_execute_48748), .Y(_abc_44694_new_n4060_));
AND2X2 AND2X2_1834 ( .A(state_q_3_bF_buf1_), .B(next_pc_r_0_), .Y(_abc_44694_new_n4063_));
AND2X2 AND2X2_1835 ( .A(_abc_44694_new_n4064__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48711_0_), .Y(_abc_44694_new_n4065_));
AND2X2 AND2X2_1836 ( .A(state_q_3_bF_buf0_), .B(next_pc_r_1_), .Y(_abc_44694_new_n4067_));
AND2X2 AND2X2_1837 ( .A(_abc_44694_new_n4064__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48711_1_), .Y(_abc_44694_new_n4068_));
AND2X2 AND2X2_1838 ( .A(_abc_44694_new_n4064__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48711_2_), .Y(_abc_44694_new_n4070_));
AND2X2 AND2X2_1839 ( .A(state_q_3_bF_buf5_), .B(pc_q_2_), .Y(_abc_44694_new_n4071_));
AND2X2 AND2X2_184 ( .A(_abc_44694_new_n951_), .B(_abc_44694_new_n673__bF_buf0), .Y(_abc_44694_new_n952_));
AND2X2 AND2X2_1840 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_2_), .B(alu_op_r_2_), .Y(_abc_44694_new_n4073_));
AND2X2 AND2X2_1841 ( .A(_abc_44694_new_n4074_), .B(_abc_44694_new_n1006_), .Y(_abc_44694_new_n4075_));
AND2X2 AND2X2_1842 ( .A(_abc_44694_new_n4072_), .B(_abc_44694_new_n4075_), .Y(_abc_44694_new_n4076_));
AND2X2 AND2X2_1843 ( .A(_abc_44694_new_n4077_), .B(_abc_44694_new_n4078_), .Y(_abc_44694_new_n4079_));
AND2X2 AND2X2_1844 ( .A(_abc_44694_new_n668__bF_buf0), .B(_abc_44694_new_n4079_), .Y(_abc_44694_new_n4080_));
AND2X2 AND2X2_1845 ( .A(_abc_44694_new_n4064__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48711_3_), .Y(_abc_44694_new_n4083_));
AND2X2 AND2X2_1846 ( .A(state_q_3_bF_buf4_), .B(pc_q_3_), .Y(_abc_44694_new_n4084_));
AND2X2 AND2X2_1847 ( .A(_abc_44694_new_n4077_), .B(_abc_44694_new_n4074_), .Y(_abc_44694_new_n4085_));
AND2X2 AND2X2_1848 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_3_), .B(alu_op_r_3_), .Y(_abc_44694_new_n4087_));
AND2X2 AND2X2_1849 ( .A(_abc_44694_new_n4088_), .B(_abc_44694_new_n1004_), .Y(_abc_44694_new_n4089_));
AND2X2 AND2X2_185 ( .A(_abc_44694_new_n953_), .B(_abc_44694_new_n954_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_));
AND2X2 AND2X2_1850 ( .A(_abc_44694_new_n4090_), .B(_abc_44694_new_n4092_), .Y(_abc_44694_new_n4093_));
AND2X2 AND2X2_1851 ( .A(_abc_44694_new_n4093_), .B(_abc_44694_new_n668__bF_buf4), .Y(_abc_44694_new_n4094_));
AND2X2 AND2X2_1852 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_4_), .B(int32_r_4_), .Y(_abc_44694_new_n4097_));
AND2X2 AND2X2_1853 ( .A(_abc_44694_new_n4098_), .B(_abc_44694_new_n994_), .Y(_abc_44694_new_n4099_));
AND2X2 AND2X2_1854 ( .A(_abc_44694_new_n4100_), .B(_abc_44694_new_n4088_), .Y(_abc_44694_new_n4101_));
AND2X2 AND2X2_1855 ( .A(_abc_44694_new_n4105_), .B(_abc_44694_new_n668__bF_buf3), .Y(_abc_44694_new_n4106_));
AND2X2 AND2X2_1856 ( .A(_abc_44694_new_n4106_), .B(_abc_44694_new_n4103_), .Y(_abc_44694_new_n4107_));
AND2X2 AND2X2_1857 ( .A(state_q_3_bF_buf3_), .B(pc_q_4_), .Y(_abc_44694_new_n4108_));
AND2X2 AND2X2_1858 ( .A(_abc_44694_new_n4064__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48711_4_), .Y(_abc_44694_new_n4109_));
AND2X2 AND2X2_1859 ( .A(_abc_44694_new_n4105_), .B(_abc_44694_new_n4098_), .Y(_abc_44694_new_n4112_));
AND2X2 AND2X2_186 ( .A(_abc_44694_new_n677__bF_buf0), .B(\mem_dat_i[30] ), .Y(_abc_44694_new_n956_));
AND2X2 AND2X2_1860 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_5_), .B(int32_r_5_), .Y(_abc_44694_new_n4113_));
AND2X2 AND2X2_1861 ( .A(_abc_44694_new_n4114_), .B(_abc_44694_new_n990_), .Y(_abc_44694_new_n4115_));
AND2X2 AND2X2_1862 ( .A(_abc_44694_new_n4119_), .B(_abc_44694_new_n668__bF_buf2), .Y(_abc_44694_new_n4120_));
AND2X2 AND2X2_1863 ( .A(_abc_44694_new_n4120_), .B(_abc_44694_new_n4117_), .Y(_abc_44694_new_n4121_));
AND2X2 AND2X2_1864 ( .A(state_q_3_bF_buf2_), .B(pc_q_5_), .Y(_abc_44694_new_n4122_));
AND2X2 AND2X2_1865 ( .A(_abc_44694_new_n4064__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48711_5_), .Y(_abc_44694_new_n4123_));
AND2X2 AND2X2_1866 ( .A(_abc_44694_new_n4117_), .B(_abc_44694_new_n4114_), .Y(_abc_44694_new_n4126_));
AND2X2 AND2X2_1867 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_6_), .B(alu_op_r_4_), .Y(_abc_44694_new_n4128_));
AND2X2 AND2X2_1868 ( .A(_abc_44694_new_n4129_), .B(_abc_44694_new_n1001_), .Y(_abc_44694_new_n4130_));
AND2X2 AND2X2_1869 ( .A(_abc_44694_new_n4127_), .B(_abc_44694_new_n4130_), .Y(_abc_44694_new_n4132_));
AND2X2 AND2X2_187 ( .A(_abc_44694_new_n957_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n958_));
AND2X2 AND2X2_1870 ( .A(_abc_44694_new_n4133_), .B(_abc_44694_new_n4131_), .Y(_abc_44694_new_n4134_));
AND2X2 AND2X2_1871 ( .A(_abc_44694_new_n4134_), .B(_abc_44694_new_n668__bF_buf1), .Y(_abc_44694_new_n4135_));
AND2X2 AND2X2_1872 ( .A(state_q_3_bF_buf1_), .B(pc_q_6_), .Y(_abc_44694_new_n4136_));
AND2X2 AND2X2_1873 ( .A(_abc_44694_new_n4064__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48711_6_), .Y(_abc_44694_new_n4137_));
AND2X2 AND2X2_1874 ( .A(state_q_5_bF_buf1_), .B(_auto_iopadmap_cc_368_execute_48711_7_), .Y(_abc_44694_new_n4140_));
AND2X2 AND2X2_1875 ( .A(_abc_44694_new_n4133_), .B(_abc_44694_new_n4129_), .Y(_abc_44694_new_n4142_));
AND2X2 AND2X2_1876 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_7_), .B(alu_op_r_5_), .Y(_abc_44694_new_n4144_));
AND2X2 AND2X2_1877 ( .A(_abc_44694_new_n4145_), .B(_abc_44694_new_n999_), .Y(_abc_44694_new_n4146_));
AND2X2 AND2X2_1878 ( .A(_abc_44694_new_n4143_), .B(_abc_44694_new_n4147_), .Y(_abc_44694_new_n4148_));
AND2X2 AND2X2_1879 ( .A(_abc_44694_new_n4142_), .B(_abc_44694_new_n4146_), .Y(_abc_44694_new_n4149_));
AND2X2 AND2X2_188 ( .A(_abc_44694_new_n959_), .B(_abc_44694_new_n960_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_));
AND2X2 AND2X2_1880 ( .A(_abc_44694_new_n4151_), .B(_abc_44694_new_n4141_), .Y(_abc_44694_new_n4152_));
AND2X2 AND2X2_1881 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_7_), .Y(_abc_44694_new_n4153_));
AND2X2 AND2X2_1882 ( .A(state_q_3_bF_buf0_), .B(pc_q_7_), .Y(_abc_44694_new_n4154_));
AND2X2 AND2X2_1883 ( .A(_abc_44694_new_n999_), .B(_abc_44694_new_n4128_), .Y(_abc_44694_new_n4157_));
AND2X2 AND2X2_1884 ( .A(_abc_44694_new_n4130_), .B(_abc_44694_new_n4146_), .Y(_abc_44694_new_n4160_));
AND2X2 AND2X2_1885 ( .A(_abc_44694_new_n4162_), .B(_abc_44694_new_n4159_), .Y(_abc_44694_new_n4163_));
AND2X2 AND2X2_1886 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_8_), .B(alu_op_r_6_), .Y(_abc_44694_new_n4165_));
AND2X2 AND2X2_1887 ( .A(_abc_44694_new_n4166_), .B(_abc_44694_new_n972_), .Y(_abc_44694_new_n4167_));
AND2X2 AND2X2_1888 ( .A(_abc_44694_new_n4164_), .B(_abc_44694_new_n4167_), .Y(_abc_44694_new_n4169_));
AND2X2 AND2X2_1889 ( .A(_abc_44694_new_n4170_), .B(_abc_44694_new_n4168_), .Y(_abc_44694_new_n4171_));
AND2X2 AND2X2_189 ( .A(_abc_44694_new_n677__bF_buf3), .B(\mem_dat_i[31] ), .Y(_abc_44694_new_n962_));
AND2X2 AND2X2_1890 ( .A(_abc_44694_new_n4171_), .B(_abc_44694_new_n668__bF_buf4), .Y(_abc_44694_new_n4172_));
AND2X2 AND2X2_1891 ( .A(state_q_3_bF_buf5_), .B(pc_q_8_), .Y(_abc_44694_new_n4173_));
AND2X2 AND2X2_1892 ( .A(_abc_44694_new_n4064__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48711_8_), .Y(_abc_44694_new_n4174_));
AND2X2 AND2X2_1893 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_9_), .B(alu_op_r_7_), .Y(_abc_44694_new_n4177_));
AND2X2 AND2X2_1894 ( .A(_abc_44694_new_n4178_), .B(_abc_44694_new_n974_), .Y(_abc_44694_new_n4179_));
AND2X2 AND2X2_1895 ( .A(_abc_44694_new_n4170_), .B(_abc_44694_new_n4166_), .Y(_abc_44694_new_n4180_));
AND2X2 AND2X2_1896 ( .A(_abc_44694_new_n4181_), .B(_abc_44694_new_n4179_), .Y(_abc_44694_new_n4182_));
AND2X2 AND2X2_1897 ( .A(_abc_44694_new_n4184_), .B(_abc_44694_new_n668__bF_buf3), .Y(_abc_44694_new_n4185_));
AND2X2 AND2X2_1898 ( .A(_abc_44694_new_n4185_), .B(_abc_44694_new_n4183_), .Y(_abc_44694_new_n4186_));
AND2X2 AND2X2_1899 ( .A(state_q_3_bF_buf4_), .B(pc_q_9_), .Y(_abc_44694_new_n4187_));
AND2X2 AND2X2_19 ( .A(_abc_44694_new_n625_), .B(inst_r_1_), .Y(_abc_44694_new_n645_));
AND2X2 AND2X2_190 ( .A(_abc_44694_new_n963_), .B(_abc_44694_new_n673__bF_buf3), .Y(_abc_44694_new_n964_));
AND2X2 AND2X2_1900 ( .A(_abc_44694_new_n4064__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48711_9_), .Y(_abc_44694_new_n4188_));
AND2X2 AND2X2_1901 ( .A(_abc_44694_new_n4167_), .B(_abc_44694_new_n4179_), .Y(_abc_44694_new_n4191_));
AND2X2 AND2X2_1902 ( .A(_abc_44694_new_n4179_), .B(_abc_44694_new_n4165_), .Y(_abc_44694_new_n4194_));
AND2X2 AND2X2_1903 ( .A(_abc_44694_new_n4193_), .B(_abc_44694_new_n4196_), .Y(_abc_44694_new_n4197_));
AND2X2 AND2X2_1904 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_10_), .B(int32_r_10_), .Y(_abc_44694_new_n4199_));
AND2X2 AND2X2_1905 ( .A(_abc_44694_new_n4200_), .B(_abc_44694_new_n985_), .Y(_abc_44694_new_n4201_));
AND2X2 AND2X2_1906 ( .A(_abc_44694_new_n4198_), .B(_abc_44694_new_n4201_), .Y(_abc_44694_new_n4202_));
AND2X2 AND2X2_1907 ( .A(_abc_44694_new_n4204_), .B(_abc_44694_new_n668__bF_buf2), .Y(_abc_44694_new_n4205_));
AND2X2 AND2X2_1908 ( .A(_abc_44694_new_n4205_), .B(_abc_44694_new_n4203_), .Y(_abc_44694_new_n4206_));
AND2X2 AND2X2_1909 ( .A(state_q_3_bF_buf3_), .B(pc_q_10_), .Y(_abc_44694_new_n4207_));
AND2X2 AND2X2_191 ( .A(_abc_44694_new_n965_), .B(_abc_44694_new_n966_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_));
AND2X2 AND2X2_1910 ( .A(_abc_44694_new_n4064__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48711_10_), .Y(_abc_44694_new_n4208_));
AND2X2 AND2X2_1911 ( .A(_abc_44694_new_n4203_), .B(_abc_44694_new_n4200_), .Y(_abc_44694_new_n4211_));
AND2X2 AND2X2_1912 ( .A(_abc_44694_new_n635_), .B(opcode_q_21_), .Y(_abc_44694_new_n4212_));
AND2X2 AND2X2_1913 ( .A(_abc_44694_new_n636_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_44694_new_n4213_));
AND2X2 AND2X2_1914 ( .A(_abc_44694_new_n4214_), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_44694_new_n4215_));
AND2X2 AND2X2_1915 ( .A(_abc_44694_new_n4216_), .B(_abc_44694_new_n4217_), .Y(_abc_44694_new_n4218_));
AND2X2 AND2X2_1916 ( .A(_abc_44694_new_n4211_), .B(_abc_44694_new_n4218_), .Y(_abc_44694_new_n4219_));
AND2X2 AND2X2_1917 ( .A(_abc_44694_new_n4220_), .B(_abc_44694_new_n4221_), .Y(_abc_44694_new_n4222_));
AND2X2 AND2X2_1918 ( .A(_abc_44694_new_n4223_), .B(_abc_44694_new_n668__bF_buf1), .Y(_abc_44694_new_n4224_));
AND2X2 AND2X2_1919 ( .A(state_q_3_bF_buf2_), .B(pc_q_11_), .Y(_abc_44694_new_n4225_));
AND2X2 AND2X2_192 ( .A(_abc_44694_new_n626_), .B(_abc_44694_new_n639_), .Y(_abc_44694_new_n969_));
AND2X2 AND2X2_1920 ( .A(_abc_44694_new_n4064__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48711_11_), .Y(_abc_44694_new_n4226_));
AND2X2 AND2X2_1921 ( .A(_abc_44694_new_n635_), .B(opcode_q_22_), .Y(_abc_44694_new_n4229_));
AND2X2 AND2X2_1922 ( .A(_abc_44694_new_n636_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_44694_new_n4230_));
AND2X2 AND2X2_1923 ( .A(_abc_44694_new_n4231_), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_44694_new_n4232_));
AND2X2 AND2X2_1924 ( .A(_abc_44694_new_n4233_), .B(_abc_44694_new_n4234_), .Y(_abc_44694_new_n4235_));
AND2X2 AND2X2_1925 ( .A(_abc_44694_new_n4236_), .B(_abc_44694_new_n4217_), .Y(_abc_44694_new_n4237_));
AND2X2 AND2X2_1926 ( .A(_abc_44694_new_n4218_), .B(_abc_44694_new_n4201_), .Y(_abc_44694_new_n4238_));
AND2X2 AND2X2_1927 ( .A(_abc_44694_new_n4238_), .B(_abc_44694_new_n4195_), .Y(_abc_44694_new_n4239_));
AND2X2 AND2X2_1928 ( .A(_abc_44694_new_n4238_), .B(_abc_44694_new_n4191_), .Y(_abc_44694_new_n4241_));
AND2X2 AND2X2_1929 ( .A(_abc_44694_new_n4164_), .B(_abc_44694_new_n4241_), .Y(_abc_44694_new_n4242_));
AND2X2 AND2X2_193 ( .A(_abc_44694_new_n969_), .B(_abc_44694_new_n633_), .Y(_abc_44694_new_n970_));
AND2X2 AND2X2_1930 ( .A(_abc_44694_new_n4243_), .B(_abc_44694_new_n4235_), .Y(_abc_44694_new_n4245_));
AND2X2 AND2X2_1931 ( .A(_abc_44694_new_n4246_), .B(_abc_44694_new_n4244_), .Y(_abc_44694_new_n4247_));
AND2X2 AND2X2_1932 ( .A(_abc_44694_new_n4247_), .B(_abc_44694_new_n668__bF_buf0), .Y(_abc_44694_new_n4248_));
AND2X2 AND2X2_1933 ( .A(state_q_3_bF_buf1_), .B(pc_q_12_), .Y(_abc_44694_new_n4249_));
AND2X2 AND2X2_1934 ( .A(_abc_44694_new_n4064__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48711_12_), .Y(_abc_44694_new_n4250_));
AND2X2 AND2X2_1935 ( .A(_abc_44694_new_n635_), .B(opcode_q_23_), .Y(_abc_44694_new_n4253_));
AND2X2 AND2X2_1936 ( .A(_abc_44694_new_n636_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_44694_new_n4254_));
AND2X2 AND2X2_1937 ( .A(_abc_44694_new_n4255_), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_44694_new_n4256_));
AND2X2 AND2X2_1938 ( .A(_abc_44694_new_n4257_), .B(_abc_44694_new_n4258_), .Y(_abc_44694_new_n4259_));
AND2X2 AND2X2_1939 ( .A(_abc_44694_new_n4235_), .B(_abc_44694_new_n4259_), .Y(_abc_44694_new_n4262_));
AND2X2 AND2X2_194 ( .A(_abc_44694_new_n973_), .B(_abc_44694_new_n975_), .Y(_abc_44694_new_n976_));
AND2X2 AND2X2_1940 ( .A(_abc_44694_new_n4243_), .B(_abc_44694_new_n4262_), .Y(_abc_44694_new_n4263_));
AND2X2 AND2X2_1941 ( .A(_abc_44694_new_n4259_), .B(_abc_44694_new_n4232_), .Y(_abc_44694_new_n4265_));
AND2X2 AND2X2_1942 ( .A(_abc_44694_new_n4266_), .B(_abc_44694_new_n668__bF_buf4), .Y(_abc_44694_new_n4267_));
AND2X2 AND2X2_1943 ( .A(_abc_44694_new_n4264_), .B(_abc_44694_new_n4267_), .Y(_abc_44694_new_n4268_));
AND2X2 AND2X2_1944 ( .A(_abc_44694_new_n4268_), .B(_abc_44694_new_n4261_), .Y(_abc_44694_new_n4269_));
AND2X2 AND2X2_1945 ( .A(state_q_3_bF_buf0_), .B(pc_q_13_), .Y(_abc_44694_new_n4270_));
AND2X2 AND2X2_1946 ( .A(_abc_44694_new_n4064__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48711_13_), .Y(_abc_44694_new_n4271_));
AND2X2 AND2X2_1947 ( .A(_abc_44694_new_n4266_), .B(_abc_44694_new_n4257_), .Y(_abc_44694_new_n4274_));
AND2X2 AND2X2_1948 ( .A(_abc_44694_new_n4264_), .B(_abc_44694_new_n4274_), .Y(_abc_44694_new_n4275_));
AND2X2 AND2X2_1949 ( .A(_abc_44694_new_n635_), .B(opcode_q_24_), .Y(_abc_44694_new_n4277_));
AND2X2 AND2X2_195 ( .A(_abc_44694_new_n978_), .B(_abc_44694_new_n979_), .Y(_abc_44694_new_n980_));
AND2X2 AND2X2_1950 ( .A(_abc_44694_new_n636_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_44694_new_n4278_));
AND2X2 AND2X2_1951 ( .A(_abc_44694_new_n4279_), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_44694_new_n4280_));
AND2X2 AND2X2_1952 ( .A(_abc_44694_new_n4281_), .B(_abc_44694_new_n4282_), .Y(_abc_44694_new_n4283_));
AND2X2 AND2X2_1953 ( .A(_abc_44694_new_n4276_), .B(_abc_44694_new_n4283_), .Y(_abc_44694_new_n4285_));
AND2X2 AND2X2_1954 ( .A(_abc_44694_new_n4286_), .B(_abc_44694_new_n668__bF_buf3), .Y(_abc_44694_new_n4287_));
AND2X2 AND2X2_1955 ( .A(_abc_44694_new_n4287_), .B(_abc_44694_new_n4284_), .Y(_abc_44694_new_n4288_));
AND2X2 AND2X2_1956 ( .A(state_q_3_bF_buf5_), .B(pc_q_14_), .Y(_abc_44694_new_n4289_));
AND2X2 AND2X2_1957 ( .A(_abc_44694_new_n4064__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48711_14_), .Y(_abc_44694_new_n4290_));
AND2X2 AND2X2_1958 ( .A(_abc_44694_new_n4286_), .B(_abc_44694_new_n4281_), .Y(_abc_44694_new_n4293_));
AND2X2 AND2X2_1959 ( .A(_abc_44694_new_n635_), .B(opcode_q_25_), .Y(_abc_44694_new_n4295_));
AND2X2 AND2X2_196 ( .A(_abc_44694_new_n980_), .B(_abc_44694_new_n977_), .Y(_abc_44694_new_n981_));
AND2X2 AND2X2_1960 ( .A(_abc_44694_new_n636_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3_), .Y(_abc_44694_new_n4296_));
AND2X2 AND2X2_1961 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_44694_new_n4298_));
AND2X2 AND2X2_1962 ( .A(_abc_44694_new_n4300_), .B(_abc_44694_new_n979_), .Y(_abc_44694_new_n4301_));
AND2X2 AND2X2_1963 ( .A(_abc_44694_new_n4302_), .B(_abc_44694_new_n4299_), .Y(_abc_44694_new_n4303_));
AND2X2 AND2X2_1964 ( .A(_abc_44694_new_n4294_), .B(_abc_44694_new_n4304_), .Y(_abc_44694_new_n4305_));
AND2X2 AND2X2_1965 ( .A(_abc_44694_new_n4293_), .B(_abc_44694_new_n4303_), .Y(_abc_44694_new_n4306_));
AND2X2 AND2X2_1966 ( .A(_abc_44694_new_n4309_), .B(state_q_5_bF_buf0_), .Y(_abc_44694_new_n4310_));
AND2X2 AND2X2_1967 ( .A(_abc_44694_new_n4308_), .B(_abc_44694_new_n4310_), .Y(_abc_44694_new_n4311_));
AND2X2 AND2X2_1968 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_15_), .Y(_abc_44694_new_n4312_));
AND2X2 AND2X2_1969 ( .A(state_q_3_bF_buf4_), .B(pc_q_15_), .Y(_abc_44694_new_n4313_));
AND2X2 AND2X2_197 ( .A(_abc_44694_new_n982_), .B(_abc_44694_new_n983_), .Y(_abc_44694_new_n984_));
AND2X2 AND2X2_1970 ( .A(_abc_44694_new_n4297__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_44694_new_n4316_));
AND2X2 AND2X2_1971 ( .A(_abc_44694_new_n4317_), .B(_abc_44694_new_n4318_), .Y(_abc_44694_new_n4319_));
AND2X2 AND2X2_1972 ( .A(_abc_44694_new_n4302_), .B(_abc_44694_new_n4280_), .Y(_abc_44694_new_n4320_));
AND2X2 AND2X2_1973 ( .A(_abc_44694_new_n4274_), .B(_abc_44694_new_n4322_), .Y(_abc_44694_new_n4323_));
AND2X2 AND2X2_1974 ( .A(_abc_44694_new_n4303_), .B(_abc_44694_new_n4283_), .Y(_abc_44694_new_n4326_));
AND2X2 AND2X2_1975 ( .A(_abc_44694_new_n4325_), .B(_abc_44694_new_n4327_), .Y(_abc_44694_new_n4328_));
AND2X2 AND2X2_1976 ( .A(_abc_44694_new_n4328_), .B(_abc_44694_new_n4319_), .Y(_abc_44694_new_n4330_));
AND2X2 AND2X2_1977 ( .A(_abc_44694_new_n4331_), .B(_abc_44694_new_n4329_), .Y(_abc_44694_new_n4332_));
AND2X2 AND2X2_1978 ( .A(_abc_44694_new_n4332_), .B(_abc_44694_new_n668__bF_buf2), .Y(_abc_44694_new_n4333_));
AND2X2 AND2X2_1979 ( .A(state_q_3_bF_buf3_), .B(pc_q_16_), .Y(_abc_44694_new_n4334_));
AND2X2 AND2X2_198 ( .A(_abc_44694_new_n986_), .B(_abc_44694_new_n984_), .Y(_abc_44694_new_n987_));
AND2X2 AND2X2_1980 ( .A(_abc_44694_new_n4064__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48711_16_), .Y(_abc_44694_new_n4335_));
AND2X2 AND2X2_1981 ( .A(_abc_44694_new_n4331_), .B(_abc_44694_new_n4317_), .Y(_abc_44694_new_n4338_));
AND2X2 AND2X2_1982 ( .A(_abc_44694_new_n4297__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_44694_new_n4340_));
AND2X2 AND2X2_1983 ( .A(_abc_44694_new_n4341_), .B(_abc_44694_new_n4342_), .Y(_abc_44694_new_n4343_));
AND2X2 AND2X2_1984 ( .A(_abc_44694_new_n4339_), .B(_abc_44694_new_n4344_), .Y(_abc_44694_new_n4345_));
AND2X2 AND2X2_1985 ( .A(_abc_44694_new_n4338_), .B(_abc_44694_new_n4343_), .Y(_abc_44694_new_n4346_));
AND2X2 AND2X2_1986 ( .A(_abc_44694_new_n4349_), .B(state_q_5_bF_buf3_), .Y(_abc_44694_new_n4350_));
AND2X2 AND2X2_1987 ( .A(_abc_44694_new_n4348_), .B(_abc_44694_new_n4350_), .Y(_abc_44694_new_n4351_));
AND2X2 AND2X2_1988 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_17_), .Y(_abc_44694_new_n4352_));
AND2X2 AND2X2_1989 ( .A(state_q_3_bF_buf2_), .B(pc_q_17_), .Y(_abc_44694_new_n4353_));
AND2X2 AND2X2_199 ( .A(_abc_44694_new_n987_), .B(_abc_44694_new_n981_), .Y(_abc_44694_new_n988_));
AND2X2 AND2X2_1990 ( .A(_abc_44694_new_n4297__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_44694_new_n4356_));
AND2X2 AND2X2_1991 ( .A(_abc_44694_new_n4357_), .B(_abc_44694_new_n4358_), .Y(_abc_44694_new_n4359_));
AND2X2 AND2X2_1992 ( .A(_abc_44694_new_n4317_), .B(_abc_44694_new_n4341_), .Y(_abc_44694_new_n4360_));
AND2X2 AND2X2_1993 ( .A(_abc_44694_new_n4319_), .B(_abc_44694_new_n4343_), .Y(_abc_44694_new_n4362_));
AND2X2 AND2X2_1994 ( .A(_abc_44694_new_n4328_), .B(_abc_44694_new_n4362_), .Y(_abc_44694_new_n4363_));
AND2X2 AND2X2_1995 ( .A(_abc_44694_new_n4364_), .B(_abc_44694_new_n4359_), .Y(_abc_44694_new_n4366_));
AND2X2 AND2X2_1996 ( .A(_abc_44694_new_n4367_), .B(_abc_44694_new_n4365_), .Y(_abc_44694_new_n4368_));
AND2X2 AND2X2_1997 ( .A(_abc_44694_new_n4368_), .B(_abc_44694_new_n668__bF_buf1), .Y(_abc_44694_new_n4369_));
AND2X2 AND2X2_1998 ( .A(state_q_3_bF_buf1_), .B(pc_q_18_), .Y(_abc_44694_new_n4370_));
AND2X2 AND2X2_1999 ( .A(_abc_44694_new_n4064__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48711_18_), .Y(_abc_44694_new_n4371_));
AND2X2 AND2X2_2 ( .A(_abc_44694_new_n620_), .B(inst_r_3_), .Y(_abc_44694_new_n621_));
AND2X2 AND2X2_20 ( .A(_abc_44694_new_n624_), .B(inst_r_0_), .Y(_abc_44694_new_n647_));
AND2X2 AND2X2_200 ( .A(_abc_44694_new_n988_), .B(_abc_44694_new_n976_), .Y(_abc_44694_new_n989_));
AND2X2 AND2X2_2000 ( .A(_abc_44694_new_n4367_), .B(_abc_44694_new_n4357_), .Y(_abc_44694_new_n4374_));
AND2X2 AND2X2_2001 ( .A(_abc_44694_new_n4297__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_44694_new_n4376_));
AND2X2 AND2X2_2002 ( .A(_abc_44694_new_n4377_), .B(_abc_44694_new_n4378_), .Y(_abc_44694_new_n4379_));
AND2X2 AND2X2_2003 ( .A(_abc_44694_new_n4375_), .B(_abc_44694_new_n4380_), .Y(_abc_44694_new_n4381_));
AND2X2 AND2X2_2004 ( .A(_abc_44694_new_n4374_), .B(_abc_44694_new_n4379_), .Y(_abc_44694_new_n4382_));
AND2X2 AND2X2_2005 ( .A(_abc_44694_new_n4385_), .B(state_q_5_bF_buf2_), .Y(_abc_44694_new_n4386_));
AND2X2 AND2X2_2006 ( .A(_abc_44694_new_n4384_), .B(_abc_44694_new_n4386_), .Y(_abc_44694_new_n4387_));
AND2X2 AND2X2_2007 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_19_), .Y(_abc_44694_new_n4388_));
AND2X2 AND2X2_2008 ( .A(state_q_3_bF_buf0_), .B(pc_q_19_), .Y(_abc_44694_new_n4389_));
AND2X2 AND2X2_2009 ( .A(_abc_44694_new_n4359_), .B(_abc_44694_new_n4379_), .Y(_abc_44694_new_n4392_));
AND2X2 AND2X2_201 ( .A(_abc_44694_new_n991_), .B(_abc_44694_new_n992_), .Y(_abc_44694_new_n993_));
AND2X2 AND2X2_2010 ( .A(_abc_44694_new_n4362_), .B(_abc_44694_new_n4392_), .Y(_abc_44694_new_n4393_));
AND2X2 AND2X2_2011 ( .A(_abc_44694_new_n4328_), .B(_abc_44694_new_n4393_), .Y(_abc_44694_new_n4394_));
AND2X2 AND2X2_2012 ( .A(_abc_44694_new_n4392_), .B(_abc_44694_new_n4361_), .Y(_abc_44694_new_n4395_));
AND2X2 AND2X2_2013 ( .A(_abc_44694_new_n4357_), .B(_abc_44694_new_n4377_), .Y(_abc_44694_new_n4397_));
AND2X2 AND2X2_2014 ( .A(_abc_44694_new_n4396_), .B(_abc_44694_new_n4397_), .Y(_abc_44694_new_n4398_));
AND2X2 AND2X2_2015 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_44694_new_n4401_));
AND2X2 AND2X2_2016 ( .A(_abc_44694_new_n4402_), .B(_abc_44694_new_n4403_), .Y(_abc_44694_new_n4404_));
AND2X2 AND2X2_2017 ( .A(_abc_44694_new_n4400_), .B(_abc_44694_new_n4404_), .Y(_abc_44694_new_n4406_));
AND2X2 AND2X2_2018 ( .A(_abc_44694_new_n4407_), .B(_abc_44694_new_n668__bF_buf0), .Y(_abc_44694_new_n4408_));
AND2X2 AND2X2_2019 ( .A(_abc_44694_new_n4408_), .B(_abc_44694_new_n4405_), .Y(_abc_44694_new_n4409_));
AND2X2 AND2X2_202 ( .A(_abc_44694_new_n996_), .B(_abc_44694_new_n994_), .Y(_abc_44694_new_n997_));
AND2X2 AND2X2_2020 ( .A(state_q_3_bF_buf5_), .B(pc_q_20_), .Y(_abc_44694_new_n4410_));
AND2X2 AND2X2_2021 ( .A(_abc_44694_new_n4064__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48711_20_), .Y(_abc_44694_new_n4411_));
AND2X2 AND2X2_2022 ( .A(_abc_44694_new_n4407_), .B(_abc_44694_new_n4402_), .Y(_abc_44694_new_n4414_));
AND2X2 AND2X2_2023 ( .A(_abc_44694_new_n4297__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_44694_new_n4415_));
AND2X2 AND2X2_2024 ( .A(_abc_44694_new_n4416_), .B(_abc_44694_new_n4417_), .Y(_abc_44694_new_n4418_));
AND2X2 AND2X2_2025 ( .A(_abc_44694_new_n4422_), .B(_abc_44694_new_n668__bF_buf4), .Y(_abc_44694_new_n4423_));
AND2X2 AND2X2_2026 ( .A(_abc_44694_new_n4423_), .B(_abc_44694_new_n4420_), .Y(_abc_44694_new_n4424_));
AND2X2 AND2X2_2027 ( .A(state_q_3_bF_buf4_), .B(pc_q_21_), .Y(_abc_44694_new_n4425_));
AND2X2 AND2X2_2028 ( .A(_abc_44694_new_n4064__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48711_21_), .Y(_abc_44694_new_n4426_));
AND2X2 AND2X2_2029 ( .A(_abc_44694_new_n4297__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_44694_new_n4429_));
AND2X2 AND2X2_203 ( .A(_abc_44694_new_n993_), .B(_abc_44694_new_n997_), .Y(_abc_44694_new_n998_));
AND2X2 AND2X2_2030 ( .A(_abc_44694_new_n4430_), .B(_abc_44694_new_n4431_), .Y(_abc_44694_new_n4432_));
AND2X2 AND2X2_2031 ( .A(_abc_44694_new_n4402_), .B(_abc_44694_new_n4416_), .Y(_abc_44694_new_n4433_));
AND2X2 AND2X2_2032 ( .A(_abc_44694_new_n4404_), .B(_abc_44694_new_n4418_), .Y(_abc_44694_new_n4435_));
AND2X2 AND2X2_2033 ( .A(_abc_44694_new_n4400_), .B(_abc_44694_new_n4435_), .Y(_abc_44694_new_n4436_));
AND2X2 AND2X2_2034 ( .A(_abc_44694_new_n4437_), .B(_abc_44694_new_n4432_), .Y(_abc_44694_new_n4439_));
AND2X2 AND2X2_2035 ( .A(_abc_44694_new_n4440_), .B(_abc_44694_new_n4438_), .Y(_abc_44694_new_n4441_));
AND2X2 AND2X2_2036 ( .A(_abc_44694_new_n4441_), .B(_abc_44694_new_n668__bF_buf3), .Y(_abc_44694_new_n4442_));
AND2X2 AND2X2_2037 ( .A(state_q_3_bF_buf3_), .B(pc_q_22_), .Y(_abc_44694_new_n4443_));
AND2X2 AND2X2_2038 ( .A(_abc_44694_new_n4064__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48711_22_), .Y(_abc_44694_new_n4444_));
AND2X2 AND2X2_2039 ( .A(_abc_44694_new_n4440_), .B(_abc_44694_new_n4430_), .Y(_abc_44694_new_n4447_));
AND2X2 AND2X2_204 ( .A(_abc_44694_new_n1000_), .B(_abc_44694_new_n1002_), .Y(_abc_44694_new_n1003_));
AND2X2 AND2X2_2040 ( .A(_abc_44694_new_n4297__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_44694_new_n4449_));
AND2X2 AND2X2_2041 ( .A(_abc_44694_new_n4450_), .B(_abc_44694_new_n4451_), .Y(_abc_44694_new_n4452_));
AND2X2 AND2X2_2042 ( .A(_abc_44694_new_n4448_), .B(_abc_44694_new_n4453_), .Y(_abc_44694_new_n4454_));
AND2X2 AND2X2_2043 ( .A(_abc_44694_new_n4447_), .B(_abc_44694_new_n4452_), .Y(_abc_44694_new_n4455_));
AND2X2 AND2X2_2044 ( .A(_abc_44694_new_n4458_), .B(state_q_5_bF_buf1_), .Y(_abc_44694_new_n4459_));
AND2X2 AND2X2_2045 ( .A(_abc_44694_new_n4457_), .B(_abc_44694_new_n4459_), .Y(_abc_44694_new_n4460_));
AND2X2 AND2X2_2046 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_23_), .Y(_abc_44694_new_n4461_));
AND2X2 AND2X2_2047 ( .A(state_q_3_bF_buf2_), .B(pc_q_23_), .Y(_abc_44694_new_n4462_));
AND2X2 AND2X2_2048 ( .A(_abc_44694_new_n4432_), .B(_abc_44694_new_n4452_), .Y(_abc_44694_new_n4465_));
AND2X2 AND2X2_2049 ( .A(_abc_44694_new_n4465_), .B(_abc_44694_new_n4434_), .Y(_abc_44694_new_n4466_));
AND2X2 AND2X2_205 ( .A(_abc_44694_new_n1005_), .B(_abc_44694_new_n1007_), .Y(_abc_44694_new_n1008_));
AND2X2 AND2X2_2050 ( .A(_abc_44694_new_n4430_), .B(_abc_44694_new_n4450_), .Y(_abc_44694_new_n4468_));
AND2X2 AND2X2_2051 ( .A(_abc_44694_new_n4467_), .B(_abc_44694_new_n4468_), .Y(_abc_44694_new_n4469_));
AND2X2 AND2X2_2052 ( .A(_abc_44694_new_n4435_), .B(_abc_44694_new_n4465_), .Y(_abc_44694_new_n4470_));
AND2X2 AND2X2_2053 ( .A(_abc_44694_new_n4472_), .B(_abc_44694_new_n4469_), .Y(_abc_44694_new_n4473_));
AND2X2 AND2X2_2054 ( .A(_abc_44694_new_n4393_), .B(_abc_44694_new_n4470_), .Y(_abc_44694_new_n4475_));
AND2X2 AND2X2_2055 ( .A(_abc_44694_new_n4477_), .B(_abc_44694_new_n4473_), .Y(_abc_44694_new_n4478_));
AND2X2 AND2X2_2056 ( .A(_abc_44694_new_n4297__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_44694_new_n4480_));
AND2X2 AND2X2_2057 ( .A(_abc_44694_new_n4481_), .B(_abc_44694_new_n4482_), .Y(_abc_44694_new_n4483_));
AND2X2 AND2X2_2058 ( .A(_abc_44694_new_n4479_), .B(_abc_44694_new_n4483_), .Y(_abc_44694_new_n4485_));
AND2X2 AND2X2_2059 ( .A(_abc_44694_new_n4486_), .B(_abc_44694_new_n4484_), .Y(_abc_44694_new_n4487_));
AND2X2 AND2X2_206 ( .A(_abc_44694_new_n1003_), .B(_abc_44694_new_n1008_), .Y(_abc_44694_new_n1009_));
AND2X2 AND2X2_2060 ( .A(_abc_44694_new_n4487_), .B(_abc_44694_new_n668__bF_buf2), .Y(_abc_44694_new_n4488_));
AND2X2 AND2X2_2061 ( .A(state_q_3_bF_buf1_), .B(pc_q_24_), .Y(_abc_44694_new_n4489_));
AND2X2 AND2X2_2062 ( .A(_abc_44694_new_n4064__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48711_24_), .Y(_abc_44694_new_n4490_));
AND2X2 AND2X2_2063 ( .A(_abc_44694_new_n4486_), .B(_abc_44694_new_n4481_), .Y(_abc_44694_new_n4493_));
AND2X2 AND2X2_2064 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_44694_new_n4495_));
AND2X2 AND2X2_2065 ( .A(_abc_44694_new_n4496_), .B(_abc_44694_new_n4497_), .Y(_abc_44694_new_n4498_));
AND2X2 AND2X2_2066 ( .A(_abc_44694_new_n4494_), .B(_abc_44694_new_n4499_), .Y(_abc_44694_new_n4500_));
AND2X2 AND2X2_2067 ( .A(_abc_44694_new_n4493_), .B(_abc_44694_new_n4498_), .Y(_abc_44694_new_n4501_));
AND2X2 AND2X2_2068 ( .A(_abc_44694_new_n4504_), .B(state_q_5_bF_buf0_), .Y(_abc_44694_new_n4505_));
AND2X2 AND2X2_2069 ( .A(_abc_44694_new_n4503_), .B(_abc_44694_new_n4505_), .Y(_abc_44694_new_n4506_));
AND2X2 AND2X2_207 ( .A(_abc_44694_new_n1009_), .B(_abc_44694_new_n998_), .Y(_abc_44694_new_n1010_));
AND2X2 AND2X2_2070 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_25_), .Y(_abc_44694_new_n4507_));
AND2X2 AND2X2_2071 ( .A(state_q_3_bF_buf0_), .B(pc_q_25_), .Y(_abc_44694_new_n4508_));
AND2X2 AND2X2_2072 ( .A(_abc_44694_new_n4483_), .B(_abc_44694_new_n4498_), .Y(_abc_44694_new_n4511_));
AND2X2 AND2X2_2073 ( .A(_abc_44694_new_n4481_), .B(_abc_44694_new_n4496_), .Y(_abc_44694_new_n4514_));
AND2X2 AND2X2_2074 ( .A(_abc_44694_new_n4513_), .B(_abc_44694_new_n4514_), .Y(_abc_44694_new_n4515_));
AND2X2 AND2X2_2075 ( .A(_abc_44694_new_n4297__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_44694_new_n4517_));
AND2X2 AND2X2_2076 ( .A(_abc_44694_new_n4518_), .B(_abc_44694_new_n4519_), .Y(_abc_44694_new_n4520_));
AND2X2 AND2X2_2077 ( .A(_abc_44694_new_n4516_), .B(_abc_44694_new_n4520_), .Y(_abc_44694_new_n4522_));
AND2X2 AND2X2_2078 ( .A(_abc_44694_new_n4523_), .B(_abc_44694_new_n4521_), .Y(_abc_44694_new_n4524_));
AND2X2 AND2X2_2079 ( .A(_abc_44694_new_n4524_), .B(_abc_44694_new_n668__bF_buf1), .Y(_abc_44694_new_n4525_));
AND2X2 AND2X2_208 ( .A(_abc_44694_new_n1010_), .B(_abc_44694_new_n989_), .Y(_abc_44694_new_n1011_));
AND2X2 AND2X2_2080 ( .A(state_q_3_bF_buf5_), .B(pc_q_26_), .Y(_abc_44694_new_n4526_));
AND2X2 AND2X2_2081 ( .A(_abc_44694_new_n4064__bF_buf4), .B(_auto_iopadmap_cc_368_execute_48711_26_), .Y(_abc_44694_new_n4527_));
AND2X2 AND2X2_2082 ( .A(_abc_44694_new_n4523_), .B(_abc_44694_new_n4518_), .Y(_abc_44694_new_n4530_));
AND2X2 AND2X2_2083 ( .A(_abc_44694_new_n4297__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_44694_new_n4532_));
AND2X2 AND2X2_2084 ( .A(_abc_44694_new_n4533_), .B(_abc_44694_new_n4534_), .Y(_abc_44694_new_n4535_));
AND2X2 AND2X2_2085 ( .A(_abc_44694_new_n4538_), .B(_abc_44694_new_n668__bF_buf0), .Y(_abc_44694_new_n4539_));
AND2X2 AND2X2_2086 ( .A(_abc_44694_new_n4539_), .B(_abc_44694_new_n4536_), .Y(_abc_44694_new_n4540_));
AND2X2 AND2X2_2087 ( .A(state_q_3_bF_buf4_), .B(pc_q_27_), .Y(_abc_44694_new_n4541_));
AND2X2 AND2X2_2088 ( .A(_abc_44694_new_n4064__bF_buf3), .B(_auto_iopadmap_cc_368_execute_48711_27_), .Y(_abc_44694_new_n4542_));
AND2X2 AND2X2_2089 ( .A(_abc_44694_new_n4520_), .B(_abc_44694_new_n4535_), .Y(_abc_44694_new_n4545_));
AND2X2 AND2X2_209 ( .A(_abc_44694_new_n1011_), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n1013_));
AND2X2 AND2X2_2090 ( .A(_abc_44694_new_n4511_), .B(_abc_44694_new_n4545_), .Y(_abc_44694_new_n4546_));
AND2X2 AND2X2_2091 ( .A(_abc_44694_new_n4479_), .B(_abc_44694_new_n4546_), .Y(_abc_44694_new_n4547_));
AND2X2 AND2X2_2092 ( .A(_abc_44694_new_n4518_), .B(_abc_44694_new_n4533_), .Y(_abc_44694_new_n4551_));
AND2X2 AND2X2_2093 ( .A(_abc_44694_new_n4550_), .B(_abc_44694_new_n4551_), .Y(_abc_44694_new_n4552_));
AND2X2 AND2X2_2094 ( .A(_abc_44694_new_n4548_), .B(_abc_44694_new_n4552_), .Y(_abc_44694_new_n4553_));
AND2X2 AND2X2_2095 ( .A(_abc_44694_new_n4297__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_44694_new_n4555_));
AND2X2 AND2X2_2096 ( .A(_abc_44694_new_n4300_), .B(_abc_44694_new_n4556_), .Y(_abc_44694_new_n4557_));
AND2X2 AND2X2_2097 ( .A(_abc_44694_new_n4554_), .B(_abc_44694_new_n4559_), .Y(_abc_44694_new_n4561_));
AND2X2 AND2X2_2098 ( .A(_abc_44694_new_n4562_), .B(_abc_44694_new_n668__bF_buf4), .Y(_abc_44694_new_n4563_));
AND2X2 AND2X2_2099 ( .A(_abc_44694_new_n4563_), .B(_abc_44694_new_n4560_), .Y(_abc_44694_new_n4564_));
AND2X2 AND2X2_21 ( .A(_abc_44694_new_n646_), .B(_abc_44694_new_n648_), .Y(_abc_44694_new_n649_));
AND2X2 AND2X2_210 ( .A(_abc_44694_new_n1014_), .B(_abc_44694_new_n1012_), .Y(_abc_44694_new_n1015_));
AND2X2 AND2X2_2100 ( .A(state_q_3_bF_buf3_), .B(pc_q_28_), .Y(_abc_44694_new_n4565_));
AND2X2 AND2X2_2101 ( .A(_abc_44694_new_n4064__bF_buf2), .B(_auto_iopadmap_cc_368_execute_48711_28_), .Y(_abc_44694_new_n4566_));
AND2X2 AND2X2_2102 ( .A(_abc_44694_new_n4297__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_44694_new_n4571_));
AND2X2 AND2X2_2103 ( .A(_abc_44694_new_n4300_), .B(_abc_44694_new_n4572_), .Y(_abc_44694_new_n4573_));
AND2X2 AND2X2_2104 ( .A(_abc_44694_new_n4570_), .B(_abc_44694_new_n4575_), .Y(_abc_44694_new_n4576_));
AND2X2 AND2X2_2105 ( .A(_abc_44694_new_n4569_), .B(_abc_44694_new_n4574_), .Y(_abc_44694_new_n4577_));
AND2X2 AND2X2_2106 ( .A(_abc_44694_new_n4580_), .B(state_q_5_bF_buf3_), .Y(_abc_44694_new_n4581_));
AND2X2 AND2X2_2107 ( .A(_abc_44694_new_n4579_), .B(_abc_44694_new_n4581_), .Y(_abc_44694_new_n4582_));
AND2X2 AND2X2_2108 ( .A(_abc_44694_new_n4047_), .B(_auto_iopadmap_cc_368_execute_48711_29_), .Y(_abc_44694_new_n4583_));
AND2X2 AND2X2_2109 ( .A(state_q_3_bF_buf2_), .B(pc_q_29_), .Y(_abc_44694_new_n4584_));
AND2X2 AND2X2_211 ( .A(_abc_44694_new_n1015_), .B(_abc_44694_new_n970_), .Y(_abc_44694_new_n1016_));
AND2X2 AND2X2_2110 ( .A(_abc_44694_new_n4297__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_44694_new_n4587_));
AND2X2 AND2X2_2111 ( .A(_abc_44694_new_n4588_), .B(_abc_44694_new_n4589_), .Y(_abc_44694_new_n4590_));
AND2X2 AND2X2_2112 ( .A(_abc_44694_new_n4556_), .B(_abc_44694_new_n4572_), .Y(_abc_44694_new_n4591_));
AND2X2 AND2X2_2113 ( .A(_abc_44694_new_n4559_), .B(_abc_44694_new_n4575_), .Y(_abc_44694_new_n4593_));
AND2X2 AND2X2_2114 ( .A(_abc_44694_new_n4595_), .B(_abc_44694_new_n4592_), .Y(_abc_44694_new_n4596_));
AND2X2 AND2X2_2115 ( .A(_abc_44694_new_n4600_), .B(_abc_44694_new_n668__bF_buf3), .Y(_abc_44694_new_n4601_));
AND2X2 AND2X2_2116 ( .A(_abc_44694_new_n4601_), .B(_abc_44694_new_n4598_), .Y(_abc_44694_new_n4602_));
AND2X2 AND2X2_2117 ( .A(state_q_3_bF_buf1_), .B(pc_q_30_), .Y(_abc_44694_new_n4603_));
AND2X2 AND2X2_2118 ( .A(_abc_44694_new_n4064__bF_buf1), .B(_auto_iopadmap_cc_368_execute_48711_30_), .Y(_abc_44694_new_n4604_));
AND2X2 AND2X2_2119 ( .A(_abc_44694_new_n4600_), .B(_abc_44694_new_n4588_), .Y(_abc_44694_new_n4607_));
AND2X2 AND2X2_212 ( .A(_abc_44694_new_n621_), .B(_abc_44694_new_n647_), .Y(_abc_44694_new_n1018_));
AND2X2 AND2X2_2120 ( .A(_abc_44694_new_n4610_), .B(_abc_44694_new_n4611_), .Y(_abc_44694_new_n4612_));
AND2X2 AND2X2_2121 ( .A(_abc_44694_new_n4608_), .B(_abc_44694_new_n4613_), .Y(_abc_44694_new_n4614_));
AND2X2 AND2X2_2122 ( .A(_abc_44694_new_n4607_), .B(_abc_44694_new_n4612_), .Y(_abc_44694_new_n4615_));
AND2X2 AND2X2_2123 ( .A(_abc_44694_new_n4616_), .B(_abc_44694_new_n668__bF_buf2), .Y(_abc_44694_new_n4617_));
AND2X2 AND2X2_2124 ( .A(state_q_3_bF_buf0_), .B(pc_q_31_), .Y(_abc_44694_new_n4618_));
AND2X2 AND2X2_2125 ( .A(_abc_44694_new_n4064__bF_buf0), .B(_auto_iopadmap_cc_368_execute_48711_31_), .Y(_abc_44694_new_n4619_));
AND2X2 AND2X2_2126 ( .A(_abc_44694_new_n657_), .B(state_q_0_), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2386));
AND2X2 AND2X2_2127 ( .A(_abc_44694_new_n1044_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n4623_));
AND2X2 AND2X2_2128 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n4623_), .Y(_0nmi_q_0_0_));
AND2X2 AND2X2_2129 ( .A(_abc_44694_new_n1205_), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .Y(_abc_44694_new_n4625_));
AND2X2 AND2X2_213 ( .A(_abc_44694_new_n1018_), .B(_abc_44694_new_n619_), .Y(_abc_44694_new_n1019_));
AND2X2 AND2X2_2130 ( .A(_abc_44694_new_n4626_), .B(enable_i_bF_buf7), .Y(_0fault_o_0_0_));
AND2X2 AND2X2_2131 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2099_));
AND2X2 AND2X2_2132 ( .A(REGFILE_SIM_reg_bank_rd_i_0_), .B(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2100_));
AND2X2 AND2X2_2133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2099_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2100_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2101_));
AND2X2 AND2X2_2134 ( .A(REGFILE_SIM_reg_bank_rd_i_4_), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2102_));
AND2X2 AND2X2_2135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2101_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103_));
AND2X2 AND2X2_2136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2106_));
AND2X2 AND2X2_2137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2107_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2104_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__0_));
AND2X2 AND2X2_2138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2111_));
AND2X2 AND2X2_2139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2112_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2109_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__1_));
AND2X2 AND2X2_214 ( .A(_abc_44694_new_n1019__bF_buf4), .B(esr_q_2_), .Y(_abc_44694_new_n1020_));
AND2X2 AND2X2_2140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2116_));
AND2X2 AND2X2_2141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2117_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2114_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__2_));
AND2X2 AND2X2_2142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2121_));
AND2X2 AND2X2_2143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2122_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2119_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__3_));
AND2X2 AND2X2_2144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2126_));
AND2X2 AND2X2_2145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2127_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2124_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__4_));
AND2X2 AND2X2_2146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2131_));
AND2X2 AND2X2_2147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2132_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2129_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__5_));
AND2X2 AND2X2_2148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2136_));
AND2X2 AND2X2_2149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2137_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2134_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__6_));
AND2X2 AND2X2_215 ( .A(_abc_44694_new_n1021_), .B(sr_q_2_), .Y(_abc_44694_new_n1022_));
AND2X2 AND2X2_2150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2141_));
AND2X2 AND2X2_2151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2142_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2139_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__7_));
AND2X2 AND2X2_2152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2146_));
AND2X2 AND2X2_2153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2147_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2144_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__8_));
AND2X2 AND2X2_2154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2151_));
AND2X2 AND2X2_2155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2152_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2149_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__9_));
AND2X2 AND2X2_2156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2156_));
AND2X2 AND2X2_2157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2157_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2154_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__10_));
AND2X2 AND2X2_2158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2161_));
AND2X2 AND2X2_2159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2162_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2159_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__11_));
AND2X2 AND2X2_216 ( .A(_abc_44694_new_n1024_), .B(_abc_44694_new_n1017_), .Y(_abc_44694_new_n1025_));
AND2X2 AND2X2_2160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2166_));
AND2X2 AND2X2_2161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2167_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2164_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__12_));
AND2X2 AND2X2_2162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2171_));
AND2X2 AND2X2_2163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2172_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2169_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__13_));
AND2X2 AND2X2_2164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2176_));
AND2X2 AND2X2_2165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2177_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2174_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__14_));
AND2X2 AND2X2_2166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2181_));
AND2X2 AND2X2_2167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2182_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2179_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__15_));
AND2X2 AND2X2_2168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2186_));
AND2X2 AND2X2_2169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2187_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2184_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__16_));
AND2X2 AND2X2_217 ( .A(_abc_44694_new_n1027_), .B(intr_i), .Y(_abc_44694_new_n1028_));
AND2X2 AND2X2_2170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2191_));
AND2X2 AND2X2_2171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2192_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2189_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__17_));
AND2X2 AND2X2_2172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2196_));
AND2X2 AND2X2_2173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2197_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2194_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__18_));
AND2X2 AND2X2_2174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2201_));
AND2X2 AND2X2_2175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2202_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2199_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__19_));
AND2X2 AND2X2_2176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2206_));
AND2X2 AND2X2_2177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2207_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2204_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__20_));
AND2X2 AND2X2_2178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2211_));
AND2X2 AND2X2_2179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2212_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2209_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__21_));
AND2X2 AND2X2_218 ( .A(_abc_44694_new_n1029_), .B(_abc_44694_new_n996_), .Y(_abc_44694_new_n1030_));
AND2X2 AND2X2_2180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2216_));
AND2X2 AND2X2_2181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2217_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2214_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__22_));
AND2X2 AND2X2_2182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2221_));
AND2X2 AND2X2_2183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2222_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2219_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__23_));
AND2X2 AND2X2_2184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2226_));
AND2X2 AND2X2_2185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2224_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__24_));
AND2X2 AND2X2_2186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2231_));
AND2X2 AND2X2_2187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2232_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2229_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__25_));
AND2X2 AND2X2_2188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2236_));
AND2X2 AND2X2_2189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2237_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2234_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__26_));
AND2X2 AND2X2_219 ( .A(_abc_44694_new_n1008_), .B(_abc_44694_new_n1030_), .Y(_abc_44694_new_n1031_));
AND2X2 AND2X2_2190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2241_));
AND2X2 AND2X2_2191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2242_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2239_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__27_));
AND2X2 AND2X2_2192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2246_));
AND2X2 AND2X2_2193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2247_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2244_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__28_));
AND2X2 AND2X2_2194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2251_));
AND2X2 AND2X2_2195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2252_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2249_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__29_));
AND2X2 AND2X2_2196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2256_));
AND2X2 AND2X2_2197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2254_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__30_));
AND2X2 AND2X2_2198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2261_));
AND2X2 AND2X2_2199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2262_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2259_), .Y(REGFILE_SIM_reg_bank__0reg_r31_31_0__31_));
AND2X2 AND2X2_22 ( .A(_abc_44694_new_n637_), .B(_abc_44694_new_n631_), .Y(_abc_44694_new_n651_));
AND2X2 AND2X2_220 ( .A(_abc_44694_new_n991_), .B(_abc_44694_new_n1032_), .Y(_abc_44694_new_n1033_));
AND2X2 AND2X2_2200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2264_), .B(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2265_));
AND2X2 AND2X2_2201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2265_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2099_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2266_));
AND2X2 AND2X2_2202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2266_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2267_));
AND2X2 AND2X2_2203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2270_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2268_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__0_));
AND2X2 AND2X2_2204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2273_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2272_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__1_));
AND2X2 AND2X2_2205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2276_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2275_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__2_));
AND2X2 AND2X2_2206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2279_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2278_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__3_));
AND2X2 AND2X2_2207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2282_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2281_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__4_));
AND2X2 AND2X2_2208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2285_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2284_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__5_));
AND2X2 AND2X2_2209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2288_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2287_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__6_));
AND2X2 AND2X2_221 ( .A(_abc_44694_new_n1000_), .B(_abc_44694_new_n1001_), .Y(_abc_44694_new_n1034_));
AND2X2 AND2X2_2210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2291_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2290_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__7_));
AND2X2 AND2X2_2211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2294_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2293_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__8_));
AND2X2 AND2X2_2212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2297_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2296_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__9_));
AND2X2 AND2X2_2213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2300_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2299_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__10_));
AND2X2 AND2X2_2214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2303_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2302_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__11_));
AND2X2 AND2X2_2215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2306_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2305_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__12_));
AND2X2 AND2X2_2216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2309_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2308_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__13_));
AND2X2 AND2X2_2217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2312_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2311_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__14_));
AND2X2 AND2X2_2218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2315_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2314_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__15_));
AND2X2 AND2X2_2219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2318_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2317_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__16_));
AND2X2 AND2X2_222 ( .A(_abc_44694_new_n1033_), .B(_abc_44694_new_n1034_), .Y(_abc_44694_new_n1035_));
AND2X2 AND2X2_2220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2321_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2320_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__17_));
AND2X2 AND2X2_2221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2324_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2323_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__18_));
AND2X2 AND2X2_2222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2327_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2326_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__19_));
AND2X2 AND2X2_2223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2330_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2329_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__20_));
AND2X2 AND2X2_2224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2333_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2332_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__21_));
AND2X2 AND2X2_2225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2336_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2335_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__22_));
AND2X2 AND2X2_2226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2339_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2338_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__23_));
AND2X2 AND2X2_2227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2342_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2341_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__24_));
AND2X2 AND2X2_2228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2345_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2344_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__25_));
AND2X2 AND2X2_2229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2348_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2347_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__26_));
AND2X2 AND2X2_223 ( .A(_abc_44694_new_n1031_), .B(_abc_44694_new_n1035_), .Y(_abc_44694_new_n1036_));
AND2X2 AND2X2_2230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2351_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2350_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__27_));
AND2X2 AND2X2_2231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2354_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2353_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__28_));
AND2X2 AND2X2_2232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2357_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2356_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__29_));
AND2X2 AND2X2_2233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2360_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2359_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__30_));
AND2X2 AND2X2_2234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2363_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2362_), .Y(REGFILE_SIM_reg_bank__0reg_r30_31_0__31_));
AND2X2 AND2X2_2235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2365_), .B(REGFILE_SIM_reg_bank_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2366_));
AND2X2 AND2X2_2236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2366_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2099_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2367_));
AND2X2 AND2X2_2237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2368_));
AND2X2 AND2X2_2238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2371_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2369_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__0_));
AND2X2 AND2X2_2239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2374_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2373_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__1_));
AND2X2 AND2X2_224 ( .A(_abc_44694_new_n1036_), .B(_abc_44694_new_n989_), .Y(_abc_44694_new_n1037_));
AND2X2 AND2X2_2240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2377_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2376_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__2_));
AND2X2 AND2X2_2241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2380_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2379_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__3_));
AND2X2 AND2X2_2242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2383_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2382_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__4_));
AND2X2 AND2X2_2243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2386_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2385_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__5_));
AND2X2 AND2X2_2244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2389_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2388_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__6_));
AND2X2 AND2X2_2245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2392_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2391_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__7_));
AND2X2 AND2X2_2246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2395_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2394_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__8_));
AND2X2 AND2X2_2247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2398_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2397_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__9_));
AND2X2 AND2X2_2248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2401_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2400_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__10_));
AND2X2 AND2X2_2249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2404_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2403_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__11_));
AND2X2 AND2X2_225 ( .A(_abc_44694_new_n1037_), .B(_abc_44694_new_n970_), .Y(_abc_44694_new_n1038_));
AND2X2 AND2X2_2250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2407_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2406_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__12_));
AND2X2 AND2X2_2251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2410_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2409_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__13_));
AND2X2 AND2X2_2252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2413_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2412_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__14_));
AND2X2 AND2X2_2253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2416_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2415_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__15_));
AND2X2 AND2X2_2254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2419_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2418_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__16_));
AND2X2 AND2X2_2255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2422_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2421_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__17_));
AND2X2 AND2X2_2256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2425_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2424_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__18_));
AND2X2 AND2X2_2257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2428_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2427_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__19_));
AND2X2 AND2X2_2258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2431_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2430_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__20_));
AND2X2 AND2X2_2259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2434_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2433_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__21_));
AND2X2 AND2X2_226 ( .A(_abc_44694_new_n1039_), .B(esr_q_2_), .Y(_abc_44694_new_n1040_));
AND2X2 AND2X2_2260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2437_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2436_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__22_));
AND2X2 AND2X2_2261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2440_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2439_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__23_));
AND2X2 AND2X2_2262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2443_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2442_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__24_));
AND2X2 AND2X2_2263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2446_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2445_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__25_));
AND2X2 AND2X2_2264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2449_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2448_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__26_));
AND2X2 AND2X2_2265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2452_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2451_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__27_));
AND2X2 AND2X2_2266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2455_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2454_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__28_));
AND2X2 AND2X2_2267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2458_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2457_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__29_));
AND2X2 AND2X2_2268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2461_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2460_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__30_));
AND2X2 AND2X2_2269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2464_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2463_), .Y(REGFILE_SIM_reg_bank__0reg_r29_31_0__31_));
AND2X2 AND2X2_227 ( .A(_abc_44694_new_n1038_), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n1041_));
AND2X2 AND2X2_2270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2264_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2365_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2466_));
AND2X2 AND2X2_2271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2466_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2467_));
AND2X2 AND2X2_2272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2467_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2099_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468_));
AND2X2 AND2X2_2273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2470_));
AND2X2 AND2X2_2274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2469_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__0_));
AND2X2 AND2X2_2275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2474_));
AND2X2 AND2X2_2276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2475_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2473_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__1_));
AND2X2 AND2X2_2277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2478_));
AND2X2 AND2X2_2278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2479_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2477_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__2_));
AND2X2 AND2X2_2279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2482_));
AND2X2 AND2X2_228 ( .A(_abc_44694_new_n627_), .B(_abc_44694_new_n1046_), .Y(_abc_44694_new_n1047_));
AND2X2 AND2X2_2280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2483_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2481_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__3_));
AND2X2 AND2X2_2281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2486_));
AND2X2 AND2X2_2282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2487_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2485_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__4_));
AND2X2 AND2X2_2283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2490_));
AND2X2 AND2X2_2284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2491_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2489_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__5_));
AND2X2 AND2X2_2285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2494_));
AND2X2 AND2X2_2286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2493_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__6_));
AND2X2 AND2X2_2287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2498_));
AND2X2 AND2X2_2288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2499_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2497_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__7_));
AND2X2 AND2X2_2289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2502_));
AND2X2 AND2X2_229 ( .A(_abc_44694_new_n1047_), .B(_abc_44694_new_n622_), .Y(_abc_44694_new_n1048_));
AND2X2 AND2X2_2290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2503_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2501_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__8_));
AND2X2 AND2X2_2291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2506_));
AND2X2 AND2X2_2292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2507_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2505_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__9_));
AND2X2 AND2X2_2293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2510_));
AND2X2 AND2X2_2294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2511_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2509_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__10_));
AND2X2 AND2X2_2295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2514_));
AND2X2 AND2X2_2296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2513_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__11_));
AND2X2 AND2X2_2297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2518_));
AND2X2 AND2X2_2298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2519_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2517_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__12_));
AND2X2 AND2X2_2299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2522_));
AND2X2 AND2X2_23 ( .A(_abc_44694_new_n650_), .B(_abc_44694_new_n651_), .Y(_abc_44694_new_n652_));
AND2X2 AND2X2_230 ( .A(_abc_44694_new_n621_), .B(_abc_44694_new_n633_), .Y(_abc_44694_new_n1051_));
AND2X2 AND2X2_2300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2523_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2521_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__13_));
AND2X2 AND2X2_2301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2526_));
AND2X2 AND2X2_2302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2527_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2525_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__14_));
AND2X2 AND2X2_2303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2530_));
AND2X2 AND2X2_2304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2531_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2529_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__15_));
AND2X2 AND2X2_2305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2534_));
AND2X2 AND2X2_2306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2535_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2533_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__16_));
AND2X2 AND2X2_2307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2538_));
AND2X2 AND2X2_2308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2539_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2537_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__17_));
AND2X2 AND2X2_2309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2542_));
AND2X2 AND2X2_231 ( .A(_abc_44694_new_n1051_), .B(_abc_44694_new_n626_), .Y(_abc_44694_new_n1052_));
AND2X2 AND2X2_2310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2543_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2541_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__18_));
AND2X2 AND2X2_2311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2546_));
AND2X2 AND2X2_2312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2547_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2545_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__19_));
AND2X2 AND2X2_2313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2550_));
AND2X2 AND2X2_2314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2551_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2549_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__20_));
AND2X2 AND2X2_2315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2554_));
AND2X2 AND2X2_2316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2555_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2553_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__21_));
AND2X2 AND2X2_2317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2558_));
AND2X2 AND2X2_2318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2559_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2557_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__22_));
AND2X2 AND2X2_2319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2562_));
AND2X2 AND2X2_232 ( .A(_abc_44694_new_n1053_), .B(_abc_44694_new_n1054_), .Y(_abc_44694_new_n1055_));
AND2X2 AND2X2_2320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2561_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__23_));
AND2X2 AND2X2_2321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2566_));
AND2X2 AND2X2_2322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2567_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2565_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__24_));
AND2X2 AND2X2_2323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2570_));
AND2X2 AND2X2_2324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2571_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2569_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__25_));
AND2X2 AND2X2_2325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2574_));
AND2X2 AND2X2_2326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2575_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2573_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__26_));
AND2X2 AND2X2_2327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2578_));
AND2X2 AND2X2_2328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2579_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2577_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__27_));
AND2X2 AND2X2_2329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2582_));
AND2X2 AND2X2_233 ( .A(_abc_44694_new_n1056_), .B(_abc_44694_new_n1057_), .Y(_abc_44694_new_n1058_));
AND2X2 AND2X2_2330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2583_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2581_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__28_));
AND2X2 AND2X2_2331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2586_));
AND2X2 AND2X2_2332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2587_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2585_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__29_));
AND2X2 AND2X2_2333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2590_));
AND2X2 AND2X2_2334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2591_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2589_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__30_));
AND2X2 AND2X2_2335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2594_));
AND2X2 AND2X2_2336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2595_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2593_), .Y(REGFILE_SIM_reg_bank__0reg_r28_31_0__31_));
AND2X2 AND2X2_2337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2597_), .B(REGFILE_SIM_reg_bank_rd_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2598_));
AND2X2 AND2X2_2338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2598_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2100_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2599_));
AND2X2 AND2X2_2339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2599_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2600_));
AND2X2 AND2X2_234 ( .A(_abc_44694_new_n1059_), .B(_abc_44694_new_n1060_), .Y(_abc_44694_new_n1061_));
AND2X2 AND2X2_2340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2603_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2601_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__0_));
AND2X2 AND2X2_2341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2606_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2605_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__1_));
AND2X2 AND2X2_2342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2609_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2608_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__2_));
AND2X2 AND2X2_2343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2612_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2611_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__3_));
AND2X2 AND2X2_2344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2615_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2614_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__4_));
AND2X2 AND2X2_2345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2618_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2617_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__5_));
AND2X2 AND2X2_2346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2621_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2620_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__6_));
AND2X2 AND2X2_2347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2623_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__7_));
AND2X2 AND2X2_2348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2627_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2626_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__8_));
AND2X2 AND2X2_2349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2630_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2629_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__9_));
AND2X2 AND2X2_235 ( .A(_abc_44694_new_n1058_), .B(_abc_44694_new_n1061_), .Y(_abc_44694_new_n1062_));
AND2X2 AND2X2_2350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2633_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2632_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__10_));
AND2X2 AND2X2_2351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2636_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2635_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__11_));
AND2X2 AND2X2_2352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2639_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2638_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__12_));
AND2X2 AND2X2_2353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2642_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2641_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__13_));
AND2X2 AND2X2_2354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2645_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2644_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__14_));
AND2X2 AND2X2_2355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2648_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2647_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__15_));
AND2X2 AND2X2_2356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2651_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2650_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__16_));
AND2X2 AND2X2_2357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2654_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2653_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__17_));
AND2X2 AND2X2_2358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2657_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2656_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__18_));
AND2X2 AND2X2_2359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2660_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2659_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__19_));
AND2X2 AND2X2_236 ( .A(_abc_44694_new_n1063_), .B(_abc_44694_new_n1064_), .Y(_abc_44694_new_n1065_));
AND2X2 AND2X2_2360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2663_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2662_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__20_));
AND2X2 AND2X2_2361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2666_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2665_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__21_));
AND2X2 AND2X2_2362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2669_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2668_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__22_));
AND2X2 AND2X2_2363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2672_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2671_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__23_));
AND2X2 AND2X2_2364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2675_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2674_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__24_));
AND2X2 AND2X2_2365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2678_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2677_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__25_));
AND2X2 AND2X2_2366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2681_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2680_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__26_));
AND2X2 AND2X2_2367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2684_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2683_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__27_));
AND2X2 AND2X2_2368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2687_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2686_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__28_));
AND2X2 AND2X2_2369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2690_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2689_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__29_));
AND2X2 AND2X2_237 ( .A(_abc_44694_new_n1062_), .B(_abc_44694_new_n1065_), .Y(_abc_44694_new_n1066_));
AND2X2 AND2X2_2370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2693_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2692_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__30_));
AND2X2 AND2X2_2371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2696_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2695_), .Y(REGFILE_SIM_reg_bank__0reg_r27_31_0__31_));
AND2X2 AND2X2_2372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2265_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2698_));
AND2X2 AND2X2_2373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2698_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699_));
AND2X2 AND2X2_2374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2701_));
AND2X2 AND2X2_2375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2702_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2700_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__0_));
AND2X2 AND2X2_2376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2705_));
AND2X2 AND2X2_2377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2706_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2704_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__1_));
AND2X2 AND2X2_2378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2709_));
AND2X2 AND2X2_2379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2710_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2708_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__2_));
AND2X2 AND2X2_238 ( .A(_abc_44694_new_n1066_), .B(_abc_44694_new_n1055_), .Y(_abc_44694_new_n1067_));
AND2X2 AND2X2_2380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2713_));
AND2X2 AND2X2_2381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2714_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2712_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__3_));
AND2X2 AND2X2_2382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2717_));
AND2X2 AND2X2_2383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2718_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2716_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__4_));
AND2X2 AND2X2_2384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2721_));
AND2X2 AND2X2_2385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2722_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2720_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__5_));
AND2X2 AND2X2_2386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2725_));
AND2X2 AND2X2_2387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2726_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2724_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__6_));
AND2X2 AND2X2_2388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2729_));
AND2X2 AND2X2_2389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2730_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2728_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__7_));
AND2X2 AND2X2_239 ( .A(_abc_44694_new_n1064_), .B(alu_op_r_0_), .Y(_abc_44694_new_n1068_));
AND2X2 AND2X2_2390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2733_));
AND2X2 AND2X2_2391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2734_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2732_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__8_));
AND2X2 AND2X2_2392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2737_));
AND2X2 AND2X2_2393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2738_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2736_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__9_));
AND2X2 AND2X2_2394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2741_));
AND2X2 AND2X2_2395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2742_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2740_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__10_));
AND2X2 AND2X2_2396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2745_));
AND2X2 AND2X2_2397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2746_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2744_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__11_));
AND2X2 AND2X2_2398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2749_));
AND2X2 AND2X2_2399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2750_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2748_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__12_));
AND2X2 AND2X2_24 ( .A(_abc_44694_new_n654_), .B(_abc_44694_new_n636_), .Y(_abc_44694_new_n655_));
AND2X2 AND2X2_240 ( .A(_abc_44694_new_n1062_), .B(_abc_44694_new_n1055_), .Y(_abc_44694_new_n1069_));
AND2X2 AND2X2_2400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2753_));
AND2X2 AND2X2_2401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2754_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2752_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__13_));
AND2X2 AND2X2_2402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2757_));
AND2X2 AND2X2_2403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2758_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2756_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__14_));
AND2X2 AND2X2_2404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2761_));
AND2X2 AND2X2_2405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2762_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2760_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__15_));
AND2X2 AND2X2_2406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2765_));
AND2X2 AND2X2_2407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2766_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2764_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__16_));
AND2X2 AND2X2_2408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2769_));
AND2X2 AND2X2_2409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2770_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2768_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__17_));
AND2X2 AND2X2_241 ( .A(_abc_44694_new_n1069_), .B(_abc_44694_new_n1068_), .Y(_abc_44694_new_n1070_));
AND2X2 AND2X2_2410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2773_));
AND2X2 AND2X2_2411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2774_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2772_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__18_));
AND2X2 AND2X2_2412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2777_));
AND2X2 AND2X2_2413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2778_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2776_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__19_));
AND2X2 AND2X2_2414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2781_));
AND2X2 AND2X2_2415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2782_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2780_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__20_));
AND2X2 AND2X2_2416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2785_));
AND2X2 AND2X2_2417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2786_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2784_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__21_));
AND2X2 AND2X2_2418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2789_));
AND2X2 AND2X2_2419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2790_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2788_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__22_));
AND2X2 AND2X2_242 ( .A(_abc_44694_new_n1071_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n1072_));
AND2X2 AND2X2_2420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2793_));
AND2X2 AND2X2_2421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2794_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2792_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__23_));
AND2X2 AND2X2_2422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2797_));
AND2X2 AND2X2_2423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2798_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2796_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__24_));
AND2X2 AND2X2_2424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2801_));
AND2X2 AND2X2_2425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2802_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2800_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__25_));
AND2X2 AND2X2_2426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2805_));
AND2X2 AND2X2_2427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2806_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2804_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__26_));
AND2X2 AND2X2_2428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2809_));
AND2X2 AND2X2_2429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2810_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2808_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__27_));
AND2X2 AND2X2_243 ( .A(_abc_44694_new_n1054_), .B(alu_op_r_2_), .Y(_abc_44694_new_n1073_));
AND2X2 AND2X2_2430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2813_));
AND2X2 AND2X2_2431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2814_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2812_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__28_));
AND2X2 AND2X2_2432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2817_));
AND2X2 AND2X2_2433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2818_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2816_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__29_));
AND2X2 AND2X2_2434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2821_));
AND2X2 AND2X2_2435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2822_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2820_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__30_));
AND2X2 AND2X2_2436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2825_));
AND2X2 AND2X2_2437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2826_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2824_), .Y(REGFILE_SIM_reg_bank__0reg_r26_31_0__31_));
AND2X2 AND2X2_2438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2366_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2828_));
AND2X2 AND2X2_2439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2828_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829_));
AND2X2 AND2X2_244 ( .A(_abc_44694_new_n1066_), .B(_abc_44694_new_n1073_), .Y(_abc_44694_new_n1074_));
AND2X2 AND2X2_2440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2831_));
AND2X2 AND2X2_2441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2832_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2830_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__0_));
AND2X2 AND2X2_2442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2835_));
AND2X2 AND2X2_2443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2836_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2834_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__1_));
AND2X2 AND2X2_2444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2839_));
AND2X2 AND2X2_2445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2840_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2838_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__2_));
AND2X2 AND2X2_2446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2843_));
AND2X2 AND2X2_2447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2844_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2842_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__3_));
AND2X2 AND2X2_2448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2847_));
AND2X2 AND2X2_2449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2848_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2846_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__4_));
AND2X2 AND2X2_245 ( .A(_abc_44694_new_n1074_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n1075_));
AND2X2 AND2X2_2450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2851_));
AND2X2 AND2X2_2451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2852_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2850_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__5_));
AND2X2 AND2X2_2452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2855_));
AND2X2 AND2X2_2453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2856_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2854_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__6_));
AND2X2 AND2X2_2454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2859_));
AND2X2 AND2X2_2455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2860_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2858_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__7_));
AND2X2 AND2X2_2456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2863_));
AND2X2 AND2X2_2457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2864_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2862_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__8_));
AND2X2 AND2X2_2458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2867_));
AND2X2 AND2X2_2459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2868_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2866_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__9_));
AND2X2 AND2X2_246 ( .A(alu_op_r_0_), .B(alu_op_r_1_), .Y(_abc_44694_new_n1076_));
AND2X2 AND2X2_2460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2871_));
AND2X2 AND2X2_2461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2872_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2870_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__10_));
AND2X2 AND2X2_2462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2875_));
AND2X2 AND2X2_2463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2876_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2874_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__11_));
AND2X2 AND2X2_2464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2879_));
AND2X2 AND2X2_2465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2880_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2878_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__12_));
AND2X2 AND2X2_2466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2883_));
AND2X2 AND2X2_2467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2884_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2882_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__13_));
AND2X2 AND2X2_2468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2887_));
AND2X2 AND2X2_2469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2888_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2886_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__14_));
AND2X2 AND2X2_247 ( .A(_abc_44694_new_n1052_), .B(_abc_44694_new_n1076_), .Y(_abc_44694_new_n1077_));
AND2X2 AND2X2_2470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2891_));
AND2X2 AND2X2_2471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2892_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2890_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__15_));
AND2X2 AND2X2_2472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2895_));
AND2X2 AND2X2_2473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2896_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2894_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__16_));
AND2X2 AND2X2_2474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2899_));
AND2X2 AND2X2_2475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2900_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2898_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__17_));
AND2X2 AND2X2_2476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2903_));
AND2X2 AND2X2_2477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2904_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2902_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__18_));
AND2X2 AND2X2_2478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2907_));
AND2X2 AND2X2_2479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2908_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2906_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__19_));
AND2X2 AND2X2_248 ( .A(_abc_44694_new_n1077_), .B(_abc_44694_new_n1069_), .Y(_abc_44694_new_n1078_));
AND2X2 AND2X2_2480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2911_));
AND2X2 AND2X2_2481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2912_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2910_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__20_));
AND2X2 AND2X2_2482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2915_));
AND2X2 AND2X2_2483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2916_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2914_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__21_));
AND2X2 AND2X2_2484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2919_));
AND2X2 AND2X2_2485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2920_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2918_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__22_));
AND2X2 AND2X2_2486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2923_));
AND2X2 AND2X2_2487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2924_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2922_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__23_));
AND2X2 AND2X2_2488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2927_));
AND2X2 AND2X2_2489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2928_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2926_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__24_));
AND2X2 AND2X2_249 ( .A(inst_r_2_), .B(inst_r_3_), .Y(_abc_44694_new_n1082_));
AND2X2 AND2X2_2490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2931_));
AND2X2 AND2X2_2491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2932_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2930_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__25_));
AND2X2 AND2X2_2492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2935_));
AND2X2 AND2X2_2493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2936_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2934_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__26_));
AND2X2 AND2X2_2494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2939_));
AND2X2 AND2X2_2495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2940_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2938_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__27_));
AND2X2 AND2X2_2496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2943_));
AND2X2 AND2X2_2497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2944_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2942_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__28_));
AND2X2 AND2X2_2498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2947_));
AND2X2 AND2X2_2499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2948_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2946_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__29_));
AND2X2 AND2X2_25 ( .A(_abc_44694_new_n655_), .B(state_q_5_bF_buf3_), .Y(_abc_44694_new_n656_));
AND2X2 AND2X2_250 ( .A(_abc_44694_new_n637_), .B(_abc_44694_new_n1082_), .Y(_abc_44694_new_n1083_));
AND2X2 AND2X2_2500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2951_));
AND2X2 AND2X2_2501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2952_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2950_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__30_));
AND2X2 AND2X2_2502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2955_));
AND2X2 AND2X2_2503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2956_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2954_), .Y(REGFILE_SIM_reg_bank__0reg_r25_31_0__31_));
AND2X2 AND2X2_2504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2467_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2958_));
AND2X2 AND2X2_2505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2961_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2959_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__0_));
AND2X2 AND2X2_2506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2964_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2963_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__1_));
AND2X2 AND2X2_2507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2967_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2966_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__2_));
AND2X2 AND2X2_2508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2970_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2969_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__3_));
AND2X2 AND2X2_2509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2973_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2972_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__4_));
AND2X2 AND2X2_251 ( .A(_abc_44694_new_n1083_), .B(_abc_44694_new_n638_), .Y(_abc_44694_new_n1084_));
AND2X2 AND2X2_2510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2976_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2975_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__5_));
AND2X2 AND2X2_2511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2979_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2978_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__6_));
AND2X2 AND2X2_2512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2982_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2981_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__7_));
AND2X2 AND2X2_2513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2985_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2984_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__8_));
AND2X2 AND2X2_2514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2988_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2987_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__9_));
AND2X2 AND2X2_2515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2991_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2990_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__10_));
AND2X2 AND2X2_2516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2994_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2993_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__11_));
AND2X2 AND2X2_2517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2997_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2996_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__12_));
AND2X2 AND2X2_2518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3000_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2999_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__13_));
AND2X2 AND2X2_2519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3003_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3002_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__14_));
AND2X2 AND2X2_252 ( .A(_abc_44694_new_n1051_), .B(_abc_44694_new_n647_), .Y(_abc_44694_new_n1086_));
AND2X2 AND2X2_2520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3006_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3005_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__15_));
AND2X2 AND2X2_2521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3009_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3008_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__16_));
AND2X2 AND2X2_2522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3012_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3011_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__17_));
AND2X2 AND2X2_2523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3015_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3014_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__18_));
AND2X2 AND2X2_2524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3018_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3017_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__19_));
AND2X2 AND2X2_2525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3021_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3020_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__20_));
AND2X2 AND2X2_2526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3024_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3023_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__21_));
AND2X2 AND2X2_2527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3027_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3026_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__22_));
AND2X2 AND2X2_2528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3030_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3029_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__23_));
AND2X2 AND2X2_2529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3033_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3032_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__24_));
AND2X2 AND2X2_253 ( .A(_abc_44694_new_n1085_), .B(_abc_44694_new_n1087__bF_buf3), .Y(_abc_44694_new_n1088_));
AND2X2 AND2X2_2530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3036_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3035_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__25_));
AND2X2 AND2X2_2531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3039_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3038_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__26_));
AND2X2 AND2X2_2532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3042_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3041_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__27_));
AND2X2 AND2X2_2533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3045_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3044_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__28_));
AND2X2 AND2X2_2534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3048_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3047_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__29_));
AND2X2 AND2X2_2535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3051_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3050_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__30_));
AND2X2 AND2X2_2536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3053_), .Y(REGFILE_SIM_reg_bank__0reg_r24_31_0__31_));
AND2X2 AND2X2_2537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3056_), .B(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3057_));
AND2X2 AND2X2_2538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3057_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2100_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3058_));
AND2X2 AND2X2_2539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3058_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3059_));
AND2X2 AND2X2_254 ( .A(_abc_44694_new_n1046_), .B(opcode_q_23_), .Y(_abc_44694_new_n1090_));
AND2X2 AND2X2_2540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3062_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3060_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__0_));
AND2X2 AND2X2_2541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3065_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3064_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__1_));
AND2X2 AND2X2_2542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3068_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3067_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__2_));
AND2X2 AND2X2_2543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3071_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3070_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__3_));
AND2X2 AND2X2_2544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3074_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3073_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__4_));
AND2X2 AND2X2_2545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3077_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3076_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__5_));
AND2X2 AND2X2_2546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3080_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3079_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__6_));
AND2X2 AND2X2_2547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3083_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3082_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__7_));
AND2X2 AND2X2_2548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3086_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3085_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__8_));
AND2X2 AND2X2_2549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3089_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3088_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__9_));
AND2X2 AND2X2_255 ( .A(inst_r_0_), .B(inst_r_3_), .Y(_abc_44694_new_n1091_));
AND2X2 AND2X2_2550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3092_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3091_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__10_));
AND2X2 AND2X2_2551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3095_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3094_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__11_));
AND2X2 AND2X2_2552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3098_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3097_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__12_));
AND2X2 AND2X2_2553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3101_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3100_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__13_));
AND2X2 AND2X2_2554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3104_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3103_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__14_));
AND2X2 AND2X2_2555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3107_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3106_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__15_));
AND2X2 AND2X2_2556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3110_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3109_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__16_));
AND2X2 AND2X2_2557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3113_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3112_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__17_));
AND2X2 AND2X2_2558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3116_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3115_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__18_));
AND2X2 AND2X2_2559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3119_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3118_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__19_));
AND2X2 AND2X2_256 ( .A(_abc_44694_new_n623_), .B(inst_r_5_), .Y(_abc_44694_new_n1092_));
AND2X2 AND2X2_2560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3122_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3121_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__20_));
AND2X2 AND2X2_2561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3125_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3124_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__21_));
AND2X2 AND2X2_2562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3128_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3127_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__22_));
AND2X2 AND2X2_2563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3131_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3130_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__23_));
AND2X2 AND2X2_2564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3134_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3133_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__24_));
AND2X2 AND2X2_2565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3137_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3136_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__25_));
AND2X2 AND2X2_2566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3140_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3139_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__26_));
AND2X2 AND2X2_2567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3143_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3142_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__27_));
AND2X2 AND2X2_2568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3146_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3145_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__28_));
AND2X2 AND2X2_2569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3149_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3148_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__29_));
AND2X2 AND2X2_257 ( .A(_abc_44694_new_n1092_), .B(_abc_44694_new_n1091_), .Y(_abc_44694_new_n1093_));
AND2X2 AND2X2_2570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3152_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3151_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__30_));
AND2X2 AND2X2_2571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3155_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3154_), .Y(REGFILE_SIM_reg_bank__0reg_r23_31_0__31_));
AND2X2 AND2X2_2572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2265_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3157_));
AND2X2 AND2X2_2573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3157_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158_));
AND2X2 AND2X2_2574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3160_));
AND2X2 AND2X2_2575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3161_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3159_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__0_));
AND2X2 AND2X2_2576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3164_));
AND2X2 AND2X2_2577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3165_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3163_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__1_));
AND2X2 AND2X2_2578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3168_));
AND2X2 AND2X2_2579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3169_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3167_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__2_));
AND2X2 AND2X2_258 ( .A(_abc_44694_new_n1094_), .B(_abc_44694_new_n1095_), .Y(_abc_44694_new_n1096_));
AND2X2 AND2X2_2580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3172_));
AND2X2 AND2X2_2581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3173_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3171_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__3_));
AND2X2 AND2X2_2582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3176_));
AND2X2 AND2X2_2583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3177_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3175_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__4_));
AND2X2 AND2X2_2584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3180_));
AND2X2 AND2X2_2585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3181_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3179_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__5_));
AND2X2 AND2X2_2586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3184_));
AND2X2 AND2X2_2587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3185_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3183_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__6_));
AND2X2 AND2X2_2588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3188_));
AND2X2 AND2X2_2589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3189_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3187_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__7_));
AND2X2 AND2X2_259 ( .A(_abc_44694_new_n1093_), .B(_abc_44694_new_n1096_), .Y(_abc_44694_new_n1097_));
AND2X2 AND2X2_2590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3192_));
AND2X2 AND2X2_2591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3193_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3191_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__8_));
AND2X2 AND2X2_2592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3196_));
AND2X2 AND2X2_2593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3197_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3195_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__9_));
AND2X2 AND2X2_2594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3200_));
AND2X2 AND2X2_2595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3201_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3199_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__10_));
AND2X2 AND2X2_2596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3204_));
AND2X2 AND2X2_2597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3205_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3203_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__11_));
AND2X2 AND2X2_2598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3208_));
AND2X2 AND2X2_2599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3209_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3207_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__12_));
AND2X2 AND2X2_26 ( .A(_abc_44694_new_n657_), .B(state_q_4_), .Y(_abc_44694_new_n658_));
AND2X2 AND2X2_260 ( .A(_abc_44694_new_n1097_), .B(_abc_44694_new_n1090_), .Y(_abc_44694_new_n1098_));
AND2X2 AND2X2_2600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3212_));
AND2X2 AND2X2_2601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3213_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3211_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__13_));
AND2X2 AND2X2_2602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3216_));
AND2X2 AND2X2_2603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3217_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3215_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__14_));
AND2X2 AND2X2_2604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3220_));
AND2X2 AND2X2_2605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3221_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3219_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__15_));
AND2X2 AND2X2_2606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3224_));
AND2X2 AND2X2_2607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3225_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3223_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__16_));
AND2X2 AND2X2_2608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3228_));
AND2X2 AND2X2_2609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3229_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3227_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__17_));
AND2X2 AND2X2_261 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1098_), .Y(_abc_44694_new_n1099_));
AND2X2 AND2X2_2610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3232_));
AND2X2 AND2X2_2611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3233_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3231_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__18_));
AND2X2 AND2X2_2612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3236_));
AND2X2 AND2X2_2613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3237_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3235_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__19_));
AND2X2 AND2X2_2614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3240_));
AND2X2 AND2X2_2615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3241_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3239_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__20_));
AND2X2 AND2X2_2616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3244_));
AND2X2 AND2X2_2617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3245_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3243_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__21_));
AND2X2 AND2X2_2618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3248_));
AND2X2 AND2X2_2619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3249_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3247_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__22_));
AND2X2 AND2X2_262 ( .A(_abc_44694_new_n1053_), .B(alu_op_r_3_), .Y(_abc_44694_new_n1100_));
AND2X2 AND2X2_2620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3252_));
AND2X2 AND2X2_2621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3253_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3251_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__23_));
AND2X2 AND2X2_2622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3256_));
AND2X2 AND2X2_2623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3255_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__24_));
AND2X2 AND2X2_2624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3260_));
AND2X2 AND2X2_2625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3261_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3259_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__25_));
AND2X2 AND2X2_2626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3264_));
AND2X2 AND2X2_2627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3265_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3263_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__26_));
AND2X2 AND2X2_2628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3268_));
AND2X2 AND2X2_2629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3269_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3267_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__27_));
AND2X2 AND2X2_263 ( .A(_abc_44694_new_n1065_), .B(_abc_44694_new_n1100_), .Y(_abc_44694_new_n1101_));
AND2X2 AND2X2_2630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3272_));
AND2X2 AND2X2_2631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3273_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3271_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__28_));
AND2X2 AND2X2_2632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3276_));
AND2X2 AND2X2_2633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3277_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3275_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__29_));
AND2X2 AND2X2_2634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3280_));
AND2X2 AND2X2_2635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3281_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3279_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__30_));
AND2X2 AND2X2_2636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3284_));
AND2X2 AND2X2_2637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3285_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3283_), .Y(REGFILE_SIM_reg_bank__0reg_r22_31_0__31_));
AND2X2 AND2X2_2638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2366_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3287_));
AND2X2 AND2X2_2639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3287_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288_));
AND2X2 AND2X2_264 ( .A(_abc_44694_new_n1052_), .B(_abc_44694_new_n1101_), .Y(_abc_44694_new_n1102_));
AND2X2 AND2X2_2640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3290_));
AND2X2 AND2X2_2641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3291_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3289_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__0_));
AND2X2 AND2X2_2642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3294_));
AND2X2 AND2X2_2643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3295_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3293_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__1_));
AND2X2 AND2X2_2644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3298_));
AND2X2 AND2X2_2645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3299_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3297_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__2_));
AND2X2 AND2X2_2646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3302_));
AND2X2 AND2X2_2647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3303_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3301_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__3_));
AND2X2 AND2X2_2648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3306_));
AND2X2 AND2X2_2649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3307_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3305_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__4_));
AND2X2 AND2X2_265 ( .A(_abc_44694_new_n1061_), .B(_abc_44694_new_n1056_), .Y(_abc_44694_new_n1103_));
AND2X2 AND2X2_2650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3310_));
AND2X2 AND2X2_2651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3311_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3309_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__5_));
AND2X2 AND2X2_2652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3314_));
AND2X2 AND2X2_2653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3315_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3313_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__6_));
AND2X2 AND2X2_2654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3318_));
AND2X2 AND2X2_2655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3319_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3317_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__7_));
AND2X2 AND2X2_2656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3322_));
AND2X2 AND2X2_2657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3323_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3321_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__8_));
AND2X2 AND2X2_2658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3326_));
AND2X2 AND2X2_2659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3327_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3325_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__9_));
AND2X2 AND2X2_266 ( .A(_abc_44694_new_n1102_), .B(_abc_44694_new_n1103_), .Y(_abc_44694_new_n1104_));
AND2X2 AND2X2_2660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3330_));
AND2X2 AND2X2_2661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3331_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3329_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__10_));
AND2X2 AND2X2_2662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3334_));
AND2X2 AND2X2_2663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3335_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3333_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__11_));
AND2X2 AND2X2_2664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3338_));
AND2X2 AND2X2_2665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3339_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3337_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__12_));
AND2X2 AND2X2_2666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3342_));
AND2X2 AND2X2_2667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3343_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3341_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__13_));
AND2X2 AND2X2_2668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3346_));
AND2X2 AND2X2_2669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3347_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3345_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__14_));
AND2X2 AND2X2_267 ( .A(_abc_44694_new_n1095_), .B(opcode_q_22_), .Y(_abc_44694_new_n1105_));
AND2X2 AND2X2_2670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3350_));
AND2X2 AND2X2_2671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3351_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3349_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__15_));
AND2X2 AND2X2_2672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3354_));
AND2X2 AND2X2_2673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3355_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3353_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__16_));
AND2X2 AND2X2_2674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3358_));
AND2X2 AND2X2_2675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3359_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3357_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__17_));
AND2X2 AND2X2_2676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3362_));
AND2X2 AND2X2_2677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3363_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3361_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__18_));
AND2X2 AND2X2_2678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3366_));
AND2X2 AND2X2_2679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3365_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__19_));
AND2X2 AND2X2_268 ( .A(_abc_44694_new_n1106_), .B(opcode_q_24_), .Y(_abc_44694_new_n1107_));
AND2X2 AND2X2_2680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3370_));
AND2X2 AND2X2_2681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3371_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3369_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__20_));
AND2X2 AND2X2_2682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3374_));
AND2X2 AND2X2_2683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3375_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3373_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__21_));
AND2X2 AND2X2_2684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3378_));
AND2X2 AND2X2_2685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3379_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3377_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__22_));
AND2X2 AND2X2_2686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3382_));
AND2X2 AND2X2_2687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3383_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3381_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__23_));
AND2X2 AND2X2_2688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3386_));
AND2X2 AND2X2_2689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3387_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3385_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__24_));
AND2X2 AND2X2_269 ( .A(_abc_44694_new_n1093_), .B(_abc_44694_new_n1107_), .Y(_abc_44694_new_n1108_));
AND2X2 AND2X2_2690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3390_));
AND2X2 AND2X2_2691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3391_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3389_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__25_));
AND2X2 AND2X2_2692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3394_));
AND2X2 AND2X2_2693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3395_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3393_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__26_));
AND2X2 AND2X2_2694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3398_));
AND2X2 AND2X2_2695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3399_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3397_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__27_));
AND2X2 AND2X2_2696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3402_));
AND2X2 AND2X2_2697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3403_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3401_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__28_));
AND2X2 AND2X2_2698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3406_));
AND2X2 AND2X2_2699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3407_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3405_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__29_));
AND2X2 AND2X2_27 ( .A(mem_ack_i), .B(state_q_1_bF_buf4_), .Y(_abc_44694_new_n660_));
AND2X2 AND2X2_270 ( .A(_abc_44694_new_n1108_), .B(_abc_44694_new_n1105_), .Y(_abc_44694_new_n1109_));
AND2X2 AND2X2_2700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3410_));
AND2X2 AND2X2_2701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3411_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3409_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__30_));
AND2X2 AND2X2_2702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3414_));
AND2X2 AND2X2_2703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3415_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3413_), .Y(REGFILE_SIM_reg_bank__0reg_r21_31_0__31_));
AND2X2 AND2X2_2704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2467_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3417_));
AND2X2 AND2X2_2705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3420_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3418_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__0_));
AND2X2 AND2X2_2706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3423_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3422_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__1_));
AND2X2 AND2X2_2707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3426_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3425_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__2_));
AND2X2 AND2X2_2708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3429_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3428_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__3_));
AND2X2 AND2X2_2709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3432_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3431_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__4_));
AND2X2 AND2X2_271 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1109_), .Y(_abc_44694_new_n1110_));
AND2X2 AND2X2_2710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3435_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3434_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__5_));
AND2X2 AND2X2_2711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3438_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3437_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__6_));
AND2X2 AND2X2_2712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3441_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3440_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__7_));
AND2X2 AND2X2_2713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3444_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3443_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__8_));
AND2X2 AND2X2_2714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3447_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3446_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__9_));
AND2X2 AND2X2_2715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3450_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3449_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__10_));
AND2X2 AND2X2_2716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3453_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3452_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__11_));
AND2X2 AND2X2_2717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3456_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3455_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__12_));
AND2X2 AND2X2_2718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3459_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3458_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__13_));
AND2X2 AND2X2_2719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3462_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3461_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__14_));
AND2X2 AND2X2_272 ( .A(_abc_44694_new_n1083_), .B(_abc_44694_new_n647_), .Y(_abc_44694_new_n1114_));
AND2X2 AND2X2_2720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3465_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3464_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__15_));
AND2X2 AND2X2_2721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3468_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3467_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__16_));
AND2X2 AND2X2_2722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3470_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__17_));
AND2X2 AND2X2_2723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3474_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3473_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__18_));
AND2X2 AND2X2_2724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3477_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3476_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__19_));
AND2X2 AND2X2_2725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3480_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3479_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__20_));
AND2X2 AND2X2_2726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3483_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3482_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__21_));
AND2X2 AND2X2_2727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3486_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3485_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__22_));
AND2X2 AND2X2_2728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3489_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3488_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__23_));
AND2X2 AND2X2_2729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3492_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3491_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__24_));
AND2X2 AND2X2_273 ( .A(_abc_44694_new_n1017_), .B(_abc_44694_new_n1115_), .Y(_abc_44694_new_n1116_));
AND2X2 AND2X2_2730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3494_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__25_));
AND2X2 AND2X2_2731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3498_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3497_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__26_));
AND2X2 AND2X2_2732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3501_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3500_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__27_));
AND2X2 AND2X2_2733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3504_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3503_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__28_));
AND2X2 AND2X2_2734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3507_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3506_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__29_));
AND2X2 AND2X2_2735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3510_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3509_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__30_));
AND2X2 AND2X2_2736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3513_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3512_), .Y(REGFILE_SIM_reg_bank__0reg_r20_31_0__31_));
AND2X2 AND2X2_2737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3056_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2597_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3515_));
AND2X2 AND2X2_2738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2100_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3516_));
AND2X2 AND2X2_2739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3516_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3517_));
AND2X2 AND2X2_274 ( .A(_abc_44694_new_n619_), .B(_abc_44694_new_n639_), .Y(_abc_44694_new_n1117_));
AND2X2 AND2X2_2740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3520_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3518_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__0_));
AND2X2 AND2X2_2741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3523_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3522_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__1_));
AND2X2 AND2X2_2742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3526_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3525_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__2_));
AND2X2 AND2X2_2743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3529_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3528_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__3_));
AND2X2 AND2X2_2744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3532_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3531_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__4_));
AND2X2 AND2X2_2745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3535_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3534_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__5_));
AND2X2 AND2X2_2746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3538_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3537_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__6_));
AND2X2 AND2X2_2747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3541_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3540_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__7_));
AND2X2 AND2X2_2748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3544_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3543_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__8_));
AND2X2 AND2X2_2749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3547_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3546_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__9_));
AND2X2 AND2X2_275 ( .A(_abc_44694_new_n649_), .B(_abc_44694_new_n1117_), .Y(_abc_44694_new_n1118_));
AND2X2 AND2X2_2750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3550_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3549_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__10_));
AND2X2 AND2X2_2751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3553_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3552_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__11_));
AND2X2 AND2X2_2752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3555_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__12_));
AND2X2 AND2X2_2753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3559_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3558_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__13_));
AND2X2 AND2X2_2754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3562_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3561_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__14_));
AND2X2 AND2X2_2755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3565_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3564_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__15_));
AND2X2 AND2X2_2756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3568_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3567_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__16_));
AND2X2 AND2X2_2757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3571_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3570_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__17_));
AND2X2 AND2X2_2758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3574_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3573_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__18_));
AND2X2 AND2X2_2759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3577_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3576_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__19_));
AND2X2 AND2X2_276 ( .A(_abc_44694_new_n639_), .B(_abc_44694_new_n647_), .Y(_abc_44694_new_n1119_));
AND2X2 AND2X2_2760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3580_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3579_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__20_));
AND2X2 AND2X2_2761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3583_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3582_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__21_));
AND2X2 AND2X2_2762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3586_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3585_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__22_));
AND2X2 AND2X2_2763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3589_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3588_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__23_));
AND2X2 AND2X2_2764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3592_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3591_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__24_));
AND2X2 AND2X2_2765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3595_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3594_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__25_));
AND2X2 AND2X2_2766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3598_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3597_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__26_));
AND2X2 AND2X2_2767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3601_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3600_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__27_));
AND2X2 AND2X2_2768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3604_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3603_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__28_));
AND2X2 AND2X2_2769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3607_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3606_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__29_));
AND2X2 AND2X2_277 ( .A(_abc_44694_new_n618_), .B(inst_r_4_), .Y(_abc_44694_new_n1120_));
AND2X2 AND2X2_2770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3610_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3609_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__30_));
AND2X2 AND2X2_2771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3613_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3612_), .Y(REGFILE_SIM_reg_bank__0reg_r19_31_0__31_));
AND2X2 AND2X2_2772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2265_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3615_));
AND2X2 AND2X2_2773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3615_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3616_));
AND2X2 AND2X2_2774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3619_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3617_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__0_));
AND2X2 AND2X2_2775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3622_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3621_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__1_));
AND2X2 AND2X2_2776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3625_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3624_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__2_));
AND2X2 AND2X2_2777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3628_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3627_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__3_));
AND2X2 AND2X2_2778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3631_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3630_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__4_));
AND2X2 AND2X2_2779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3634_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3633_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__5_));
AND2X2 AND2X2_278 ( .A(_abc_44694_new_n1119_), .B(_abc_44694_new_n1120_), .Y(_abc_44694_new_n1121_));
AND2X2 AND2X2_2780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3637_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3636_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__6_));
AND2X2 AND2X2_2781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3640_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3639_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__7_));
AND2X2 AND2X2_2782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3643_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3642_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__8_));
AND2X2 AND2X2_2783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3646_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3645_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__9_));
AND2X2 AND2X2_2784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3649_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3648_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__10_));
AND2X2 AND2X2_2785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3652_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3651_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__11_));
AND2X2 AND2X2_2786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3655_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3654_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__12_));
AND2X2 AND2X2_2787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3658_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3657_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__13_));
AND2X2 AND2X2_2788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3661_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3660_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__14_));
AND2X2 AND2X2_2789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3664_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3663_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__15_));
AND2X2 AND2X2_279 ( .A(_abc_44694_new_n619_), .B(_abc_44694_new_n632_), .Y(_abc_44694_new_n1122_));
AND2X2 AND2X2_2790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3667_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3666_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__16_));
AND2X2 AND2X2_2791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3670_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3669_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__17_));
AND2X2 AND2X2_2792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3673_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3672_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__18_));
AND2X2 AND2X2_2793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3676_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3675_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__19_));
AND2X2 AND2X2_2794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3679_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3678_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__20_));
AND2X2 AND2X2_2795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3682_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3681_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__21_));
AND2X2 AND2X2_2796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3685_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3684_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__22_));
AND2X2 AND2X2_2797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3688_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3687_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__23_));
AND2X2 AND2X2_2798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3691_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3690_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__24_));
AND2X2 AND2X2_2799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3694_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3693_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__25_));
AND2X2 AND2X2_28 ( .A(_abc_44694_new_n661_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n662_));
AND2X2 AND2X2_280 ( .A(_abc_44694_new_n1122_), .B(_abc_44694_new_n624_), .Y(_abc_44694_new_n1123_));
AND2X2 AND2X2_2800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3697_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3696_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__26_));
AND2X2 AND2X2_2801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3700_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3699_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__27_));
AND2X2 AND2X2_2802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3703_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3702_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__28_));
AND2X2 AND2X2_2803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3706_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3705_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__29_));
AND2X2 AND2X2_2804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3709_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3708_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__30_));
AND2X2 AND2X2_2805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3712_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3711_), .Y(REGFILE_SIM_reg_bank__0reg_r18_31_0__31_));
AND2X2 AND2X2_2806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2366_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3714_));
AND2X2 AND2X2_2807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3714_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3715_));
AND2X2 AND2X2_2808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3718_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3716_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__0_));
AND2X2 AND2X2_2809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3721_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3720_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__1_));
AND2X2 AND2X2_281 ( .A(_abc_44694_new_n1126_), .B(_abc_44694_new_n1116_), .Y(_abc_44694_new_n1127_));
AND2X2 AND2X2_2810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3724_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3723_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__2_));
AND2X2 AND2X2_2811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3727_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3726_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__3_));
AND2X2 AND2X2_2812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3730_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3729_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__4_));
AND2X2 AND2X2_2813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3733_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3732_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__5_));
AND2X2 AND2X2_2814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3736_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3735_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__6_));
AND2X2 AND2X2_2815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3739_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3738_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__7_));
AND2X2 AND2X2_2816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3742_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3741_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__8_));
AND2X2 AND2X2_2817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3745_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3744_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__9_));
AND2X2 AND2X2_2818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3748_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3747_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__10_));
AND2X2 AND2X2_2819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3751_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3750_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__11_));
AND2X2 AND2X2_282 ( .A(_abc_44694_new_n1093_), .B(_abc_44694_new_n1129_), .Y(_abc_44694_new_n1130_));
AND2X2 AND2X2_2820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3754_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3753_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__12_));
AND2X2 AND2X2_2821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3757_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3756_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__13_));
AND2X2 AND2X2_2822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3760_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3759_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__14_));
AND2X2 AND2X2_2823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3763_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3762_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__15_));
AND2X2 AND2X2_2824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3766_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3765_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__16_));
AND2X2 AND2X2_2825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3769_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3768_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__17_));
AND2X2 AND2X2_2826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3772_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3771_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__18_));
AND2X2 AND2X2_2827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3775_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3774_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__19_));
AND2X2 AND2X2_2828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3778_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3777_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__20_));
AND2X2 AND2X2_2829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3781_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3780_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__21_));
AND2X2 AND2X2_283 ( .A(_abc_44694_new_n1130_), .B(_abc_44694_new_n1090_), .Y(_abc_44694_new_n1131_));
AND2X2 AND2X2_2830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3784_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3783_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__22_));
AND2X2 AND2X2_2831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3787_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3786_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__23_));
AND2X2 AND2X2_2832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3790_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3789_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__24_));
AND2X2 AND2X2_2833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3793_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3792_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__25_));
AND2X2 AND2X2_2834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3796_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3795_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__26_));
AND2X2 AND2X2_2835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3799_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3798_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__27_));
AND2X2 AND2X2_2836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3802_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3801_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__28_));
AND2X2 AND2X2_2837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3805_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3804_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__29_));
AND2X2 AND2X2_2838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3808_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3807_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__30_));
AND2X2 AND2X2_2839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3811_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3810_), .Y(REGFILE_SIM_reg_bank__0reg_r17_31_0__31_));
AND2X2 AND2X2_284 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1131_), .Y(_abc_44694_new_n1132_));
AND2X2 AND2X2_2840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2467_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3515_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3813_));
AND2X2 AND2X2_2841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3816_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3814_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__0_));
AND2X2 AND2X2_2842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3819_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3818_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__1_));
AND2X2 AND2X2_2843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3822_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3821_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__2_));
AND2X2 AND2X2_2844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3825_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3824_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__3_));
AND2X2 AND2X2_2845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3828_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3827_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__4_));
AND2X2 AND2X2_2846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3831_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3830_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__5_));
AND2X2 AND2X2_2847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3834_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3833_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__6_));
AND2X2 AND2X2_2848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3837_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3836_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__7_));
AND2X2 AND2X2_2849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3840_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3839_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__8_));
AND2X2 AND2X2_285 ( .A(opcode_q_22_), .B(opcode_q_21_), .Y(_abc_44694_new_n1134_));
AND2X2 AND2X2_2850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3843_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3842_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__9_));
AND2X2 AND2X2_2851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3846_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3845_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__10_));
AND2X2 AND2X2_2852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3849_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3848_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__11_));
AND2X2 AND2X2_2853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3852_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3851_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__12_));
AND2X2 AND2X2_2854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3855_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3854_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__13_));
AND2X2 AND2X2_2855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3858_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3857_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__14_));
AND2X2 AND2X2_2856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3861_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3860_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__15_));
AND2X2 AND2X2_2857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3864_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3863_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__16_));
AND2X2 AND2X2_2858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3867_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3866_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__17_));
AND2X2 AND2X2_2859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3870_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3869_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__18_));
AND2X2 AND2X2_286 ( .A(_abc_44694_new_n1108_), .B(_abc_44694_new_n1134_), .Y(_abc_44694_new_n1135_));
AND2X2 AND2X2_2860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3873_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3872_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__19_));
AND2X2 AND2X2_2861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3876_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3875_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__20_));
AND2X2 AND2X2_2862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3879_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3878_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__21_));
AND2X2 AND2X2_2863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3882_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3881_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__22_));
AND2X2 AND2X2_2864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3885_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3884_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__23_));
AND2X2 AND2X2_2865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3888_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3887_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__24_));
AND2X2 AND2X2_2866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3891_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3890_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__25_));
AND2X2 AND2X2_2867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3894_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3893_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__26_));
AND2X2 AND2X2_2868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3897_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3896_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__27_));
AND2X2 AND2X2_2869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3900_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3899_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__28_));
AND2X2 AND2X2_287 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1135_), .Y(_abc_44694_new_n1136_));
AND2X2 AND2X2_2870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3903_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3902_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__29_));
AND2X2 AND2X2_2871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3906_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3905_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__30_));
AND2X2 AND2X2_2872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3909_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3908_), .Y(REGFILE_SIM_reg_bank__0reg_r16_31_0__31_));
AND2X2 AND2X2_2873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3911_), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3912_));
AND2X2 AND2X2_2874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2101_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913_));
AND2X2 AND2X2_2875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3915_));
AND2X2 AND2X2_2876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3916_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3914_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__0_));
AND2X2 AND2X2_2877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3919_));
AND2X2 AND2X2_2878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3920_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3918_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__1_));
AND2X2 AND2X2_2879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3923_));
AND2X2 AND2X2_288 ( .A(_abc_44694_new_n1137_), .B(_abc_44694_new_n1133_), .Y(_abc_44694_new_n1138_));
AND2X2 AND2X2_2880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3924_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3922_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__2_));
AND2X2 AND2X2_2881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3927_));
AND2X2 AND2X2_2882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3928_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3926_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__3_));
AND2X2 AND2X2_2883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3931_));
AND2X2 AND2X2_2884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3932_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3930_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__4_));
AND2X2 AND2X2_2885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3935_));
AND2X2 AND2X2_2886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3936_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3934_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__5_));
AND2X2 AND2X2_2887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3939_));
AND2X2 AND2X2_2888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3940_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3938_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__6_));
AND2X2 AND2X2_2889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3943_));
AND2X2 AND2X2_289 ( .A(_abc_44694_new_n1138_), .B(_abc_44694_new_n1127_), .Y(_abc_44694_new_n1139_));
AND2X2 AND2X2_2890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3944_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3942_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__7_));
AND2X2 AND2X2_2891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3947_));
AND2X2 AND2X2_2892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3948_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3946_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__8_));
AND2X2 AND2X2_2893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3951_));
AND2X2 AND2X2_2894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3952_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3950_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__9_));
AND2X2 AND2X2_2895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3955_));
AND2X2 AND2X2_2896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3956_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3954_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__10_));
AND2X2 AND2X2_2897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3959_));
AND2X2 AND2X2_2898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3960_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3958_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__11_));
AND2X2 AND2X2_2899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3963_));
AND2X2 AND2X2_29 ( .A(_abc_44694_new_n664_), .B(state_q_2_), .Y(_abc_44694_new_n665_));
AND2X2 AND2X2_290 ( .A(_abc_44694_new_n1113_), .B(_abc_44694_new_n1139_), .Y(_abc_44694_new_n1140_));
AND2X2 AND2X2_2900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3964_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3962_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__12_));
AND2X2 AND2X2_2901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3967_));
AND2X2 AND2X2_2902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3968_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3966_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__13_));
AND2X2 AND2X2_2903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3971_));
AND2X2 AND2X2_2904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3972_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3970_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__14_));
AND2X2 AND2X2_2905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3975_));
AND2X2 AND2X2_2906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3976_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3974_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__15_));
AND2X2 AND2X2_2907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3979_));
AND2X2 AND2X2_2908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3980_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3978_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__16_));
AND2X2 AND2X2_2909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3983_));
AND2X2 AND2X2_291 ( .A(_abc_44694_new_n1140_), .B(_abc_44694_new_n1081_), .Y(_abc_44694_new_n1141_));
AND2X2 AND2X2_2910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3984_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3982_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__17_));
AND2X2 AND2X2_2911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3987_));
AND2X2 AND2X2_2912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3988_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3986_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__18_));
AND2X2 AND2X2_2913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3991_));
AND2X2 AND2X2_2914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3992_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3990_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__19_));
AND2X2 AND2X2_2915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3995_));
AND2X2 AND2X2_2916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3996_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3994_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__20_));
AND2X2 AND2X2_2917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3999_));
AND2X2 AND2X2_2918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4000_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3998_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__21_));
AND2X2 AND2X2_2919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4003_));
AND2X2 AND2X2_292 ( .A(_abc_44694_new_n1083_), .B(_abc_44694_new_n645_), .Y(_abc_44694_new_n1142_));
AND2X2 AND2X2_2920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4004_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4002_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__22_));
AND2X2 AND2X2_2921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4007_));
AND2X2 AND2X2_2922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4008_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4006_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__23_));
AND2X2 AND2X2_2923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4011_));
AND2X2 AND2X2_2924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4012_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4010_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__24_));
AND2X2 AND2X2_2925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4015_));
AND2X2 AND2X2_2926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4016_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4014_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__25_));
AND2X2 AND2X2_2927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4019_));
AND2X2 AND2X2_2928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4020_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4018_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__26_));
AND2X2 AND2X2_2929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4023_));
AND2X2 AND2X2_293 ( .A(_abc_44694_new_n1057_), .B(alu_op_r_4_), .Y(_abc_44694_new_n1143_));
AND2X2 AND2X2_2930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4024_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4022_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__27_));
AND2X2 AND2X2_2931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4027_));
AND2X2 AND2X2_2932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4028_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4026_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__28_));
AND2X2 AND2X2_2933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4031_));
AND2X2 AND2X2_2934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4032_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4030_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__29_));
AND2X2 AND2X2_2935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4035_));
AND2X2 AND2X2_2936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4036_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4034_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__30_));
AND2X2 AND2X2_2937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4039_));
AND2X2 AND2X2_2938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4040_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4038_), .Y(REGFILE_SIM_reg_bank__0reg_r15_31_0__31_));
AND2X2 AND2X2_2939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2266_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4042_));
AND2X2 AND2X2_294 ( .A(_abc_44694_new_n1142_), .B(_abc_44694_new_n1143_), .Y(_abc_44694_new_n1144_));
AND2X2 AND2X2_2940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4045_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4043_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__0_));
AND2X2 AND2X2_2941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4048_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4047_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__1_));
AND2X2 AND2X2_2942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4051_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4050_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__2_));
AND2X2 AND2X2_2943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4053_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__3_));
AND2X2 AND2X2_2944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4057_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4056_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__4_));
AND2X2 AND2X2_2945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4060_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4059_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__5_));
AND2X2 AND2X2_2946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4063_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4062_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__6_));
AND2X2 AND2X2_2947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4066_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4065_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__7_));
AND2X2 AND2X2_2948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4069_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4068_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__8_));
AND2X2 AND2X2_2949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4072_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4071_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__9_));
AND2X2 AND2X2_295 ( .A(_abc_44694_new_n621_), .B(_abc_44694_new_n637_), .Y(_abc_44694_new_n1145_));
AND2X2 AND2X2_2950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4075_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4074_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__10_));
AND2X2 AND2X2_2951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4078_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4077_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__11_));
AND2X2 AND2X2_2952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4081_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4080_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__12_));
AND2X2 AND2X2_2953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4084_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4083_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__13_));
AND2X2 AND2X2_2954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4087_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4086_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__14_));
AND2X2 AND2X2_2955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4090_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4089_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__15_));
AND2X2 AND2X2_2956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4093_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4092_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__16_));
AND2X2 AND2X2_2957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4096_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4095_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__17_));
AND2X2 AND2X2_2958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4099_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4098_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__18_));
AND2X2 AND2X2_2959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4102_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4101_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__19_));
AND2X2 AND2X2_296 ( .A(_abc_44694_new_n1145_), .B(_abc_44694_new_n638_), .Y(_abc_44694_new_n1146_));
AND2X2 AND2X2_2960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4105_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4104_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__20_));
AND2X2 AND2X2_2961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4108_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4107_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__21_));
AND2X2 AND2X2_2962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4111_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4110_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__22_));
AND2X2 AND2X2_2963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4114_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4113_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__23_));
AND2X2 AND2X2_2964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4117_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4116_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__24_));
AND2X2 AND2X2_2965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4120_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4119_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__25_));
AND2X2 AND2X2_2966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4123_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4122_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__26_));
AND2X2 AND2X2_2967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4126_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4125_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__27_));
AND2X2 AND2X2_2968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4129_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4128_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__28_));
AND2X2 AND2X2_2969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4132_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4131_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__29_));
AND2X2 AND2X2_297 ( .A(_abc_44694_new_n1142_), .B(_abc_44694_new_n1056_), .Y(_abc_44694_new_n1147_));
AND2X2 AND2X2_2970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4135_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4134_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__30_));
AND2X2 AND2X2_2971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4138_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4137_), .Y(REGFILE_SIM_reg_bank__0reg_r14_31_0__31_));
AND2X2 AND2X2_2972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4140_));
AND2X2 AND2X2_2973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4143_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4141_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__0_));
AND2X2 AND2X2_2974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4146_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4145_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__1_));
AND2X2 AND2X2_2975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4149_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4148_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__2_));
AND2X2 AND2X2_2976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4152_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4151_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__3_));
AND2X2 AND2X2_2977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4155_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4154_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__4_));
AND2X2 AND2X2_2978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4158_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4157_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__5_));
AND2X2 AND2X2_2979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4161_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4160_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__6_));
AND2X2 AND2X2_298 ( .A(_abc_44694_new_n1061_), .B(_abc_44694_new_n1143_), .Y(_abc_44694_new_n1150_));
AND2X2 AND2X2_2980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4164_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4163_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__7_));
AND2X2 AND2X2_2981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4167_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4166_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__8_));
AND2X2 AND2X2_2982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4170_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4169_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__9_));
AND2X2 AND2X2_2983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4173_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4172_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__10_));
AND2X2 AND2X2_2984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4176_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4175_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__11_));
AND2X2 AND2X2_2985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4179_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4178_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__12_));
AND2X2 AND2X2_2986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4182_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4181_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__13_));
AND2X2 AND2X2_2987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4185_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4184_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__14_));
AND2X2 AND2X2_2988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4188_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4187_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__15_));
AND2X2 AND2X2_2989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4191_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4190_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__16_));
AND2X2 AND2X2_299 ( .A(_abc_44694_new_n1101_), .B(_abc_44694_new_n1150_), .Y(_abc_44694_new_n1151_));
AND2X2 AND2X2_2990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4194_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4193_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__17_));
AND2X2 AND2X2_2991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4197_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4196_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__18_));
AND2X2 AND2X2_2992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4200_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4199_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__19_));
AND2X2 AND2X2_2993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4203_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4202_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__20_));
AND2X2 AND2X2_2994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4206_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4205_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__21_));
AND2X2 AND2X2_2995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4209_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4208_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__22_));
AND2X2 AND2X2_2996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4212_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4211_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__23_));
AND2X2 AND2X2_2997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4215_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4214_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__24_));
AND2X2 AND2X2_2998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4218_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4217_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__25_));
AND2X2 AND2X2_2999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4221_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4220_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__26_));
AND2X2 AND2X2_3 ( .A(_abc_44694_new_n619_), .B(_abc_44694_new_n621_), .Y(_abc_44694_new_n622_));
AND2X2 AND2X2_30 ( .A(_abc_44694_new_n667_), .B(state_q_5_bF_buf2_), .Y(_abc_44694_new_n668_));
AND2X2 AND2X2_300 ( .A(_abc_44694_new_n1151_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n1152_));
AND2X2 AND2X2_3000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4224_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4223_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__27_));
AND2X2 AND2X2_3001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4226_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__28_));
AND2X2 AND2X2_3002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4230_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4229_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__29_));
AND2X2 AND2X2_3003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4233_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4232_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__30_));
AND2X2 AND2X2_3004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4236_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4235_), .Y(REGFILE_SIM_reg_bank__0reg_r13_31_0__31_));
AND2X2 AND2X2_3005 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2466_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4238_));
AND2X2 AND2X2_3006 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4238_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2099_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4239_));
AND2X2 AND2X2_3007 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4242_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4240_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__0_));
AND2X2 AND2X2_3008 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4245_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4244_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__1_));
AND2X2 AND2X2_3009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4248_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4247_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__2_));
AND2X2 AND2X2_301 ( .A(_abc_44694_new_n1068_), .B(_abc_44694_new_n1073_), .Y(_abc_44694_new_n1153_));
AND2X2 AND2X2_3010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4251_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4250_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__3_));
AND2X2 AND2X2_3011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4254_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4253_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__4_));
AND2X2 AND2X2_3012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4256_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__5_));
AND2X2 AND2X2_3013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4260_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4259_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__6_));
AND2X2 AND2X2_3014 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4263_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4262_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__7_));
AND2X2 AND2X2_3015 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4266_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4265_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__8_));
AND2X2 AND2X2_3016 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4269_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4268_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__9_));
AND2X2 AND2X2_3017 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4272_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4271_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__10_));
AND2X2 AND2X2_3018 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4275_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4274_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__11_));
AND2X2 AND2X2_3019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4278_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4277_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__12_));
AND2X2 AND2X2_302 ( .A(_abc_44694_new_n1062_), .B(_abc_44694_new_n1153_), .Y(_abc_44694_new_n1154_));
AND2X2 AND2X2_3020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4281_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4280_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__13_));
AND2X2 AND2X2_3021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4284_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4283_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__14_));
AND2X2 AND2X2_3022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4287_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4286_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__15_));
AND2X2 AND2X2_3023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4290_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4289_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__16_));
AND2X2 AND2X2_3024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4293_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4292_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__17_));
AND2X2 AND2X2_3025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4296_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4295_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__18_));
AND2X2 AND2X2_3026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4299_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4298_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__19_));
AND2X2 AND2X2_3027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4302_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4301_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__20_));
AND2X2 AND2X2_3028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4305_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4304_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__21_));
AND2X2 AND2X2_3029 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4308_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4307_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__22_));
AND2X2 AND2X2_303 ( .A(_abc_44694_new_n1154_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n1155_));
AND2X2 AND2X2_3030 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4311_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4310_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__23_));
AND2X2 AND2X2_3031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4314_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4313_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__24_));
AND2X2 AND2X2_3032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4317_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4316_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__25_));
AND2X2 AND2X2_3033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4320_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4319_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__26_));
AND2X2 AND2X2_3034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4323_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4322_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__27_));
AND2X2 AND2X2_3035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4326_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4325_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__28_));
AND2X2 AND2X2_3036 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4329_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4328_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__29_));
AND2X2 AND2X2_3037 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4332_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4331_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__30_));
AND2X2 AND2X2_3038 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4335_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4334_), .Y(REGFILE_SIM_reg_bank__0reg_r12_31_0__31_));
AND2X2 AND2X2_3039 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2599_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4337_));
AND2X2 AND2X2_304 ( .A(_abc_44694_new_n1063_), .B(alu_op_r_1_), .Y(_abc_44694_new_n1156_));
AND2X2 AND2X2_3040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4340_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4338_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__0_));
AND2X2 AND2X2_3041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4343_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4342_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__1_));
AND2X2 AND2X2_3042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4346_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4345_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__2_));
AND2X2 AND2X2_3043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4349_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4348_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__3_));
AND2X2 AND2X2_3044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4352_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4351_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__4_));
AND2X2 AND2X2_3045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4355_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4354_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__5_));
AND2X2 AND2X2_3046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4358_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4357_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__6_));
AND2X2 AND2X2_3047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4361_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4360_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__7_));
AND2X2 AND2X2_3048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4364_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4363_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__8_));
AND2X2 AND2X2_3049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4366_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__9_));
AND2X2 AND2X2_305 ( .A(_abc_44694_new_n1055_), .B(_abc_44694_new_n1156_), .Y(_abc_44694_new_n1157_));
AND2X2 AND2X2_3050 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4370_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4369_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__10_));
AND2X2 AND2X2_3051 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4373_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4372_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__11_));
AND2X2 AND2X2_3052 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4376_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4375_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__12_));
AND2X2 AND2X2_3053 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4379_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4378_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__13_));
AND2X2 AND2X2_3054 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4382_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4381_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__14_));
AND2X2 AND2X2_3055 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4385_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4384_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__15_));
AND2X2 AND2X2_3056 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4388_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4387_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__16_));
AND2X2 AND2X2_3057 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4391_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4390_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__17_));
AND2X2 AND2X2_3058 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4394_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4393_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__18_));
AND2X2 AND2X2_3059 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4397_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4396_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__19_));
AND2X2 AND2X2_306 ( .A(_abc_44694_new_n1062_), .B(_abc_44694_new_n1157_), .Y(_abc_44694_new_n1158_));
AND2X2 AND2X2_3060 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4400_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4399_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__20_));
AND2X2 AND2X2_3061 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4403_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4402_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__21_));
AND2X2 AND2X2_3062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4406_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4405_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__22_));
AND2X2 AND2X2_3063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4409_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4408_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__23_));
AND2X2 AND2X2_3064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4412_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4411_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__24_));
AND2X2 AND2X2_3065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4415_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4414_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__25_));
AND2X2 AND2X2_3066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4418_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4417_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__26_));
AND2X2 AND2X2_3067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4421_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4420_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__27_));
AND2X2 AND2X2_3068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4424_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4423_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__28_));
AND2X2 AND2X2_3069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4427_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4426_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__29_));
AND2X2 AND2X2_307 ( .A(_abc_44694_new_n1158_), .B(_abc_44694_new_n1052_), .Y(_abc_44694_new_n1159_));
AND2X2 AND2X2_3070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4430_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4429_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__30_));
AND2X2 AND2X2_3071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4433_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4432_), .Y(REGFILE_SIM_reg_bank__0reg_r11_31_0__31_));
AND2X2 AND2X2_3072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2698_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435_));
AND2X2 AND2X2_3073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4437_));
AND2X2 AND2X2_3074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4438_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4436_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__0_));
AND2X2 AND2X2_3075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4441_));
AND2X2 AND2X2_3076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4442_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4440_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__1_));
AND2X2 AND2X2_3077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4445_));
AND2X2 AND2X2_3078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4446_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4444_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__2_));
AND2X2 AND2X2_3079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4449_));
AND2X2 AND2X2_308 ( .A(opcode_q_24_), .B(opcode_q_23_), .Y(_abc_44694_new_n1164_));
AND2X2 AND2X2_3080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4450_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4448_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__3_));
AND2X2 AND2X2_3081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4453_));
AND2X2 AND2X2_3082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4454_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4452_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__4_));
AND2X2 AND2X2_3083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4457_));
AND2X2 AND2X2_3084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4458_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4456_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__5_));
AND2X2 AND2X2_3085 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4461_));
AND2X2 AND2X2_3086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4462_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4460_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__6_));
AND2X2 AND2X2_3087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4465_));
AND2X2 AND2X2_3088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4466_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4464_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__7_));
AND2X2 AND2X2_3089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4469_));
AND2X2 AND2X2_309 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1164_), .Y(_abc_44694_new_n1165_));
AND2X2 AND2X2_3090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4470_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4468_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__8_));
AND2X2 AND2X2_3091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4473_));
AND2X2 AND2X2_3092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4474_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4472_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__9_));
AND2X2 AND2X2_3093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4477_));
AND2X2 AND2X2_3094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4478_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4476_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__10_));
AND2X2 AND2X2_3095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4481_));
AND2X2 AND2X2_3096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4482_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4480_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__11_));
AND2X2 AND2X2_3097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4485_));
AND2X2 AND2X2_3098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4486_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4484_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__12_));
AND2X2 AND2X2_3099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4489_));
AND2X2 AND2X2_31 ( .A(_abc_44694_new_n664_), .B(state_q_1_bF_buf3_), .Y(_abc_44694_new_n669_));
AND2X2 AND2X2_310 ( .A(_abc_44694_new_n1165_), .B(_abc_44694_new_n1130_), .Y(_abc_44694_new_n1166_));
AND2X2 AND2X2_3100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4490_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4488_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__13_));
AND2X2 AND2X2_3101 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4493_));
AND2X2 AND2X2_3102 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4494_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4492_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__14_));
AND2X2 AND2X2_3103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4497_));
AND2X2 AND2X2_3104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4498_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4496_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__15_));
AND2X2 AND2X2_3105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4501_));
AND2X2 AND2X2_3106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4502_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4500_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__16_));
AND2X2 AND2X2_3107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4505_));
AND2X2 AND2X2_3108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4506_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4504_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__17_));
AND2X2 AND2X2_3109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4509_));
AND2X2 AND2X2_311 ( .A(_abc_44694_new_n1046_), .B(_abc_44694_new_n1106_), .Y(_abc_44694_new_n1167_));
AND2X2 AND2X2_3110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4510_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4508_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__18_));
AND2X2 AND2X2_3111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4513_));
AND2X2 AND2X2_3112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4514_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4512_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__19_));
AND2X2 AND2X2_3113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4517_));
AND2X2 AND2X2_3114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4518_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4516_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__20_));
AND2X2 AND2X2_3115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4521_));
AND2X2 AND2X2_3116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4522_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4520_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__21_));
AND2X2 AND2X2_3117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4525_));
AND2X2 AND2X2_3118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4526_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4524_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__22_));
AND2X2 AND2X2_3119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4529_));
AND2X2 AND2X2_312 ( .A(_abc_44694_new_n1093_), .B(_abc_44694_new_n1167_), .Y(_abc_44694_new_n1168_));
AND2X2 AND2X2_3120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4530_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4528_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__23_));
AND2X2 AND2X2_3121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4533_));
AND2X2 AND2X2_3122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4534_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4532_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__24_));
AND2X2 AND2X2_3123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4537_));
AND2X2 AND2X2_3124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4538_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4536_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__25_));
AND2X2 AND2X2_3125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4541_));
AND2X2 AND2X2_3126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4542_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4540_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__26_));
AND2X2 AND2X2_3127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4545_));
AND2X2 AND2X2_3128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4546_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4544_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__27_));
AND2X2 AND2X2_3129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4549_));
AND2X2 AND2X2_313 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1168_), .Y(_abc_44694_new_n1169_));
AND2X2 AND2X2_3130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4550_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4548_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__28_));
AND2X2 AND2X2_3131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4553_));
AND2X2 AND2X2_3132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4554_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4552_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__29_));
AND2X2 AND2X2_3133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4557_));
AND2X2 AND2X2_3134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4558_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4556_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__30_));
AND2X2 AND2X2_3135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4561_));
AND2X2 AND2X2_3136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4562_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4560_), .Y(REGFILE_SIM_reg_bank__0reg_r10_31_0__31_));
AND2X2 AND2X2_3137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3714_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4564_));
AND2X2 AND2X2_3138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4567_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4565_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__0_));
AND2X2 AND2X2_3139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4570_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4569_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__1_));
AND2X2 AND2X2_314 ( .A(_abc_44694_new_n1169_), .B(_abc_44694_new_n1095_), .Y(_abc_44694_new_n1170_));
AND2X2 AND2X2_3140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4573_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4572_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__2_));
AND2X2 AND2X2_3141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4576_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4575_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__3_));
AND2X2 AND2X2_3142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4579_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4578_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__4_));
AND2X2 AND2X2_3143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4582_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4581_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__5_));
AND2X2 AND2X2_3144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4585_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4584_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__6_));
AND2X2 AND2X2_3145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4588_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4587_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__7_));
AND2X2 AND2X2_3146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4591_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4590_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__8_));
AND2X2 AND2X2_3147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4594_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4593_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__9_));
AND2X2 AND2X2_3148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4597_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4596_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__10_));
AND2X2 AND2X2_3149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4600_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4599_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__11_));
AND2X2 AND2X2_315 ( .A(_abc_44694_new_n1169_), .B(_abc_44694_new_n1134_), .Y(_abc_44694_new_n1173_));
AND2X2 AND2X2_3150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4603_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4602_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__12_));
AND2X2 AND2X2_3151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4606_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4605_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__13_));
AND2X2 AND2X2_3152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4609_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4608_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__14_));
AND2X2 AND2X2_3153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4612_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4611_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__15_));
AND2X2 AND2X2_3154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4615_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4614_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__16_));
AND2X2 AND2X2_3155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4618_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4617_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__17_));
AND2X2 AND2X2_3156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4621_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4620_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__18_));
AND2X2 AND2X2_3157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4623_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__19_));
AND2X2 AND2X2_3158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4627_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4626_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__20_));
AND2X2 AND2X2_3159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4630_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4629_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__21_));
AND2X2 AND2X2_316 ( .A(_abc_44694_new_n639_), .B(_abc_44694_new_n645_), .Y(_abc_44694_new_n1175_));
AND2X2 AND2X2_3160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4633_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4632_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__22_));
AND2X2 AND2X2_3161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4636_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4635_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__23_));
AND2X2 AND2X2_3162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4639_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4638_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__24_));
AND2X2 AND2X2_3163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4642_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4641_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__25_));
AND2X2 AND2X2_3164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4645_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4644_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__26_));
AND2X2 AND2X2_3165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4648_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4647_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__27_));
AND2X2 AND2X2_3166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4651_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4650_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__28_));
AND2X2 AND2X2_3167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4654_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4653_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__29_));
AND2X2 AND2X2_3168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4657_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4656_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__30_));
AND2X2 AND2X2_3169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4660_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4659_), .Y(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__31_));
AND2X2 AND2X2_317 ( .A(_abc_44694_new_n1175_), .B(_abc_44694_new_n1120_), .Y(_abc_44694_new_n1176_));
AND2X2 AND2X2_3170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2828_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662_));
AND2X2 AND2X2_3171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4664_));
AND2X2 AND2X2_3172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4665_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4663_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__0_));
AND2X2 AND2X2_3173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4668_));
AND2X2 AND2X2_3174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4669_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4667_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__1_));
AND2X2 AND2X2_3175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4672_));
AND2X2 AND2X2_3176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4673_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4671_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__2_));
AND2X2 AND2X2_3177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4676_));
AND2X2 AND2X2_3178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4677_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4675_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__3_));
AND2X2 AND2X2_3179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4680_));
AND2X2 AND2X2_318 ( .A(_abc_44694_new_n1119_), .B(_abc_44694_new_n619_), .Y(_abc_44694_new_n1177_));
AND2X2 AND2X2_3180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4681_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4679_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__4_));
AND2X2 AND2X2_3181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4684_));
AND2X2 AND2X2_3182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4685_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4683_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__5_));
AND2X2 AND2X2_3183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4688_));
AND2X2 AND2X2_3184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4689_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4687_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__6_));
AND2X2 AND2X2_3185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4692_));
AND2X2 AND2X2_3186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4693_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4691_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__7_));
AND2X2 AND2X2_3187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4696_));
AND2X2 AND2X2_3188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4697_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4695_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__8_));
AND2X2 AND2X2_3189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4700_));
AND2X2 AND2X2_319 ( .A(_abc_44694_new_n632_), .B(_abc_44694_new_n638_), .Y(_abc_44694_new_n1180_));
AND2X2 AND2X2_3190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4701_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4699_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__9_));
AND2X2 AND2X2_3191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4704_));
AND2X2 AND2X2_3192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4705_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4703_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__10_));
AND2X2 AND2X2_3193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4708_));
AND2X2 AND2X2_3194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4709_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4707_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__11_));
AND2X2 AND2X2_3195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4712_));
AND2X2 AND2X2_3196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4713_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4711_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__12_));
AND2X2 AND2X2_3197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4716_));
AND2X2 AND2X2_3198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4717_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4715_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__13_));
AND2X2 AND2X2_3199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4720_));
AND2X2 AND2X2_32 ( .A(_abc_44694_new_n671_), .B(alu_p_o_0_), .Y(_abc_44694_new_n672_));
AND2X2 AND2X2_320 ( .A(_abc_44694_new_n1180_), .B(_abc_44694_new_n637_), .Y(_abc_44694_new_n1181_));
AND2X2 AND2X2_3200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4721_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4719_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__14_));
AND2X2 AND2X2_3201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4724_));
AND2X2 AND2X2_3202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4725_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4723_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__15_));
AND2X2 AND2X2_3203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4728_));
AND2X2 AND2X2_3204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4729_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4727_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__16_));
AND2X2 AND2X2_3205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4732_));
AND2X2 AND2X2_3206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4733_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4731_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__17_));
AND2X2 AND2X2_3207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4736_));
AND2X2 AND2X2_3208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4737_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4735_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__18_));
AND2X2 AND2X2_3209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4740_));
AND2X2 AND2X2_321 ( .A(_abc_44694_new_n1018_), .B(_abc_44694_new_n637_), .Y(_abc_44694_new_n1182_));
AND2X2 AND2X2_3210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4741_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4739_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__19_));
AND2X2 AND2X2_3211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4744_));
AND2X2 AND2X2_3212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4745_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4743_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__20_));
AND2X2 AND2X2_3213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4748_));
AND2X2 AND2X2_3214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4749_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4747_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__21_));
AND2X2 AND2X2_3215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4752_));
AND2X2 AND2X2_3216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4753_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4751_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__22_));
AND2X2 AND2X2_3217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4756_));
AND2X2 AND2X2_3218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4757_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4755_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__23_));
AND2X2 AND2X2_3219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4760_));
AND2X2 AND2X2_322 ( .A(_abc_44694_new_n869_), .B(_abc_44694_new_n619_), .Y(_abc_44694_new_n1185_));
AND2X2 AND2X2_3220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4761_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4759_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__24_));
AND2X2 AND2X2_3221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4764_));
AND2X2 AND2X2_3222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4765_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4763_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__25_));
AND2X2 AND2X2_3223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4768_));
AND2X2 AND2X2_3224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4769_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4767_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__26_));
AND2X2 AND2X2_3225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4772_));
AND2X2 AND2X2_3226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4773_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4771_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__27_));
AND2X2 AND2X2_3227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4776_));
AND2X2 AND2X2_3228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4777_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4775_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__28_));
AND2X2 AND2X2_3229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4780_));
AND2X2 AND2X2_323 ( .A(_abc_44694_new_n1145_), .B(_abc_44694_new_n645_), .Y(_abc_44694_new_n1187_));
AND2X2 AND2X2_3230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4781_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4779_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__29_));
AND2X2 AND2X2_3231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4784_));
AND2X2 AND2X2_3232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4785_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4783_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__30_));
AND2X2 AND2X2_3233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4788_));
AND2X2 AND2X2_3234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4789_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4787_), .Y(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__31_));
AND2X2 AND2X2_3235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4238_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4791_));
AND2X2 AND2X2_3236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4794_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4792_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__0_));
AND2X2 AND2X2_3237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4797_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4796_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__1_));
AND2X2 AND2X2_3238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4800_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4799_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__2_));
AND2X2 AND2X2_3239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4803_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4802_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__3_));
AND2X2 AND2X2_324 ( .A(_abc_44694_new_n1188_), .B(_abc_44694_new_n1186__bF_buf3), .Y(_abc_44694_new_n1189_));
AND2X2 AND2X2_3240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4806_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4805_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__4_));
AND2X2 AND2X2_3241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4809_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4808_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__5_));
AND2X2 AND2X2_3242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4812_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4811_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__6_));
AND2X2 AND2X2_3243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4815_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4814_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__7_));
AND2X2 AND2X2_3244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4818_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4817_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__8_));
AND2X2 AND2X2_3245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4821_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4820_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__9_));
AND2X2 AND2X2_3246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4824_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4823_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__10_));
AND2X2 AND2X2_3247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4827_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4826_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__11_));
AND2X2 AND2X2_3248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4830_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4829_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__12_));
AND2X2 AND2X2_3249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4833_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4832_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__13_));
AND2X2 AND2X2_325 ( .A(_abc_44694_new_n1184_), .B(_abc_44694_new_n1189_), .Y(_abc_44694_new_n1190_));
AND2X2 AND2X2_3250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4836_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4835_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__14_));
AND2X2 AND2X2_3251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4839_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4838_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__15_));
AND2X2 AND2X2_3252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4842_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4841_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__16_));
AND2X2 AND2X2_3253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4845_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4844_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__17_));
AND2X2 AND2X2_3254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4848_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4847_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__18_));
AND2X2 AND2X2_3255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4851_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4850_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__19_));
AND2X2 AND2X2_3256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4854_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4853_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__20_));
AND2X2 AND2X2_3257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4857_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4856_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__21_));
AND2X2 AND2X2_3258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4860_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4859_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__22_));
AND2X2 AND2X2_3259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4863_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4862_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__23_));
AND2X2 AND2X2_326 ( .A(_abc_44694_new_n1190_), .B(_abc_44694_new_n1179__bF_buf3), .Y(_abc_44694_new_n1191_));
AND2X2 AND2X2_3260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4866_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4865_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__24_));
AND2X2 AND2X2_3261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4869_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4868_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__25_));
AND2X2 AND2X2_3262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4872_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4871_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__26_));
AND2X2 AND2X2_3263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4875_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4874_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__27_));
AND2X2 AND2X2_3264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4878_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4877_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__28_));
AND2X2 AND2X2_3265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4881_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4880_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__29_));
AND2X2 AND2X2_3266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4884_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4883_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__30_));
AND2X2 AND2X2_3267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4887_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4886_), .Y(REGFILE_SIM_reg_bank__0reg_r8_31_0__31_));
AND2X2 AND2X2_3268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3058_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4889_));
AND2X2 AND2X2_3269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4892_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4890_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__0_));
AND2X2 AND2X2_327 ( .A(_abc_44694_new_n1174_), .B(_abc_44694_new_n1191_), .Y(_abc_44694_new_n1192_));
AND2X2 AND2X2_3270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4895_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4894_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__1_));
AND2X2 AND2X2_3271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4898_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4897_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__2_));
AND2X2 AND2X2_3272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4901_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4900_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__3_));
AND2X2 AND2X2_3273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4904_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4903_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__4_));
AND2X2 AND2X2_3274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4907_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4906_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__5_));
AND2X2 AND2X2_3275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4910_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4909_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__6_));
AND2X2 AND2X2_3276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4913_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4912_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__7_));
AND2X2 AND2X2_3277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4916_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4915_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__8_));
AND2X2 AND2X2_3278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4919_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4918_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__9_));
AND2X2 AND2X2_3279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4922_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4921_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__10_));
AND2X2 AND2X2_328 ( .A(_abc_44694_new_n1172_), .B(_abc_44694_new_n1192_), .Y(_abc_44694_new_n1193_));
AND2X2 AND2X2_3280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4925_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4924_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__11_));
AND2X2 AND2X2_3281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4928_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4927_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__12_));
AND2X2 AND2X2_3282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4931_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4930_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__13_));
AND2X2 AND2X2_3283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4934_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4933_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__14_));
AND2X2 AND2X2_3284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4937_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4936_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__15_));
AND2X2 AND2X2_3285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4940_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4939_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__16_));
AND2X2 AND2X2_3286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4943_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4942_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__17_));
AND2X2 AND2X2_3287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4946_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4945_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__18_));
AND2X2 AND2X2_3288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4949_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4948_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__19_));
AND2X2 AND2X2_3289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4952_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4951_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__20_));
AND2X2 AND2X2_329 ( .A(_abc_44694_new_n1050_), .B(_abc_44694_new_n1021_), .Y(_abc_44694_new_n1194_));
AND2X2 AND2X2_3290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4955_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4954_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__21_));
AND2X2 AND2X2_3291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4958_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4957_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__22_));
AND2X2 AND2X2_3292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4961_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4960_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__23_));
AND2X2 AND2X2_3293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4964_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4963_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__24_));
AND2X2 AND2X2_3294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4967_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4966_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__25_));
AND2X2 AND2X2_3295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4970_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4969_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__26_));
AND2X2 AND2X2_3296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4973_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4972_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__27_));
AND2X2 AND2X2_3297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4976_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4975_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__28_));
AND2X2 AND2X2_3298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4979_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4978_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__29_));
AND2X2 AND2X2_3299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4982_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4981_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__30_));
AND2X2 AND2X2_33 ( .A(_abc_44694_new_n674_), .B(mem_offset_q_1_), .Y(_abc_44694_new_n675_));
AND2X2 AND2X2_330 ( .A(_abc_44694_new_n655_), .B(_abc_44694_new_n1194__bF_buf4), .Y(_abc_44694_new_n1195_));
AND2X2 AND2X2_3300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4985_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4984_), .Y(REGFILE_SIM_reg_bank__0reg_r7_31_0__31_));
AND2X2 AND2X2_3301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3157_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987_));
AND2X2 AND2X2_3302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4989_));
AND2X2 AND2X2_3303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4990_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4988_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__0_));
AND2X2 AND2X2_3304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4993_));
AND2X2 AND2X2_3305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4994_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4992_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__1_));
AND2X2 AND2X2_3306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4997_));
AND2X2 AND2X2_3307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4998_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n4996_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__2_));
AND2X2 AND2X2_3308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5001_));
AND2X2 AND2X2_3309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5002_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5000_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__3_));
AND2X2 AND2X2_331 ( .A(_abc_44694_new_n1169_), .B(_abc_44694_new_n1129_), .Y(_abc_44694_new_n1196_));
AND2X2 AND2X2_3310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5005_));
AND2X2 AND2X2_3311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5006_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5004_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__4_));
AND2X2 AND2X2_3312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5009_));
AND2X2 AND2X2_3313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5010_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5008_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__5_));
AND2X2 AND2X2_3314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5013_));
AND2X2 AND2X2_3315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5014_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5012_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__6_));
AND2X2 AND2X2_3316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5017_));
AND2X2 AND2X2_3317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5018_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5016_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__7_));
AND2X2 AND2X2_3318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5021_));
AND2X2 AND2X2_3319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5022_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5020_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__8_));
AND2X2 AND2X2_332 ( .A(_abc_44694_new_n1165_), .B(_abc_44694_new_n1097_), .Y(_abc_44694_new_n1197_));
AND2X2 AND2X2_3320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5025_));
AND2X2 AND2X2_3321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5026_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5024_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__9_));
AND2X2 AND2X2_3322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5029_));
AND2X2 AND2X2_3323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5030_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5028_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__10_));
AND2X2 AND2X2_3324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5033_));
AND2X2 AND2X2_3325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5034_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5032_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__11_));
AND2X2 AND2X2_3326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5037_));
AND2X2 AND2X2_3327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5038_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5036_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__12_));
AND2X2 AND2X2_3328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5041_));
AND2X2 AND2X2_3329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5042_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5040_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__13_));
AND2X2 AND2X2_333 ( .A(_abc_44694_new_n1199_), .B(_abc_44694_new_n1195_), .Y(_abc_44694_new_n1200_));
AND2X2 AND2X2_3330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5045_));
AND2X2 AND2X2_3331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5046_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5044_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__14_));
AND2X2 AND2X2_3332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5049_));
AND2X2 AND2X2_3333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5050_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5048_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__15_));
AND2X2 AND2X2_3334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5053_));
AND2X2 AND2X2_3335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5052_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__16_));
AND2X2 AND2X2_3336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5057_));
AND2X2 AND2X2_3337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5058_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5056_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__17_));
AND2X2 AND2X2_3338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5061_));
AND2X2 AND2X2_3339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5062_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5060_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__18_));
AND2X2 AND2X2_334 ( .A(_abc_44694_new_n1200_), .B(_abc_44694_new_n1193_), .Y(_abc_44694_new_n1201_));
AND2X2 AND2X2_3340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5065_));
AND2X2 AND2X2_3341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5066_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5064_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__19_));
AND2X2 AND2X2_3342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5069_));
AND2X2 AND2X2_3343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5070_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5068_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__20_));
AND2X2 AND2X2_3344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5073_));
AND2X2 AND2X2_3345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5074_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5072_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__21_));
AND2X2 AND2X2_3346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5077_));
AND2X2 AND2X2_3347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5078_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5076_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__22_));
AND2X2 AND2X2_3348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5081_));
AND2X2 AND2X2_3349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5082_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5080_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__23_));
AND2X2 AND2X2_335 ( .A(_abc_44694_new_n1201_), .B(_abc_44694_new_n1163_), .Y(_abc_44694_new_n1202_));
AND2X2 AND2X2_3350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5085_));
AND2X2 AND2X2_3351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5086_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5084_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__24_));
AND2X2 AND2X2_3352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5089_));
AND2X2 AND2X2_3353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5090_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5088_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__25_));
AND2X2 AND2X2_3354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5093_));
AND2X2 AND2X2_3355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5094_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5092_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__26_));
AND2X2 AND2X2_3356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5097_));
AND2X2 AND2X2_3357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5098_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5096_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__27_));
AND2X2 AND2X2_3358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5101_));
AND2X2 AND2X2_3359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5102_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5100_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__28_));
AND2X2 AND2X2_336 ( .A(_abc_44694_new_n1202_), .B(_abc_44694_new_n1141_), .Y(_abc_44694_new_n1203_));
AND2X2 AND2X2_3360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5105_));
AND2X2 AND2X2_3361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5106_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5104_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__29_));
AND2X2 AND2X2_3362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5109_));
AND2X2 AND2X2_3363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5110_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5108_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__30_));
AND2X2 AND2X2_3364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5113_));
AND2X2 AND2X2_3365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5114_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5112_), .Y(REGFILE_SIM_reg_bank__0reg_r6_31_0__31_));
AND2X2 AND2X2_3366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3287_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116_));
AND2X2 AND2X2_3367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5118_));
AND2X2 AND2X2_3368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5119_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5117_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__0_));
AND2X2 AND2X2_3369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5122_));
AND2X2 AND2X2_337 ( .A(_abc_44694_new_n1206_), .B(_abc_44694_new_n1050_), .Y(_abc_44694_new_n1207_));
AND2X2 AND2X2_3370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5123_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5121_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__1_));
AND2X2 AND2X2_3371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2115_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5126_));
AND2X2 AND2X2_3372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5127_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5125_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__2_));
AND2X2 AND2X2_3373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5130_));
AND2X2 AND2X2_3374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5131_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5129_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__3_));
AND2X2 AND2X2_3375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5134_));
AND2X2 AND2X2_3376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5135_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5133_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__4_));
AND2X2 AND2X2_3377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5138_));
AND2X2 AND2X2_3378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5139_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5137_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__5_));
AND2X2 AND2X2_3379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5142_));
AND2X2 AND2X2_338 ( .A(_abc_44694_new_n1207__bF_buf5), .B(_abc_44694_new_n1045_), .Y(_abc_44694_new_n1208_));
AND2X2 AND2X2_3380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5143_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5141_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__6_));
AND2X2 AND2X2_3381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5146_));
AND2X2 AND2X2_3382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5147_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5145_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__7_));
AND2X2 AND2X2_3383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5150_));
AND2X2 AND2X2_3384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5151_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5149_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__8_));
AND2X2 AND2X2_3385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5154_));
AND2X2 AND2X2_3386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5155_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5153_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__9_));
AND2X2 AND2X2_3387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5158_));
AND2X2 AND2X2_3388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5159_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5157_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__10_));
AND2X2 AND2X2_3389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5162_));
AND2X2 AND2X2_339 ( .A(_abc_44694_new_n1208_), .B(_abc_44694_new_n1043_), .Y(_abc_44694_new_n1209_));
AND2X2 AND2X2_3390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5163_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5161_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__11_));
AND2X2 AND2X2_3391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5166_));
AND2X2 AND2X2_3392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5167_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5165_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__12_));
AND2X2 AND2X2_3393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5170_));
AND2X2 AND2X2_3394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5171_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5169_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__13_));
AND2X2 AND2X2_3395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5174_));
AND2X2 AND2X2_3396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5175_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5173_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__14_));
AND2X2 AND2X2_3397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5178_));
AND2X2 AND2X2_3398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5179_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5177_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__15_));
AND2X2 AND2X2_3399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5182_));
AND2X2 AND2X2_34 ( .A(_abc_44694_new_n652_), .B(inst_r_2_), .Y(_abc_44694_new_n676_));
AND2X2 AND2X2_340 ( .A(_abc_44694_new_n1211_), .B(_abc_44694_new_n1027_), .Y(_abc_44694_new_n1212_));
AND2X2 AND2X2_3400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5183_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5181_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__16_));
AND2X2 AND2X2_3401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5186_));
AND2X2 AND2X2_3402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5187_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5185_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__17_));
AND2X2 AND2X2_3403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5190_));
AND2X2 AND2X2_3404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5191_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5189_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__18_));
AND2X2 AND2X2_3405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5194_));
AND2X2 AND2X2_3406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5195_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5193_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__19_));
AND2X2 AND2X2_3407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5198_));
AND2X2 AND2X2_3408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5199_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5197_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__20_));
AND2X2 AND2X2_3409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5202_));
AND2X2 AND2X2_341 ( .A(_abc_44694_new_n1215_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n1216_));
AND2X2 AND2X2_3410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5203_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5201_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__21_));
AND2X2 AND2X2_3411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5206_));
AND2X2 AND2X2_3412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5207_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5205_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__22_));
AND2X2 AND2X2_3413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5210_));
AND2X2 AND2X2_3414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5211_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5209_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__23_));
AND2X2 AND2X2_3415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5214_));
AND2X2 AND2X2_3416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5215_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5213_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__24_));
AND2X2 AND2X2_3417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5218_));
AND2X2 AND2X2_3418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5219_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5217_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__25_));
AND2X2 AND2X2_3419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5222_));
AND2X2 AND2X2_342 ( .A(_abc_44694_new_n1214_), .B(_abc_44694_new_n1216_), .Y(_0esr_q_31_0__2_));
AND2X2 AND2X2_3420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5223_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5221_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__26_));
AND2X2 AND2X2_3421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5226_));
AND2X2 AND2X2_3422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5225_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__27_));
AND2X2 AND2X2_3423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5230_));
AND2X2 AND2X2_3424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5231_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5229_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__28_));
AND2X2 AND2X2_3425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5234_));
AND2X2 AND2X2_3426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5235_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5233_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__29_));
AND2X2 AND2X2_3427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5238_));
AND2X2 AND2X2_3428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5239_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5237_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__30_));
AND2X2 AND2X2_3429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0), .B(REGFILE_SIM_reg_bank__abc_34819_new_n2260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5242_));
AND2X2 AND2X2_343 ( .A(_abc_44694_new_n1218_), .B(sr_q_9_), .Y(_abc_44694_new_n1219_));
AND2X2 AND2X2_3430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5243_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5241_), .Y(REGFILE_SIM_reg_bank__0reg_r5_31_0__31_));
AND2X2 AND2X2_3431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4238_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5245_));
AND2X2 AND2X2_3432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5248_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5246_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__0_));
AND2X2 AND2X2_3433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5251_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5250_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__1_));
AND2X2 AND2X2_3434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5254_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5253_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__2_));
AND2X2 AND2X2_3435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5256_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__3_));
AND2X2 AND2X2_3436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5260_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5259_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__4_));
AND2X2 AND2X2_3437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5263_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5262_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__5_));
AND2X2 AND2X2_3438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5266_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5265_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__6_));
AND2X2 AND2X2_3439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5269_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5268_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__7_));
AND2X2 AND2X2_344 ( .A(_abc_44694_new_n1169_), .B(_abc_44694_new_n1105_), .Y(_abc_44694_new_n1220_));
AND2X2 AND2X2_3440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5272_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5271_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__8_));
AND2X2 AND2X2_3441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5275_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5274_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__9_));
AND2X2 AND2X2_3442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5278_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5277_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__10_));
AND2X2 AND2X2_3443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5281_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5280_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__11_));
AND2X2 AND2X2_3444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5284_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5283_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__12_));
AND2X2 AND2X2_3445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5287_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5286_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__13_));
AND2X2 AND2X2_3446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5290_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5289_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__14_));
AND2X2 AND2X2_3447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5293_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5292_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__15_));
AND2X2 AND2X2_3448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5296_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5295_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__16_));
AND2X2 AND2X2_3449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5299_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5298_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__17_));
AND2X2 AND2X2_345 ( .A(_abc_44694_new_n1196_), .B(alu_equal_o), .Y(_abc_44694_new_n1222_));
AND2X2 AND2X2_3450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5302_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5301_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__18_));
AND2X2 AND2X2_3451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5305_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5304_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__19_));
AND2X2 AND2X2_3452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5308_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5307_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__20_));
AND2X2 AND2X2_3453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5311_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5310_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__21_));
AND2X2 AND2X2_3454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5314_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5313_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__22_));
AND2X2 AND2X2_3455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5317_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5316_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__23_));
AND2X2 AND2X2_3456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5320_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5319_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__24_));
AND2X2 AND2X2_3457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5323_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5322_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__25_));
AND2X2 AND2X2_3458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5326_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5325_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__26_));
AND2X2 AND2X2_3459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5329_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5328_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__27_));
AND2X2 AND2X2_346 ( .A(_abc_44694_new_n1223_), .B(_abc_44694_new_n1221_), .Y(_abc_44694_new_n1224_));
AND2X2 AND2X2_3460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5332_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5331_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__28_));
AND2X2 AND2X2_3461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5335_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5334_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__29_));
AND2X2 AND2X2_3462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5338_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5337_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__30_));
AND2X2 AND2X2_3463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5341_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5340_), .Y(REGFILE_SIM_reg_bank__0reg_r4_31_0__31_));
AND2X2 AND2X2_3464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3516_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5343_));
AND2X2 AND2X2_3465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5346_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5344_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__0_));
AND2X2 AND2X2_3466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5349_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5348_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__1_));
AND2X2 AND2X2_3467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5352_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5351_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__2_));
AND2X2 AND2X2_3468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5355_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5354_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__3_));
AND2X2 AND2X2_3469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5358_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5357_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__4_));
AND2X2 AND2X2_347 ( .A(_abc_44694_new_n1225_), .B(_abc_44694_new_n1227_), .Y(_abc_44694_new_n1228_));
AND2X2 AND2X2_3470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5361_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5360_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__5_));
AND2X2 AND2X2_3471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5364_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5363_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__6_));
AND2X2 AND2X2_3472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5366_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__7_));
AND2X2 AND2X2_3473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5370_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5369_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__8_));
AND2X2 AND2X2_3474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5373_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5372_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__9_));
AND2X2 AND2X2_3475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5376_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5375_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__10_));
AND2X2 AND2X2_3476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5379_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5378_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__11_));
AND2X2 AND2X2_3477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5382_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5381_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__12_));
AND2X2 AND2X2_3478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5385_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5384_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__13_));
AND2X2 AND2X2_3479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5388_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5387_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__14_));
AND2X2 AND2X2_348 ( .A(_abc_44694_new_n1197_), .B(_abc_44694_new_n1230_), .Y(_abc_44694_new_n1231_));
AND2X2 AND2X2_3480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5391_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5390_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__15_));
AND2X2 AND2X2_3481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5394_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5393_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__16_));
AND2X2 AND2X2_3482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5397_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5396_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__17_));
AND2X2 AND2X2_3483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5400_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5399_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__18_));
AND2X2 AND2X2_3484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5403_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5402_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__19_));
AND2X2 AND2X2_3485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5406_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5405_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__20_));
AND2X2 AND2X2_3486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5409_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5408_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__21_));
AND2X2 AND2X2_3487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5412_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5411_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__22_));
AND2X2 AND2X2_3488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5415_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5414_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__23_));
AND2X2 AND2X2_3489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5418_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5417_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__24_));
AND2X2 AND2X2_349 ( .A(_abc_44694_new_n1232_), .B(_abc_44694_new_n1133_), .Y(_abc_44694_new_n1233_));
AND2X2 AND2X2_3490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5421_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5420_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__25_));
AND2X2 AND2X2_3491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5424_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5423_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__26_));
AND2X2 AND2X2_3492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5427_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5426_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__27_));
AND2X2 AND2X2_3493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5430_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5429_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__28_));
AND2X2 AND2X2_3494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5433_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5432_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__29_));
AND2X2 AND2X2_3495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5436_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5435_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__30_));
AND2X2 AND2X2_3496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5439_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5438_), .Y(REGFILE_SIM_reg_bank__0reg_r3_31_0__31_));
AND2X2 AND2X2_3497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3615_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n3912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5441_));
AND2X2 AND2X2_3498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5444_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5442_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__0_));
AND2X2 AND2X2_3499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5447_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5446_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__1_));
AND2X2 AND2X2_35 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[0] ), .Y(_abc_44694_new_n679_));
AND2X2 AND2X2_350 ( .A(_abc_44694_new_n1229_), .B(_abc_44694_new_n1233_), .Y(_abc_44694_new_n1234_));
AND2X2 AND2X2_3500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5450_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5449_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__2_));
AND2X2 AND2X2_3501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5453_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5452_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__3_));
AND2X2 AND2X2_3502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5456_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5455_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__4_));
AND2X2 AND2X2_3503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5459_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5458_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__5_));
AND2X2 AND2X2_3504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5462_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5461_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__6_));
AND2X2 AND2X2_3505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5465_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5464_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__7_));
AND2X2 AND2X2_3506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5468_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5467_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__8_));
AND2X2 AND2X2_3507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5470_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__9_));
AND2X2 AND2X2_3508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5474_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5473_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__10_));
AND2X2 AND2X2_3509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5477_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5476_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__11_));
AND2X2 AND2X2_351 ( .A(_abc_44694_new_n1132_), .B(_abc_44694_new_n1235_), .Y(_abc_44694_new_n1236_));
AND2X2 AND2X2_3510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5480_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5479_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__12_));
AND2X2 AND2X2_3511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5483_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5482_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__13_));
AND2X2 AND2X2_3512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5486_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5485_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__14_));
AND2X2 AND2X2_3513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5489_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5488_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__15_));
AND2X2 AND2X2_3514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5492_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5491_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__16_));
AND2X2 AND2X2_3515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5494_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__17_));
AND2X2 AND2X2_3516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5498_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5497_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__18_));
AND2X2 AND2X2_3517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5501_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5500_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__19_));
AND2X2 AND2X2_3518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5504_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5503_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__20_));
AND2X2 AND2X2_3519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5507_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5506_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__21_));
AND2X2 AND2X2_352 ( .A(_abc_44694_new_n1239_), .B(_abc_44694_new_n1230_), .Y(_abc_44694_new_n1240_));
AND2X2 AND2X2_3520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5510_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5509_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__22_));
AND2X2 AND2X2_3521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5513_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5512_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__23_));
AND2X2 AND2X2_3522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5516_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5515_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__24_));
AND2X2 AND2X2_3523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5519_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5518_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__25_));
AND2X2 AND2X2_3524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5522_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5521_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__26_));
AND2X2 AND2X2_3525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5525_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5524_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__27_));
AND2X2 AND2X2_3526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5528_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5527_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__28_));
AND2X2 AND2X2_3527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5531_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5530_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__29_));
AND2X2 AND2X2_3528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5534_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5533_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__30_));
AND2X2 AND2X2_3529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5537_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5536_), .Y(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__31_));
AND2X2 AND2X2_353 ( .A(_abc_44694_new_n1166_), .B(_abc_44694_new_n1240_), .Y(_abc_44694_new_n1241_));
AND2X2 AND2X2_3530 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5540_));
AND2X2 AND2X2_3531 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5541_));
AND2X2 AND2X2_3532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5540_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5542_));
AND2X2 AND2X2_3533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5542_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5543_));
AND2X2 AND2X2_3534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5544_));
AND2X2 AND2X2_3535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5545_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5546_));
AND2X2 AND2X2_3536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5546_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5547_));
AND2X2 AND2X2_3537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5547_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5548_));
AND2X2 AND2X2_3538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5549_));
AND2X2 AND2X2_3539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5551_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5545_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5552_));
AND2X2 AND2X2_354 ( .A(_abc_44694_new_n1238_), .B(_abc_44694_new_n1242_), .Y(_abc_44694_new_n1243_));
AND2X2 AND2X2_3540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5552_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5553_));
AND2X2 AND2X2_3541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5553_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5554_));
AND2X2 AND2X2_3542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5555_));
AND2X2 AND2X2_3543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5551_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5556_));
AND2X2 AND2X2_3544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5557_));
AND2X2 AND2X2_3545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5557_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5558_));
AND2X2 AND2X2_3546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5559_));
AND2X2 AND2X2_3547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5562_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5563_));
AND2X2 AND2X2_3548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5546_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5564_));
AND2X2 AND2X2_3549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5564_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5565_));
AND2X2 AND2X2_355 ( .A(_abc_44694_new_n1220_), .B(_abc_44694_new_n1246_), .Y(_abc_44694_new_n1247_));
AND2X2 AND2X2_3550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5566_));
AND2X2 AND2X2_3551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5540_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5567_));
AND2X2 AND2X2_3552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5567_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5568_));
AND2X2 AND2X2_3553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5569_));
AND2X2 AND2X2_3554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5563_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5571_));
AND2X2 AND2X2_3555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5571_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5572_));
AND2X2 AND2X2_3556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5573_));
AND2X2 AND2X2_3557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5553_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5563_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5574_));
AND2X2 AND2X2_3558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5575_));
AND2X2 AND2X2_3559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5579_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5562_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5580_));
AND2X2 AND2X2_356 ( .A(_abc_44694_new_n1248_), .B(_abc_44694_new_n1245_), .Y(_abc_44694_new_n1249_));
AND2X2 AND2X2_3560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5580_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5556_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5581_));
AND2X2 AND2X2_3561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5581_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5582_));
AND2X2 AND2X2_3562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5583_));
AND2X2 AND2X2_3563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5580_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5546_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5584_));
AND2X2 AND2X2_3564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5584_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5585_));
AND2X2 AND2X2_3565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5586_));
AND2X2 AND2X2_3566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5580_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5540_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5587_));
AND2X2 AND2X2_3567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5587_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5588_));
AND2X2 AND2X2_3568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5589_));
AND2X2 AND2X2_3569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5579_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5592_));
AND2X2 AND2X2_357 ( .A(_abc_44694_new_n1244_), .B(_abc_44694_new_n1249_), .Y(_abc_44694_new_n1250_));
AND2X2 AND2X2_3570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5593_));
AND2X2 AND2X2_3571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5593_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5594_));
AND2X2 AND2X2_3572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5595_));
AND2X2 AND2X2_3573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5553_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5596_));
AND2X2 AND2X2_3574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5597_));
AND2X2 AND2X2_3575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5592_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5540_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5599_));
AND2X2 AND2X2_3576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5599_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5600_));
AND2X2 AND2X2_3577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5601_));
AND2X2 AND2X2_3578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5546_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5602_));
AND2X2 AND2X2_3579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5602_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5603_));
AND2X2 AND2X2_358 ( .A(_abc_44694_new_n1110_), .B(alu_greater_than_signed_o), .Y(_abc_44694_new_n1251_));
AND2X2 AND2X2_3580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5604_));
AND2X2 AND2X2_3581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5542_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5609_));
AND2X2 AND2X2_3582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5610_));
AND2X2 AND2X2_3583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5547_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5611_));
AND2X2 AND2X2_3584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5612_));
AND2X2 AND2X2_3585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5552_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5614_));
AND2X2 AND2X2_3586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5614_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5615_));
AND2X2 AND2X2_3587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5616_));
AND2X2 AND2X2_3588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5557_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5617_));
AND2X2 AND2X2_3589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5618_));
AND2X2 AND2X2_359 ( .A(_abc_44694_new_n1255_), .B(_abc_44694_new_n1137_), .Y(_abc_44694_new_n1256_));
AND2X2 AND2X2_3590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5571_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5621_));
AND2X2 AND2X2_3591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5622_));
AND2X2 AND2X2_3592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5614_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5563_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5623_));
AND2X2 AND2X2_3593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5624_));
AND2X2 AND2X2_3594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5564_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5626_));
AND2X2 AND2X2_3595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5627_));
AND2X2 AND2X2_3596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5567_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5628_));
AND2X2 AND2X2_3597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5629_));
AND2X2 AND2X2_3598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5581_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5633_));
AND2X2 AND2X2_3599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5634_));
AND2X2 AND2X2_36 ( .A(_abc_44694_new_n680_), .B(_abc_44694_new_n674_), .Y(_abc_44694_new_n681_));
AND2X2 AND2X2_360 ( .A(_abc_44694_new_n1253_), .B(_abc_44694_new_n1256_), .Y(_abc_44694_new_n1257_));
AND2X2 AND2X2_3600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5614_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5580_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5635_));
AND2X2 AND2X2_3601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5636_));
AND2X2 AND2X2_3602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5584_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5638_));
AND2X2 AND2X2_3603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5639_));
AND2X2 AND2X2_3604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5587_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5640_));
AND2X2 AND2X2_3605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5641_));
AND2X2 AND2X2_3606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5614_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5644_));
AND2X2 AND2X2_3607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5645_));
AND2X2 AND2X2_3608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5593_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5646_));
AND2X2 AND2X2_3609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5647_));
AND2X2 AND2X2_361 ( .A(_abc_44694_new_n1136_), .B(_abc_44694_new_n1258_), .Y(_abc_44694_new_n1259_));
AND2X2 AND2X2_3610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5602_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5649_));
AND2X2 AND2X2_3611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5650_));
AND2X2 AND2X2_3612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5599_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5651_));
AND2X2 AND2X2_3613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5652_));
AND2X2 AND2X2_3614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5658_));
AND2X2 AND2X2_3615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5659_));
AND2X2 AND2X2_3616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5661_));
AND2X2 AND2X2_3617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5662_));
AND2X2 AND2X2_3618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5665_));
AND2X2 AND2X2_3619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5666_));
AND2X2 AND2X2_362 ( .A(_abc_44694_new_n1260_), .B(alu_flag_update_o), .Y(_abc_44694_new_n1261_));
AND2X2 AND2X2_3620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5668_));
AND2X2 AND2X2_3621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5669_));
AND2X2 AND2X2_3622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5673_));
AND2X2 AND2X2_3623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5674_));
AND2X2 AND2X2_3624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5675_));
AND2X2 AND2X2_3625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5678_));
AND2X2 AND2X2_3626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5679_));
AND2X2 AND2X2_3627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5681_));
AND2X2 AND2X2_3628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5682_));
AND2X2 AND2X2_3629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5687_));
AND2X2 AND2X2_363 ( .A(_abc_44694_new_n1262_), .B(_abc_44694_new_n1088_), .Y(_abc_44694_new_n1263_));
AND2X2 AND2X2_3630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5688_));
AND2X2 AND2X2_3631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5690_));
AND2X2 AND2X2_3632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5691_));
AND2X2 AND2X2_3633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5694_));
AND2X2 AND2X2_3634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5695_));
AND2X2 AND2X2_3635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5697_));
AND2X2 AND2X2_3636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5698_));
AND2X2 AND2X2_3637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5702_));
AND2X2 AND2X2_3638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5703_));
AND2X2 AND2X2_3639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5705_));
AND2X2 AND2X2_364 ( .A(_abc_44694_new_n1260_), .B(_abc_44694_new_n1089_), .Y(_abc_44694_new_n1264_));
AND2X2 AND2X2_3640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5706_));
AND2X2 AND2X2_3641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5709_));
AND2X2 AND2X2_3642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5710_));
AND2X2 AND2X2_3643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5712_));
AND2X2 AND2X2_3644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5713_));
AND2X2 AND2X2_3645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5719_));
AND2X2 AND2X2_3646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5720_));
AND2X2 AND2X2_3647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5722_));
AND2X2 AND2X2_3648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5723_));
AND2X2 AND2X2_3649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5726_));
AND2X2 AND2X2_365 ( .A(_abc_44694_new_n1267_), .B(_abc_44694_new_n1017_), .Y(_abc_44694_new_n1268_));
AND2X2 AND2X2_3650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5727_));
AND2X2 AND2X2_3651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5729_));
AND2X2 AND2X2_3652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5730_));
AND2X2 AND2X2_3653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5734_));
AND2X2 AND2X2_3654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5735_));
AND2X2 AND2X2_3655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5736_));
AND2X2 AND2X2_3656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5739_));
AND2X2 AND2X2_3657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5740_));
AND2X2 AND2X2_3658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5742_));
AND2X2 AND2X2_3659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5743_));
AND2X2 AND2X2_366 ( .A(_abc_44694_new_n1266_), .B(_abc_44694_new_n1268_), .Y(_abc_44694_new_n1269_));
AND2X2 AND2X2_3660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5748_));
AND2X2 AND2X2_3661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5749_));
AND2X2 AND2X2_3662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5751_));
AND2X2 AND2X2_3663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5752_));
AND2X2 AND2X2_3664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5755_));
AND2X2 AND2X2_3665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5756_));
AND2X2 AND2X2_3666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5758_));
AND2X2 AND2X2_3667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5759_));
AND2X2 AND2X2_3668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5763_));
AND2X2 AND2X2_3669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5764_));
AND2X2 AND2X2_367 ( .A(_abc_44694_new_n1011_), .B(_abc_44694_new_n1271_), .Y(_abc_44694_new_n1272_));
AND2X2 AND2X2_3670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5766_));
AND2X2 AND2X2_3671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5767_));
AND2X2 AND2X2_3672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5770_));
AND2X2 AND2X2_3673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5771_));
AND2X2 AND2X2_3674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5773_));
AND2X2 AND2X2_3675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5774_));
AND2X2 AND2X2_3676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5780_));
AND2X2 AND2X2_3677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5781_));
AND2X2 AND2X2_3678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5783_));
AND2X2 AND2X2_3679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5784_));
AND2X2 AND2X2_368 ( .A(_abc_44694_new_n1273_), .B(_abc_44694_new_n970_), .Y(_abc_44694_new_n1274_));
AND2X2 AND2X2_3680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5787_));
AND2X2 AND2X2_3681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5788_));
AND2X2 AND2X2_3682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5790_));
AND2X2 AND2X2_3683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5791_));
AND2X2 AND2X2_3684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5795_));
AND2X2 AND2X2_3685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5796_));
AND2X2 AND2X2_3686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5797_));
AND2X2 AND2X2_3687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5800_));
AND2X2 AND2X2_3688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5801_));
AND2X2 AND2X2_3689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5803_));
AND2X2 AND2X2_369 ( .A(_abc_44694_new_n1270_), .B(_abc_44694_new_n1274_), .Y(_abc_44694_new_n1275_));
AND2X2 AND2X2_3690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5804_));
AND2X2 AND2X2_3691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5809_));
AND2X2 AND2X2_3692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5810_));
AND2X2 AND2X2_3693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5812_));
AND2X2 AND2X2_3694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5813_));
AND2X2 AND2X2_3695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5816_));
AND2X2 AND2X2_3696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5817_));
AND2X2 AND2X2_3697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5819_));
AND2X2 AND2X2_3698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5820_));
AND2X2 AND2X2_3699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5824_));
AND2X2 AND2X2_37 ( .A(_abc_44694_new_n676_), .B(_abc_44694_new_n681_), .Y(_abc_44694_new_n682_));
AND2X2 AND2X2_370 ( .A(_abc_44694_new_n1277_), .B(_abc_44694_new_n1045_), .Y(_abc_44694_new_n1278_));
AND2X2 AND2X2_3700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5825_));
AND2X2 AND2X2_3701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5827_));
AND2X2 AND2X2_3702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5828_));
AND2X2 AND2X2_3703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5831_));
AND2X2 AND2X2_3704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5832_));
AND2X2 AND2X2_3705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5834_));
AND2X2 AND2X2_3706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5835_));
AND2X2 AND2X2_3707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5841_));
AND2X2 AND2X2_3708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5842_));
AND2X2 AND2X2_3709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5844_));
AND2X2 AND2X2_371 ( .A(_abc_44694_new_n1207__bF_buf4), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n1279_));
AND2X2 AND2X2_3710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5845_));
AND2X2 AND2X2_3711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5848_));
AND2X2 AND2X2_3712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5849_));
AND2X2 AND2X2_3713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5851_));
AND2X2 AND2X2_3714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5852_));
AND2X2 AND2X2_3715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5856_));
AND2X2 AND2X2_3716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5857_));
AND2X2 AND2X2_3717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5858_));
AND2X2 AND2X2_3718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5861_));
AND2X2 AND2X2_3719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5862_));
AND2X2 AND2X2_372 ( .A(_abc_44694_new_n1276_), .B(_abc_44694_new_n1280_), .Y(_abc_44694_new_n1281_));
AND2X2 AND2X2_3720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5864_));
AND2X2 AND2X2_3721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5865_));
AND2X2 AND2X2_3722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5870_));
AND2X2 AND2X2_3723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5871_));
AND2X2 AND2X2_3724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5873_));
AND2X2 AND2X2_3725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5874_));
AND2X2 AND2X2_3726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5877_));
AND2X2 AND2X2_3727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5878_));
AND2X2 AND2X2_3728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5880_));
AND2X2 AND2X2_3729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5881_));
AND2X2 AND2X2_373 ( .A(_abc_44694_new_n1039_), .B(esr_q_9_), .Y(_abc_44694_new_n1282_));
AND2X2 AND2X2_3730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5885_));
AND2X2 AND2X2_3731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5886_));
AND2X2 AND2X2_3732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5888_));
AND2X2 AND2X2_3733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5889_));
AND2X2 AND2X2_3734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5892_));
AND2X2 AND2X2_3735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5893_));
AND2X2 AND2X2_3736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5895_));
AND2X2 AND2X2_3737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5896_));
AND2X2 AND2X2_3738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5902_));
AND2X2 AND2X2_3739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5903_));
AND2X2 AND2X2_374 ( .A(_abc_44694_new_n1038_), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n1283_));
AND2X2 AND2X2_3740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5905_));
AND2X2 AND2X2_3741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5906_));
AND2X2 AND2X2_3742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5909_));
AND2X2 AND2X2_3743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5910_));
AND2X2 AND2X2_3744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5912_));
AND2X2 AND2X2_3745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5913_));
AND2X2 AND2X2_3746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5917_));
AND2X2 AND2X2_3747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5918_));
AND2X2 AND2X2_3748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5919_));
AND2X2 AND2X2_3749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5922_));
AND2X2 AND2X2_375 ( .A(_abc_44694_new_n1279_), .B(_abc_44694_new_n1284_), .Y(_abc_44694_new_n1285_));
AND2X2 AND2X2_3750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5923_));
AND2X2 AND2X2_3751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5925_));
AND2X2 AND2X2_3752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5926_));
AND2X2 AND2X2_3753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5931_));
AND2X2 AND2X2_3754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5932_));
AND2X2 AND2X2_3755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5934_));
AND2X2 AND2X2_3756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5935_));
AND2X2 AND2X2_3757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5938_));
AND2X2 AND2X2_3758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5939_));
AND2X2 AND2X2_3759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5941_));
AND2X2 AND2X2_376 ( .A(_abc_44694_new_n1288_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n1289_));
AND2X2 AND2X2_3760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5942_));
AND2X2 AND2X2_3761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5946_));
AND2X2 AND2X2_3762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5947_));
AND2X2 AND2X2_3763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5949_));
AND2X2 AND2X2_3764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5950_));
AND2X2 AND2X2_3765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5953_));
AND2X2 AND2X2_3766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5954_));
AND2X2 AND2X2_3767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5956_));
AND2X2 AND2X2_3768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5957_));
AND2X2 AND2X2_3769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5963_));
AND2X2 AND2X2_377 ( .A(_abc_44694_new_n1287_), .B(_abc_44694_new_n1289_), .Y(_0esr_q_31_0__9_));
AND2X2 AND2X2_3770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5964_));
AND2X2 AND2X2_3771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5966_));
AND2X2 AND2X2_3772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5967_));
AND2X2 AND2X2_3773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5970_));
AND2X2 AND2X2_3774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5971_));
AND2X2 AND2X2_3775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5973_));
AND2X2 AND2X2_3776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5974_));
AND2X2 AND2X2_3777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5978_));
AND2X2 AND2X2_3778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5979_));
AND2X2 AND2X2_3779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5980_));
AND2X2 AND2X2_378 ( .A(_abc_44694_new_n1039_), .B(esr_q_10_), .Y(_abc_44694_new_n1291_));
AND2X2 AND2X2_3780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5983_));
AND2X2 AND2X2_3781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5984_));
AND2X2 AND2X2_3782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5986_));
AND2X2 AND2X2_3783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5987_));
AND2X2 AND2X2_3784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5992_));
AND2X2 AND2X2_3785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5993_));
AND2X2 AND2X2_3786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5995_));
AND2X2 AND2X2_3787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5996_));
AND2X2 AND2X2_3788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5999_));
AND2X2 AND2X2_3789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6000_));
AND2X2 AND2X2_379 ( .A(_abc_44694_new_n1038_), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n1292_));
AND2X2 AND2X2_3790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6002_));
AND2X2 AND2X2_3791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6003_));
AND2X2 AND2X2_3792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6007_));
AND2X2 AND2X2_3793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6008_));
AND2X2 AND2X2_3794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6010_));
AND2X2 AND2X2_3795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6011_));
AND2X2 AND2X2_3796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6014_));
AND2X2 AND2X2_3797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6015_));
AND2X2 AND2X2_3798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6017_));
AND2X2 AND2X2_3799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6018_));
AND2X2 AND2X2_38 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[16] ), .Y(_abc_44694_new_n683_));
AND2X2 AND2X2_380 ( .A(_abc_44694_new_n1279_), .B(_abc_44694_new_n1293_), .Y(_abc_44694_new_n1294_));
AND2X2 AND2X2_3800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6024_));
AND2X2 AND2X2_3801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6025_));
AND2X2 AND2X2_3802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6027_));
AND2X2 AND2X2_3803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6028_));
AND2X2 AND2X2_3804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6031_));
AND2X2 AND2X2_3805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6032_));
AND2X2 AND2X2_3806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6034_));
AND2X2 AND2X2_3807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6035_));
AND2X2 AND2X2_3808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6039_));
AND2X2 AND2X2_3809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6040_));
AND2X2 AND2X2_381 ( .A(_abc_44694_new_n1297_), .B(_abc_44694_new_n1295_), .Y(_abc_44694_new_n1298_));
AND2X2 AND2X2_3810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6041_));
AND2X2 AND2X2_3811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6044_));
AND2X2 AND2X2_3812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6045_));
AND2X2 AND2X2_3813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6047_));
AND2X2 AND2X2_3814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6048_));
AND2X2 AND2X2_3815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6053_));
AND2X2 AND2X2_3816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6054_));
AND2X2 AND2X2_3817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6056_));
AND2X2 AND2X2_3818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6057_));
AND2X2 AND2X2_3819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6060_));
AND2X2 AND2X2_382 ( .A(_abc_44694_new_n1300_), .B(_abc_44694_new_n1299_), .Y(_abc_44694_new_n1301_));
AND2X2 AND2X2_3820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6061_));
AND2X2 AND2X2_3821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6063_));
AND2X2 AND2X2_3822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6064_));
AND2X2 AND2X2_3823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6068_));
AND2X2 AND2X2_3824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6069_));
AND2X2 AND2X2_3825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6071_));
AND2X2 AND2X2_3826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6072_));
AND2X2 AND2X2_3827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6075_));
AND2X2 AND2X2_3828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6076_));
AND2X2 AND2X2_3829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6078_));
AND2X2 AND2X2_383 ( .A(_abc_44694_new_n1011_), .B(_abc_44694_new_n1304_), .Y(_abc_44694_new_n1305_));
AND2X2 AND2X2_3830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6079_));
AND2X2 AND2X2_3831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6085_));
AND2X2 AND2X2_3832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6086_));
AND2X2 AND2X2_3833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6088_));
AND2X2 AND2X2_3834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6089_));
AND2X2 AND2X2_3835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6092_));
AND2X2 AND2X2_3836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6093_));
AND2X2 AND2X2_3837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6095_));
AND2X2 AND2X2_3838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6096_));
AND2X2 AND2X2_3839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6100_));
AND2X2 AND2X2_384 ( .A(_abc_44694_new_n1306_), .B(_abc_44694_new_n1303_), .Y(_abc_44694_new_n1307_));
AND2X2 AND2X2_3840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6101_));
AND2X2 AND2X2_3841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6102_));
AND2X2 AND2X2_3842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6105_));
AND2X2 AND2X2_3843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6106_));
AND2X2 AND2X2_3844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6108_));
AND2X2 AND2X2_3845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6109_));
AND2X2 AND2X2_3846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6114_));
AND2X2 AND2X2_3847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6115_));
AND2X2 AND2X2_3848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6117_));
AND2X2 AND2X2_3849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6118_));
AND2X2 AND2X2_385 ( .A(_abc_44694_new_n1308_), .B(_abc_44694_new_n1302_), .Y(_abc_44694_new_n1309_));
AND2X2 AND2X2_3850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6121_));
AND2X2 AND2X2_3851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6122_));
AND2X2 AND2X2_3852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6124_));
AND2X2 AND2X2_3853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6125_));
AND2X2 AND2X2_3854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6129_));
AND2X2 AND2X2_3855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6130_));
AND2X2 AND2X2_3856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6132_));
AND2X2 AND2X2_3857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6133_));
AND2X2 AND2X2_3858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6136_));
AND2X2 AND2X2_3859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6137_));
AND2X2 AND2X2_386 ( .A(_abc_44694_new_n1280_), .B(_abc_44694_new_n1309_), .Y(_abc_44694_new_n1310_));
AND2X2 AND2X2_3860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6139_));
AND2X2 AND2X2_3861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6140_));
AND2X2 AND2X2_3862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6146_));
AND2X2 AND2X2_3863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6147_));
AND2X2 AND2X2_3864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6149_));
AND2X2 AND2X2_3865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6150_));
AND2X2 AND2X2_3866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6153_));
AND2X2 AND2X2_3867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6154_));
AND2X2 AND2X2_3868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6156_));
AND2X2 AND2X2_3869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6157_));
AND2X2 AND2X2_387 ( .A(_abc_44694_new_n1313_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n1314_));
AND2X2 AND2X2_3870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6161_));
AND2X2 AND2X2_3871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6162_));
AND2X2 AND2X2_3872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6163_));
AND2X2 AND2X2_3873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6166_));
AND2X2 AND2X2_3874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6167_));
AND2X2 AND2X2_3875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6169_));
AND2X2 AND2X2_3876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6170_));
AND2X2 AND2X2_3877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6175_));
AND2X2 AND2X2_3878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6176_));
AND2X2 AND2X2_3879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6178_));
AND2X2 AND2X2_388 ( .A(_abc_44694_new_n1312_), .B(_abc_44694_new_n1314_), .Y(_0esr_q_31_0__10_));
AND2X2 AND2X2_3880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6179_));
AND2X2 AND2X2_3881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6182_));
AND2X2 AND2X2_3882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6183_));
AND2X2 AND2X2_3883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6185_));
AND2X2 AND2X2_3884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6186_));
AND2X2 AND2X2_3885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6190_));
AND2X2 AND2X2_3886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6191_));
AND2X2 AND2X2_3887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6193_));
AND2X2 AND2X2_3888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6194_));
AND2X2 AND2X2_3889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6197_));
AND2X2 AND2X2_389 ( .A(_abc_44694_new_n1027_), .B(_abc_44694_new_n1316_), .Y(_abc_44694_new_n1317_));
AND2X2 AND2X2_3890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6198_));
AND2X2 AND2X2_3891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6200_));
AND2X2 AND2X2_3892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6201_));
AND2X2 AND2X2_3893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6207_));
AND2X2 AND2X2_3894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6208_));
AND2X2 AND2X2_3895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6210_));
AND2X2 AND2X2_3896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6211_));
AND2X2 AND2X2_3897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6214_));
AND2X2 AND2X2_3898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6215_));
AND2X2 AND2X2_3899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6217_));
AND2X2 AND2X2_39 ( .A(_abc_44694_new_n684_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n685_));
AND2X2 AND2X2_390 ( .A(_abc_44694_new_n1208_), .B(_abc_44694_new_n1317_), .Y(_abc_44694_new_n1318_));
AND2X2 AND2X2_3900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6218_));
AND2X2 AND2X2_3901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6222_));
AND2X2 AND2X2_3902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6223_));
AND2X2 AND2X2_3903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6224_));
AND2X2 AND2X2_3904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6227_));
AND2X2 AND2X2_3905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6228_));
AND2X2 AND2X2_3906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6230_));
AND2X2 AND2X2_3907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6231_));
AND2X2 AND2X2_3908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6236_));
AND2X2 AND2X2_3909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6237_));
AND2X2 AND2X2_391 ( .A(_abc_44694_new_n1320_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n1321_));
AND2X2 AND2X2_3910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6239_));
AND2X2 AND2X2_3911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6240_));
AND2X2 AND2X2_3912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6243_));
AND2X2 AND2X2_3913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6244_));
AND2X2 AND2X2_3914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6246_));
AND2X2 AND2X2_3915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6247_));
AND2X2 AND2X2_3916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6251_));
AND2X2 AND2X2_3917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6252_));
AND2X2 AND2X2_3918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6254_));
AND2X2 AND2X2_3919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6255_));
AND2X2 AND2X2_392 ( .A(_abc_44694_new_n1319_), .B(_abc_44694_new_n1321_), .Y(_0sr_q_31_0__2_));
AND2X2 AND2X2_3920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6258_));
AND2X2 AND2X2_3921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6259_));
AND2X2 AND2X2_3922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6261_));
AND2X2 AND2X2_3923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6262_));
AND2X2 AND2X2_3924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6268_));
AND2X2 AND2X2_3925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6269_));
AND2X2 AND2X2_3926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6271_));
AND2X2 AND2X2_3927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6272_));
AND2X2 AND2X2_3928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6275_));
AND2X2 AND2X2_3929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6276_));
AND2X2 AND2X2_393 ( .A(_abc_44694_new_n1276_), .B(_abc_44694_new_n1279_), .Y(_abc_44694_new_n1323_));
AND2X2 AND2X2_3930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6278_));
AND2X2 AND2X2_3931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6279_));
AND2X2 AND2X2_3932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6283_));
AND2X2 AND2X2_3933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6284_));
AND2X2 AND2X2_3934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6285_));
AND2X2 AND2X2_3935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6288_));
AND2X2 AND2X2_3936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6289_));
AND2X2 AND2X2_3937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6291_));
AND2X2 AND2X2_3938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6292_));
AND2X2 AND2X2_3939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6297_));
AND2X2 AND2X2_394 ( .A(_abc_44694_new_n1325_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n1326_));
AND2X2 AND2X2_3940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6298_));
AND2X2 AND2X2_3941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6300_));
AND2X2 AND2X2_3942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6301_));
AND2X2 AND2X2_3943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6304_));
AND2X2 AND2X2_3944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6305_));
AND2X2 AND2X2_3945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6307_));
AND2X2 AND2X2_3946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6308_));
AND2X2 AND2X2_3947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6312_));
AND2X2 AND2X2_3948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6313_));
AND2X2 AND2X2_3949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6315_));
AND2X2 AND2X2_395 ( .A(_abc_44694_new_n1324_), .B(_abc_44694_new_n1326_), .Y(_0sr_q_31_0__9_));
AND2X2 AND2X2_3950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6316_));
AND2X2 AND2X2_3951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6319_));
AND2X2 AND2X2_3952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6320_));
AND2X2 AND2X2_3953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6322_));
AND2X2 AND2X2_3954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6323_));
AND2X2 AND2X2_3955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6329_));
AND2X2 AND2X2_3956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6330_));
AND2X2 AND2X2_3957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6332_));
AND2X2 AND2X2_3958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6333_));
AND2X2 AND2X2_3959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6336_));
AND2X2 AND2X2_396 ( .A(_abc_44694_new_n1210__bF_buf2), .B(alu_c_i), .Y(_abc_44694_new_n1328_));
AND2X2 AND2X2_3960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6337_));
AND2X2 AND2X2_3961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6339_));
AND2X2 AND2X2_3962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6340_));
AND2X2 AND2X2_3963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6344_));
AND2X2 AND2X2_3964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6345_));
AND2X2 AND2X2_3965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6346_));
AND2X2 AND2X2_3966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6349_));
AND2X2 AND2X2_3967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6350_));
AND2X2 AND2X2_3968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6352_));
AND2X2 AND2X2_3969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6353_));
AND2X2 AND2X2_397 ( .A(_abc_44694_new_n1278__bF_buf4), .B(_abc_44694_new_n1309_), .Y(_abc_44694_new_n1329_));
AND2X2 AND2X2_3970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6358_));
AND2X2 AND2X2_3971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6359_));
AND2X2 AND2X2_3972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6361_));
AND2X2 AND2X2_3973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6362_));
AND2X2 AND2X2_3974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6365_));
AND2X2 AND2X2_3975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6366_));
AND2X2 AND2X2_3976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6368_));
AND2X2 AND2X2_3977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6369_));
AND2X2 AND2X2_3978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6373_));
AND2X2 AND2X2_3979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6374_));
AND2X2 AND2X2_398 ( .A(_abc_44694_new_n1207__bF_buf3), .B(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .Y(_abc_44694_new_n1330_));
AND2X2 AND2X2_3980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6376_));
AND2X2 AND2X2_3981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6377_));
AND2X2 AND2X2_3982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6380_));
AND2X2 AND2X2_3983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6381_));
AND2X2 AND2X2_3984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6383_));
AND2X2 AND2X2_3985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6384_));
AND2X2 AND2X2_3986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6390_));
AND2X2 AND2X2_3987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6391_));
AND2X2 AND2X2_3988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6393_));
AND2X2 AND2X2_3989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6394_));
AND2X2 AND2X2_399 ( .A(_abc_44694_new_n1330_), .B(_abc_44694_new_n1329_), .Y(_abc_44694_new_n1331_));
AND2X2 AND2X2_3990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6397_));
AND2X2 AND2X2_3991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6398_));
AND2X2 AND2X2_3992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6400_));
AND2X2 AND2X2_3993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6401_));
AND2X2 AND2X2_3994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6405_));
AND2X2 AND2X2_3995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6406_));
AND2X2 AND2X2_3996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6407_));
AND2X2 AND2X2_3997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6410_));
AND2X2 AND2X2_3998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6411_));
AND2X2 AND2X2_3999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6413_));
AND2X2 AND2X2_4 ( .A(_abc_44694_new_n624_), .B(_abc_44694_new_n625_), .Y(_abc_44694_new_n626_));
AND2X2 AND2X2_40 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[24] ), .Y(_abc_44694_new_n686_));
AND2X2 AND2X2_400 ( .A(_abc_44694_new_n1332_), .B(enable_i_bF_buf0), .Y(_0sr_q_31_0__10_));
AND2X2 AND2X2_4000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6414_));
AND2X2 AND2X2_4001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6419_));
AND2X2 AND2X2_4002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6420_));
AND2X2 AND2X2_4003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6422_));
AND2X2 AND2X2_4004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6423_));
AND2X2 AND2X2_4005 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6426_));
AND2X2 AND2X2_4006 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6427_));
AND2X2 AND2X2_4007 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6429_));
AND2X2 AND2X2_4008 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6430_));
AND2X2 AND2X2_4009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6434_));
AND2X2 AND2X2_401 ( .A(_abc_44694_new_n1194__bF_buf3), .B(next_pc_r_0_), .Y(_abc_44694_new_n1335_));
AND2X2 AND2X2_4010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6435_));
AND2X2 AND2X2_4011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6437_));
AND2X2 AND2X2_4012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6438_));
AND2X2 AND2X2_4013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6441_));
AND2X2 AND2X2_4014 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6442_));
AND2X2 AND2X2_4015 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6444_));
AND2X2 AND2X2_4016 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6445_));
AND2X2 AND2X2_4017 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6451_));
AND2X2 AND2X2_4018 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6452_));
AND2X2 AND2X2_4019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6454_));
AND2X2 AND2X2_402 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_0_), .Y(_abc_44694_new_n1336_));
AND2X2 AND2X2_4020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6455_));
AND2X2 AND2X2_4021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6458_));
AND2X2 AND2X2_4022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6459_));
AND2X2 AND2X2_4023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6461_));
AND2X2 AND2X2_4024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6462_));
AND2X2 AND2X2_4025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6466_));
AND2X2 AND2X2_4026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6467_));
AND2X2 AND2X2_4027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6468_));
AND2X2 AND2X2_4028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6471_));
AND2X2 AND2X2_4029 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6472_));
AND2X2 AND2X2_403 ( .A(_abc_44694_new_n1339_), .B(_abc_44694_new_n1341_), .Y(_abc_44694_new_n1342_));
AND2X2 AND2X2_4030 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6474_));
AND2X2 AND2X2_4031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6475_));
AND2X2 AND2X2_4032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6480_));
AND2X2 AND2X2_4033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6481_));
AND2X2 AND2X2_4034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6483_));
AND2X2 AND2X2_4035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6484_));
AND2X2 AND2X2_4036 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6487_));
AND2X2 AND2X2_4037 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6488_));
AND2X2 AND2X2_4038 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6490_));
AND2X2 AND2X2_4039 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6491_));
AND2X2 AND2X2_404 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n1342_), .Y(_abc_44694_new_n1343_));
AND2X2 AND2X2_4040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6495_));
AND2X2 AND2X2_4041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6496_));
AND2X2 AND2X2_4042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6498_));
AND2X2 AND2X2_4043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6499_));
AND2X2 AND2X2_4044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6502_));
AND2X2 AND2X2_4045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6503_));
AND2X2 AND2X2_4046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6505_));
AND2X2 AND2X2_4047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6506_));
AND2X2 AND2X2_4048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6512_));
AND2X2 AND2X2_4049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6513_));
AND2X2 AND2X2_405 ( .A(_abc_44694_new_n1032_), .B(_abc_44694_new_n990_), .Y(_abc_44694_new_n1344_));
AND2X2 AND2X2_4050 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6515_));
AND2X2 AND2X2_4051 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6516_));
AND2X2 AND2X2_4052 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6519_));
AND2X2 AND2X2_4053 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6520_));
AND2X2 AND2X2_4054 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6522_));
AND2X2 AND2X2_4055 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6523_));
AND2X2 AND2X2_4056 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6527_));
AND2X2 AND2X2_4057 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6528_));
AND2X2 AND2X2_4058 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6529_));
AND2X2 AND2X2_4059 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6532_));
AND2X2 AND2X2_406 ( .A(_abc_44694_new_n1003_), .B(_abc_44694_new_n1344_), .Y(_abc_44694_new_n1345_));
AND2X2 AND2X2_4060 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6533_));
AND2X2 AND2X2_4061 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6535_));
AND2X2 AND2X2_4062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6536_));
AND2X2 AND2X2_4063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6541_));
AND2X2 AND2X2_4064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6542_));
AND2X2 AND2X2_4065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6544_));
AND2X2 AND2X2_4066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6545_));
AND2X2 AND2X2_4067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6548_));
AND2X2 AND2X2_4068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6549_));
AND2X2 AND2X2_4069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6551_));
AND2X2 AND2X2_407 ( .A(_abc_44694_new_n1031_), .B(_abc_44694_new_n1345_), .Y(_abc_44694_new_n1346_));
AND2X2 AND2X2_4070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6552_));
AND2X2 AND2X2_4071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6556_));
AND2X2 AND2X2_4072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6557_));
AND2X2 AND2X2_4073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6559_));
AND2X2 AND2X2_4074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6560_));
AND2X2 AND2X2_4075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6563_));
AND2X2 AND2X2_4076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6564_));
AND2X2 AND2X2_4077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6566_));
AND2X2 AND2X2_4078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6567_));
AND2X2 AND2X2_4079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6573_));
AND2X2 AND2X2_408 ( .A(_abc_44694_new_n1346_), .B(_abc_44694_new_n989_), .Y(_abc_44694_new_n1347_));
AND2X2 AND2X2_4080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6574_));
AND2X2 AND2X2_4081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6576_));
AND2X2 AND2X2_4082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6577_));
AND2X2 AND2X2_4083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6580_));
AND2X2 AND2X2_4084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6581_));
AND2X2 AND2X2_4085 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6583_));
AND2X2 AND2X2_4086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6584_));
AND2X2 AND2X2_4087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6588_));
AND2X2 AND2X2_4088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6589_));
AND2X2 AND2X2_4089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6590_));
AND2X2 AND2X2_409 ( .A(_abc_44694_new_n1347__bF_buf4), .B(_abc_44694_new_n970_), .Y(_abc_44694_new_n1348_));
AND2X2 AND2X2_4090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6593_));
AND2X2 AND2X2_4091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6594_));
AND2X2 AND2X2_4092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6596_));
AND2X2 AND2X2_4093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6597_));
AND2X2 AND2X2_4094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6602_));
AND2X2 AND2X2_4095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6603_));
AND2X2 AND2X2_4096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6605_));
AND2X2 AND2X2_4097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6606_));
AND2X2 AND2X2_4098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6609_));
AND2X2 AND2X2_4099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6610_));
AND2X2 AND2X2_41 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[8] ), .Y(_abc_44694_new_n687_));
AND2X2 AND2X2_410 ( .A(_abc_44694_new_n1348__bF_buf4), .B(_abc_44694_new_n1350_), .Y(_abc_44694_new_n1351_));
AND2X2 AND2X2_4100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6612_));
AND2X2 AND2X2_4101 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6613_));
AND2X2 AND2X2_4102 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6617_));
AND2X2 AND2X2_4103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6618_));
AND2X2 AND2X2_4104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6620_));
AND2X2 AND2X2_4105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6621_));
AND2X2 AND2X2_4106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6624_));
AND2X2 AND2X2_4107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6625_));
AND2X2 AND2X2_4108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6627_));
AND2X2 AND2X2_4109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6628_));
AND2X2 AND2X2_411 ( .A(_abc_44694_new_n1352_), .B(_abc_44694_new_n1349_), .Y(_abc_44694_new_n1353_));
AND2X2 AND2X2_4110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6634_));
AND2X2 AND2X2_4111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6635_));
AND2X2 AND2X2_4112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6637_));
AND2X2 AND2X2_4113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6638_));
AND2X2 AND2X2_4114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6641_));
AND2X2 AND2X2_4115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6642_));
AND2X2 AND2X2_4116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6644_));
AND2X2 AND2X2_4117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6645_));
AND2X2 AND2X2_4118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6649_));
AND2X2 AND2X2_4119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6650_));
AND2X2 AND2X2_412 ( .A(_abc_44694_new_n1278__bF_buf2), .B(_abc_44694_new_n1353_), .Y(_abc_44694_new_n1354_));
AND2X2 AND2X2_4120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6651_));
AND2X2 AND2X2_4121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6654_));
AND2X2 AND2X2_4122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6655_));
AND2X2 AND2X2_4123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6657_));
AND2X2 AND2X2_4124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6658_));
AND2X2 AND2X2_4125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6663_));
AND2X2 AND2X2_4126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6664_));
AND2X2 AND2X2_4127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6666_));
AND2X2 AND2X2_4128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6667_));
AND2X2 AND2X2_4129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6670_));
AND2X2 AND2X2_413 ( .A(_abc_44694_new_n1355_), .B(_abc_44694_new_n1207__bF_buf2), .Y(_abc_44694_new_n1356_));
AND2X2 AND2X2_4130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6671_));
AND2X2 AND2X2_4131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6673_));
AND2X2 AND2X2_4132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6674_));
AND2X2 AND2X2_4133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6678_));
AND2X2 AND2X2_4134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6679_));
AND2X2 AND2X2_4135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6681_));
AND2X2 AND2X2_4136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6682_));
AND2X2 AND2X2_4137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6685_));
AND2X2 AND2X2_4138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6686_));
AND2X2 AND2X2_4139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6688_));
AND2X2 AND2X2_414 ( .A(_abc_44694_new_n1359_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n1360_));
AND2X2 AND2X2_4140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6689_));
AND2X2 AND2X2_4141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6695_));
AND2X2 AND2X2_4142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6696_));
AND2X2 AND2X2_4143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6698_));
AND2X2 AND2X2_4144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6699_));
AND2X2 AND2X2_4145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6702_));
AND2X2 AND2X2_4146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6703_));
AND2X2 AND2X2_4147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6705_));
AND2X2 AND2X2_4148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6706_));
AND2X2 AND2X2_4149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6710_));
AND2X2 AND2X2_415 ( .A(_abc_44694_new_n1358_), .B(_abc_44694_new_n1360_), .Y(_0epc_q_31_0__0_));
AND2X2 AND2X2_4150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6711_));
AND2X2 AND2X2_4151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6712_));
AND2X2 AND2X2_4152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6715_));
AND2X2 AND2X2_4153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6716_));
AND2X2 AND2X2_4154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6718_));
AND2X2 AND2X2_4155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6719_));
AND2X2 AND2X2_4156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6724_));
AND2X2 AND2X2_4157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6725_));
AND2X2 AND2X2_4158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6727_));
AND2X2 AND2X2_4159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6728_));
AND2X2 AND2X2_416 ( .A(_abc_44694_new_n1194__bF_buf2), .B(next_pc_r_1_), .Y(_abc_44694_new_n1362_));
AND2X2 AND2X2_4160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6731_));
AND2X2 AND2X2_4161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6732_));
AND2X2 AND2X2_4162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6734_));
AND2X2 AND2X2_4163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6735_));
AND2X2 AND2X2_4164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6739_));
AND2X2 AND2X2_4165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6740_));
AND2X2 AND2X2_4166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6742_));
AND2X2 AND2X2_4167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6743_));
AND2X2 AND2X2_4168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6746_));
AND2X2 AND2X2_4169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6747_));
AND2X2 AND2X2_417 ( .A(_abc_44694_new_n1019__bF_buf4), .B(epc_q_1_), .Y(_abc_44694_new_n1363_));
AND2X2 AND2X2_4170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6749_));
AND2X2 AND2X2_4171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6750_));
AND2X2 AND2X2_4172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6756_));
AND2X2 AND2X2_4173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6757_));
AND2X2 AND2X2_4174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6759_));
AND2X2 AND2X2_4175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6760_));
AND2X2 AND2X2_4176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6763_));
AND2X2 AND2X2_4177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6764_));
AND2X2 AND2X2_4178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6766_));
AND2X2 AND2X2_4179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6767_));
AND2X2 AND2X2_418 ( .A(_abc_44694_new_n1365_), .B(_abc_44694_new_n1366_), .Y(_abc_44694_new_n1367_));
AND2X2 AND2X2_4180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6771_));
AND2X2 AND2X2_4181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6772_));
AND2X2 AND2X2_4182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6773_));
AND2X2 AND2X2_4183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6776_));
AND2X2 AND2X2_4184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6777_));
AND2X2 AND2X2_4185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6779_));
AND2X2 AND2X2_4186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6780_));
AND2X2 AND2X2_4187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6785_));
AND2X2 AND2X2_4188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6786_));
AND2X2 AND2X2_4189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6788_));
AND2X2 AND2X2_419 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n1367_), .Y(_abc_44694_new_n1368_));
AND2X2 AND2X2_4190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6789_));
AND2X2 AND2X2_4191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6792_));
AND2X2 AND2X2_4192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6793_));
AND2X2 AND2X2_4193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6795_));
AND2X2 AND2X2_4194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6796_));
AND2X2 AND2X2_4195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6800_));
AND2X2 AND2X2_4196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6801_));
AND2X2 AND2X2_4197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6803_));
AND2X2 AND2X2_4198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6804_));
AND2X2 AND2X2_4199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6807_));
AND2X2 AND2X2_42 ( .A(_abc_44694_new_n680_), .B(mem_offset_q_0_), .Y(_abc_44694_new_n689_));
AND2X2 AND2X2_420 ( .A(_abc_44694_new_n1348__bF_buf2), .B(_abc_44694_new_n1370_), .Y(_abc_44694_new_n1371_));
AND2X2 AND2X2_4200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6808_));
AND2X2 AND2X2_4201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6810_));
AND2X2 AND2X2_4202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6811_));
AND2X2 AND2X2_4203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6817_));
AND2X2 AND2X2_4204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6818_));
AND2X2 AND2X2_4205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6820_));
AND2X2 AND2X2_4206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6821_));
AND2X2 AND2X2_4207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6824_));
AND2X2 AND2X2_4208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6825_));
AND2X2 AND2X2_4209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6827_));
AND2X2 AND2X2_421 ( .A(_abc_44694_new_n1372_), .B(_abc_44694_new_n1369_), .Y(_abc_44694_new_n1373_));
AND2X2 AND2X2_4210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6828_));
AND2X2 AND2X2_4211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6832_));
AND2X2 AND2X2_4212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6833_));
AND2X2 AND2X2_4213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6834_));
AND2X2 AND2X2_4214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6837_));
AND2X2 AND2X2_4215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6838_));
AND2X2 AND2X2_4216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6840_));
AND2X2 AND2X2_4217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6841_));
AND2X2 AND2X2_4218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6846_));
AND2X2 AND2X2_4219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6847_));
AND2X2 AND2X2_422 ( .A(_abc_44694_new_n1278__bF_buf1), .B(_abc_44694_new_n1373_), .Y(_abc_44694_new_n1374_));
AND2X2 AND2X2_4220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6849_));
AND2X2 AND2X2_4221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6850_));
AND2X2 AND2X2_4222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6853_));
AND2X2 AND2X2_4223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6854_));
AND2X2 AND2X2_4224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6856_));
AND2X2 AND2X2_4225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6857_));
AND2X2 AND2X2_4226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6861_));
AND2X2 AND2X2_4227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6862_));
AND2X2 AND2X2_4228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6864_));
AND2X2 AND2X2_4229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6865_));
AND2X2 AND2X2_423 ( .A(_abc_44694_new_n1375_), .B(_abc_44694_new_n1207__bF_buf1), .Y(_abc_44694_new_n1376_));
AND2X2 AND2X2_4230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6868_));
AND2X2 AND2X2_4231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6869_));
AND2X2 AND2X2_4232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6871_));
AND2X2 AND2X2_4233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6872_));
AND2X2 AND2X2_4234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6878_));
AND2X2 AND2X2_4235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6879_));
AND2X2 AND2X2_4236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6881_));
AND2X2 AND2X2_4237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6882_));
AND2X2 AND2X2_4238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6885_));
AND2X2 AND2X2_4239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6886_));
AND2X2 AND2X2_424 ( .A(_abc_44694_new_n1379_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n1380_));
AND2X2 AND2X2_4240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6888_));
AND2X2 AND2X2_4241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6889_));
AND2X2 AND2X2_4242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6893_));
AND2X2 AND2X2_4243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6894_));
AND2X2 AND2X2_4244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6895_));
AND2X2 AND2X2_4245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6898_));
AND2X2 AND2X2_4246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6899_));
AND2X2 AND2X2_4247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6901_));
AND2X2 AND2X2_4248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6902_));
AND2X2 AND2X2_4249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6907_));
AND2X2 AND2X2_425 ( .A(_abc_44694_new_n1378_), .B(_abc_44694_new_n1380_), .Y(_0epc_q_31_0__1_));
AND2X2 AND2X2_4250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6908_));
AND2X2 AND2X2_4251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6910_));
AND2X2 AND2X2_4252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6911_));
AND2X2 AND2X2_4253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6914_));
AND2X2 AND2X2_4254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6915_));
AND2X2 AND2X2_4255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6917_));
AND2X2 AND2X2_4256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6918_));
AND2X2 AND2X2_4257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6922_));
AND2X2 AND2X2_4258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6923_));
AND2X2 AND2X2_4259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6925_));
AND2X2 AND2X2_426 ( .A(_abc_44694_new_n1348__bF_buf1), .B(_abc_44694_new_n1383_), .Y(_abc_44694_new_n1384_));
AND2X2 AND2X2_4260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6926_));
AND2X2 AND2X2_4261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6929_));
AND2X2 AND2X2_4262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6930_));
AND2X2 AND2X2_4263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6932_));
AND2X2 AND2X2_4264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6933_));
AND2X2 AND2X2_4265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6939_));
AND2X2 AND2X2_4266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6940_));
AND2X2 AND2X2_4267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6942_));
AND2X2 AND2X2_4268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6943_));
AND2X2 AND2X2_4269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6946_));
AND2X2 AND2X2_427 ( .A(_abc_44694_new_n1385_), .B(_abc_44694_new_n1386_), .Y(_abc_44694_new_n1387_));
AND2X2 AND2X2_4270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6947_));
AND2X2 AND2X2_4271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6949_));
AND2X2 AND2X2_4272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6950_));
AND2X2 AND2X2_4273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6954_));
AND2X2 AND2X2_4274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6955_));
AND2X2 AND2X2_4275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6956_));
AND2X2 AND2X2_4276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6959_));
AND2X2 AND2X2_4277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6960_));
AND2X2 AND2X2_4278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6962_));
AND2X2 AND2X2_4279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6963_));
AND2X2 AND2X2_428 ( .A(_abc_44694_new_n1117_), .B(_abc_44694_new_n646_), .Y(_abc_44694_new_n1390_));
AND2X2 AND2X2_4280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6968_));
AND2X2 AND2X2_4281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6969_));
AND2X2 AND2X2_4282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6971_));
AND2X2 AND2X2_4283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6972_));
AND2X2 AND2X2_4284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6975_));
AND2X2 AND2X2_4285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6976_));
AND2X2 AND2X2_4286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6978_));
AND2X2 AND2X2_4287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6979_));
AND2X2 AND2X2_4288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6983_));
AND2X2 AND2X2_4289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6984_));
AND2X2 AND2X2_429 ( .A(_abc_44694_new_n640_), .B(_abc_44694_new_n619_), .Y(_abc_44694_new_n1393_));
AND2X2 AND2X2_4290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6986_));
AND2X2 AND2X2_4291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6987_));
AND2X2 AND2X2_4292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6990_));
AND2X2 AND2X2_4293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6991_));
AND2X2 AND2X2_4294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6993_));
AND2X2 AND2X2_4295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6994_));
AND2X2 AND2X2_4296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7000_));
AND2X2 AND2X2_4297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7001_));
AND2X2 AND2X2_4298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7003_));
AND2X2 AND2X2_4299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7004_));
AND2X2 AND2X2_43 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[16] ), .Y(_abc_44694_new_n690_));
AND2X2 AND2X2_430 ( .A(_abc_44694_new_n1393_), .B(sr_q_9_), .Y(_abc_44694_new_n1394_));
AND2X2 AND2X2_4300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7007_));
AND2X2 AND2X2_4301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7008_));
AND2X2 AND2X2_4302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7010_));
AND2X2 AND2X2_4303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7011_));
AND2X2 AND2X2_4304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7015_));
AND2X2 AND2X2_4305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7016_));
AND2X2 AND2X2_4306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7017_));
AND2X2 AND2X2_4307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7020_));
AND2X2 AND2X2_4308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7021_));
AND2X2 AND2X2_4309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7023_));
AND2X2 AND2X2_431 ( .A(_abc_44694_new_n1392_), .B(_abc_44694_new_n1395_), .Y(_abc_44694_new_n1396_));
AND2X2 AND2X2_4310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7024_));
AND2X2 AND2X2_4311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7029_));
AND2X2 AND2X2_4312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7030_));
AND2X2 AND2X2_4313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7032_));
AND2X2 AND2X2_4314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7033_));
AND2X2 AND2X2_4315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7036_));
AND2X2 AND2X2_4316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7037_));
AND2X2 AND2X2_4317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7039_));
AND2X2 AND2X2_4318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7040_));
AND2X2 AND2X2_4319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7044_));
AND2X2 AND2X2_432 ( .A(_abc_44694_new_n619_), .B(sr_q_9_), .Y(_abc_44694_new_n1397_));
AND2X2 AND2X2_4320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7045_));
AND2X2 AND2X2_4321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7047_));
AND2X2 AND2X2_4322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7048_));
AND2X2 AND2X2_4323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7051_));
AND2X2 AND2X2_4324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7052_));
AND2X2 AND2X2_4325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7054_));
AND2X2 AND2X2_4326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7055_));
AND2X2 AND2X2_4327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7061_));
AND2X2 AND2X2_4328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7062_));
AND2X2 AND2X2_4329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7064_));
AND2X2 AND2X2_433 ( .A(_abc_44694_new_n642_), .B(_abc_44694_new_n1397_), .Y(_abc_44694_new_n1398_));
AND2X2 AND2X2_4330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7065_));
AND2X2 AND2X2_4331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7068_));
AND2X2 AND2X2_4332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7069_));
AND2X2 AND2X2_4333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7071_));
AND2X2 AND2X2_4334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7072_));
AND2X2 AND2X2_4335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7076_));
AND2X2 AND2X2_4336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7077_));
AND2X2 AND2X2_4337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7078_));
AND2X2 AND2X2_4338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7081_));
AND2X2 AND2X2_4339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7082_));
AND2X2 AND2X2_434 ( .A(alu_op_r_0_), .B(pc_q_2_), .Y(_abc_44694_new_n1403_));
AND2X2 AND2X2_4340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7084_));
AND2X2 AND2X2_4341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7085_));
AND2X2 AND2X2_4342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7090_));
AND2X2 AND2X2_4343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7091_));
AND2X2 AND2X2_4344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7093_));
AND2X2 AND2X2_4345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7094_));
AND2X2 AND2X2_4346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7097_));
AND2X2 AND2X2_4347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7098_));
AND2X2 AND2X2_4348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7100_));
AND2X2 AND2X2_4349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7101_));
AND2X2 AND2X2_435 ( .A(_abc_44694_new_n1404_), .B(_abc_44694_new_n1402_), .Y(_abc_44694_new_n1405_));
AND2X2 AND2X2_4350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7105_));
AND2X2 AND2X2_4351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7106_));
AND2X2 AND2X2_4352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7108_));
AND2X2 AND2X2_4353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7109_));
AND2X2 AND2X2_4354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7112_));
AND2X2 AND2X2_4355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7113_));
AND2X2 AND2X2_4356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7115_));
AND2X2 AND2X2_4357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7116_));
AND2X2 AND2X2_4358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7122_));
AND2X2 AND2X2_4359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7123_));
AND2X2 AND2X2_436 ( .A(_abc_44694_new_n1194__bF_buf0), .B(_abc_44694_new_n1405_), .Y(_abc_44694_new_n1406_));
AND2X2 AND2X2_4360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7125_));
AND2X2 AND2X2_4361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7126_));
AND2X2 AND2X2_4362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7129_));
AND2X2 AND2X2_4363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7130_));
AND2X2 AND2X2_4364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7132_));
AND2X2 AND2X2_4365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7133_));
AND2X2 AND2X2_4366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7137_));
AND2X2 AND2X2_4367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7138_));
AND2X2 AND2X2_4368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7139_));
AND2X2 AND2X2_4369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7142_));
AND2X2 AND2X2_437 ( .A(_abc_44694_new_n1019__bF_buf3), .B(epc_q_2_), .Y(_abc_44694_new_n1407_));
AND2X2 AND2X2_4370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7143_));
AND2X2 AND2X2_4371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7145_));
AND2X2 AND2X2_4372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7146_));
AND2X2 AND2X2_4373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7151_));
AND2X2 AND2X2_4374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7152_));
AND2X2 AND2X2_4375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7154_));
AND2X2 AND2X2_4376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7155_));
AND2X2 AND2X2_4377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7158_));
AND2X2 AND2X2_4378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7159_));
AND2X2 AND2X2_4379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7161_));
AND2X2 AND2X2_438 ( .A(_abc_44694_new_n1409_), .B(_abc_44694_new_n1401_), .Y(_abc_44694_new_n1410_));
AND2X2 AND2X2_4380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7162_));
AND2X2 AND2X2_4381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7166_));
AND2X2 AND2X2_4382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7167_));
AND2X2 AND2X2_4383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7169_));
AND2X2 AND2X2_4384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7170_));
AND2X2 AND2X2_4385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7173_));
AND2X2 AND2X2_4386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7174_));
AND2X2 AND2X2_4387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7176_));
AND2X2 AND2X2_4388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7177_));
AND2X2 AND2X2_4389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7183_));
AND2X2 AND2X2_439 ( .A(_abc_44694_new_n1411_), .B(_abc_44694_new_n1413_), .Y(_abc_44694_new_n1414_));
AND2X2 AND2X2_4390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7184_));
AND2X2 AND2X2_4391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7186_));
AND2X2 AND2X2_4392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7187_));
AND2X2 AND2X2_4393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7190_));
AND2X2 AND2X2_4394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7191_));
AND2X2 AND2X2_4395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7193_));
AND2X2 AND2X2_4396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7194_));
AND2X2 AND2X2_4397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7198_));
AND2X2 AND2X2_4398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7199_));
AND2X2 AND2X2_4399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7200_));
AND2X2 AND2X2_44 ( .A(mem_offset_q_1_), .B(mem_offset_q_0_), .Y(_abc_44694_new_n691_));
AND2X2 AND2X2_440 ( .A(_abc_44694_new_n1388_), .B(_abc_44694_new_n1415_), .Y(_abc_44694_new_n1416_));
AND2X2 AND2X2_4400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7203_));
AND2X2 AND2X2_4401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7204_));
AND2X2 AND2X2_4402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7206_));
AND2X2 AND2X2_4403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7207_));
AND2X2 AND2X2_4404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7212_));
AND2X2 AND2X2_4405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7213_));
AND2X2 AND2X2_4406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7215_));
AND2X2 AND2X2_4407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7216_));
AND2X2 AND2X2_4408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7219_));
AND2X2 AND2X2_4409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7220_));
AND2X2 AND2X2_441 ( .A(_abc_44694_new_n1417_), .B(_abc_44694_new_n1418_), .Y(_abc_44694_new_n1419_));
AND2X2 AND2X2_4410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7222_));
AND2X2 AND2X2_4411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7223_));
AND2X2 AND2X2_4412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7227_));
AND2X2 AND2X2_4413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7228_));
AND2X2 AND2X2_4414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7230_));
AND2X2 AND2X2_4415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7231_));
AND2X2 AND2X2_4416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7234_));
AND2X2 AND2X2_4417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7235_));
AND2X2 AND2X2_4418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7237_));
AND2X2 AND2X2_4419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7238_));
AND2X2 AND2X2_442 ( .A(_abc_44694_new_n1421_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n1422_));
AND2X2 AND2X2_4420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7244_));
AND2X2 AND2X2_4421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7245_));
AND2X2 AND2X2_4422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7247_));
AND2X2 AND2X2_4423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7248_));
AND2X2 AND2X2_4424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7251_));
AND2X2 AND2X2_4425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7252_));
AND2X2 AND2X2_4426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7254_));
AND2X2 AND2X2_4427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7255_));
AND2X2 AND2X2_4428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7259_));
AND2X2 AND2X2_4429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7260_));
AND2X2 AND2X2_443 ( .A(_abc_44694_new_n1420_), .B(_abc_44694_new_n1422_), .Y(_0epc_q_31_0__2_));
AND2X2 AND2X2_4430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7261_));
AND2X2 AND2X2_4431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7264_));
AND2X2 AND2X2_4432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7265_));
AND2X2 AND2X2_4433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7267_));
AND2X2 AND2X2_4434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7268_));
AND2X2 AND2X2_4435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7273_));
AND2X2 AND2X2_4436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7274_));
AND2X2 AND2X2_4437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7276_));
AND2X2 AND2X2_4438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7277_));
AND2X2 AND2X2_4439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7280_));
AND2X2 AND2X2_444 ( .A(_abc_44694_new_n1348__bF_buf5), .B(_abc_44694_new_n1424_), .Y(_abc_44694_new_n1425_));
AND2X2 AND2X2_4440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7281_));
AND2X2 AND2X2_4441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7283_));
AND2X2 AND2X2_4442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7284_));
AND2X2 AND2X2_4443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7288_));
AND2X2 AND2X2_4444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7289_));
AND2X2 AND2X2_4445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7291_));
AND2X2 AND2X2_4446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7292_));
AND2X2 AND2X2_4447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7295_));
AND2X2 AND2X2_4448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7296_));
AND2X2 AND2X2_4449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7298_));
AND2X2 AND2X2_445 ( .A(_abc_44694_new_n1426_), .B(_abc_44694_new_n1427_), .Y(_abc_44694_new_n1428_));
AND2X2 AND2X2_4450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7299_));
AND2X2 AND2X2_4451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7305_));
AND2X2 AND2X2_4452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7306_));
AND2X2 AND2X2_4453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7308_));
AND2X2 AND2X2_4454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7309_));
AND2X2 AND2X2_4455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7312_));
AND2X2 AND2X2_4456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7313_));
AND2X2 AND2X2_4457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7315_));
AND2X2 AND2X2_4458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7316_));
AND2X2 AND2X2_4459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7320_));
AND2X2 AND2X2_446 ( .A(alu_op_r_1_), .B(pc_q_3_), .Y(_abc_44694_new_n1431_));
AND2X2 AND2X2_4460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7321_));
AND2X2 AND2X2_4461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7322_));
AND2X2 AND2X2_4462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7325_));
AND2X2 AND2X2_4463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7326_));
AND2X2 AND2X2_4464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7328_));
AND2X2 AND2X2_4465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7329_));
AND2X2 AND2X2_4466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7334_));
AND2X2 AND2X2_4467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7335_));
AND2X2 AND2X2_4468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7337_));
AND2X2 AND2X2_4469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7338_));
AND2X2 AND2X2_447 ( .A(_abc_44694_new_n1432_), .B(_abc_44694_new_n1430_), .Y(_abc_44694_new_n1433_));
AND2X2 AND2X2_4470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7341_));
AND2X2 AND2X2_4471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7342_));
AND2X2 AND2X2_4472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7344_));
AND2X2 AND2X2_4473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7345_));
AND2X2 AND2X2_4474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7349_));
AND2X2 AND2X2_4475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7350_));
AND2X2 AND2X2_4476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7352_));
AND2X2 AND2X2_4477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7353_));
AND2X2 AND2X2_4478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7356_));
AND2X2 AND2X2_4479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7357_));
AND2X2 AND2X2_448 ( .A(_abc_44694_new_n1433_), .B(_abc_44694_new_n1403_), .Y(_abc_44694_new_n1435_));
AND2X2 AND2X2_4480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7359_));
AND2X2 AND2X2_4481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7360_));
AND2X2 AND2X2_4482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7366_));
AND2X2 AND2X2_4483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7367_));
AND2X2 AND2X2_4484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7369_));
AND2X2 AND2X2_4485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7370_));
AND2X2 AND2X2_4486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7373_));
AND2X2 AND2X2_4487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7374_));
AND2X2 AND2X2_4488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7376_));
AND2X2 AND2X2_4489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7377_));
AND2X2 AND2X2_449 ( .A(_abc_44694_new_n1436_), .B(_abc_44694_new_n1434_), .Y(_abc_44694_new_n1437_));
AND2X2 AND2X2_4490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7381_));
AND2X2 AND2X2_4491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7382_));
AND2X2 AND2X2_4492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7383_));
AND2X2 AND2X2_4493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7386_));
AND2X2 AND2X2_4494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7387_));
AND2X2 AND2X2_4495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7389_));
AND2X2 AND2X2_4496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7390_));
AND2X2 AND2X2_4497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7395_));
AND2X2 AND2X2_4498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7396_));
AND2X2 AND2X2_4499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7398_));
AND2X2 AND2X2_45 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[0] ), .Y(_abc_44694_new_n692_));
AND2X2 AND2X2_450 ( .A(_abc_44694_new_n1194__bF_buf4), .B(_abc_44694_new_n1437_), .Y(_abc_44694_new_n1438_));
AND2X2 AND2X2_4500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7399_));
AND2X2 AND2X2_4501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7402_));
AND2X2 AND2X2_4502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7403_));
AND2X2 AND2X2_4503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7405_));
AND2X2 AND2X2_4504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7406_));
AND2X2 AND2X2_4505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7410_));
AND2X2 AND2X2_4506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7411_));
AND2X2 AND2X2_4507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7413_));
AND2X2 AND2X2_4508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7414_));
AND2X2 AND2X2_4509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7417_));
AND2X2 AND2X2_451 ( .A(_abc_44694_new_n1019__bF_buf2), .B(epc_q_3_), .Y(_abc_44694_new_n1439_));
AND2X2 AND2X2_4510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7418_));
AND2X2 AND2X2_4511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7420_));
AND2X2 AND2X2_4512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7421_));
AND2X2 AND2X2_4513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7427_));
AND2X2 AND2X2_4514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7428_));
AND2X2 AND2X2_4515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7430_));
AND2X2 AND2X2_4516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7431_));
AND2X2 AND2X2_4517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7434_));
AND2X2 AND2X2_4518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7435_));
AND2X2 AND2X2_4519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7437_));
AND2X2 AND2X2_452 ( .A(_abc_44694_new_n1441_), .B(_abc_44694_new_n1442_), .Y(_abc_44694_new_n1443_));
AND2X2 AND2X2_4520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7438_));
AND2X2 AND2X2_4521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7442_));
AND2X2 AND2X2_4522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7443_));
AND2X2 AND2X2_4523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7444_));
AND2X2 AND2X2_4524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7447_));
AND2X2 AND2X2_4525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7448_));
AND2X2 AND2X2_4526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7450_));
AND2X2 AND2X2_4527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7451_));
AND2X2 AND2X2_4528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7456_));
AND2X2 AND2X2_4529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7457_));
AND2X2 AND2X2_453 ( .A(_abc_44694_new_n1399__bF_buf2), .B(_abc_44694_new_n1443_), .Y(_abc_44694_new_n1444_));
AND2X2 AND2X2_4530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7459_));
AND2X2 AND2X2_4531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7460_));
AND2X2 AND2X2_4532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7463_));
AND2X2 AND2X2_4533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7464_));
AND2X2 AND2X2_4534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7466_));
AND2X2 AND2X2_4535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7467_));
AND2X2 AND2X2_4536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7471_));
AND2X2 AND2X2_4537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7472_));
AND2X2 AND2X2_4538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7474_));
AND2X2 AND2X2_4539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7475_));
AND2X2 AND2X2_454 ( .A(pc_q_2_), .B(pc_q_3_), .Y(_abc_44694_new_n1446_));
AND2X2 AND2X2_4540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7478_));
AND2X2 AND2X2_4541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7479_));
AND2X2 AND2X2_4542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7481_));
AND2X2 AND2X2_4543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7482_));
AND2X2 AND2X2_4544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7488_));
AND2X2 AND2X2_4545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7489_));
AND2X2 AND2X2_4546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7491_));
AND2X2 AND2X2_4547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7492_));
AND2X2 AND2X2_4548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7495_));
AND2X2 AND2X2_4549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7496_));
AND2X2 AND2X2_455 ( .A(_abc_44694_new_n1447_), .B(_abc_44694_new_n1445_), .Y(_abc_44694_new_n1448_));
AND2X2 AND2X2_4550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7498_));
AND2X2 AND2X2_4551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7499_));
AND2X2 AND2X2_4552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7503_));
AND2X2 AND2X2_4553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7504_));
AND2X2 AND2X2_4554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7505_));
AND2X2 AND2X2_4555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7508_));
AND2X2 AND2X2_4556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7509_));
AND2X2 AND2X2_4557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7511_));
AND2X2 AND2X2_4558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7512_));
AND2X2 AND2X2_4559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7517_));
AND2X2 AND2X2_456 ( .A(_abc_44694_new_n1400__bF_buf3), .B(_abc_44694_new_n1448_), .Y(_abc_44694_new_n1449_));
AND2X2 AND2X2_4560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7518_));
AND2X2 AND2X2_4561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7520_));
AND2X2 AND2X2_4562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7521_));
AND2X2 AND2X2_4563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7524_));
AND2X2 AND2X2_4564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7525_));
AND2X2 AND2X2_4565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7527_));
AND2X2 AND2X2_4566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7528_));
AND2X2 AND2X2_4567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7532_));
AND2X2 AND2X2_4568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7533_));
AND2X2 AND2X2_4569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7535_));
AND2X2 AND2X2_457 ( .A(_abc_44694_new_n1429_), .B(_abc_44694_new_n1451_), .Y(_abc_44694_new_n1452_));
AND2X2 AND2X2_4570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7536_));
AND2X2 AND2X2_4571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7539_));
AND2X2 AND2X2_4572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7540_));
AND2X2 AND2X2_4573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7542_));
AND2X2 AND2X2_4574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7543_));
AND2X2 AND2X2_4575 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7550_));
AND2X2 AND2X2_4576 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7551_));
AND2X2 AND2X2_4577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7550_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7551_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7552_));
AND2X2 AND2X2_4578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7552_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7553_));
AND2X2 AND2X2_4579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7554_));
AND2X2 AND2X2_458 ( .A(_abc_44694_new_n1453_), .B(_abc_44694_new_n1454_), .Y(_abc_44694_new_n1455_));
AND2X2 AND2X2_4580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7555_), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7556_));
AND2X2 AND2X2_4581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7551_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7557_));
AND2X2 AND2X2_4582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7557_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7558_));
AND2X2 AND2X2_4583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7559_));
AND2X2 AND2X2_4584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7561_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7555_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7562_));
AND2X2 AND2X2_4585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7562_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7563_));
AND2X2 AND2X2_4586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7551_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7564_));
AND2X2 AND2X2_4587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7565_));
AND2X2 AND2X2_4588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7561_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7566_));
AND2X2 AND2X2_4589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7566_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7551_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7567_));
AND2X2 AND2X2_459 ( .A(_abc_44694_new_n1457_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n1458_));
AND2X2 AND2X2_4590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7567_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7568_));
AND2X2 AND2X2_4591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7569_));
AND2X2 AND2X2_4592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7572_), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7573_));
AND2X2 AND2X2_4593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7573_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7556_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7574_));
AND2X2 AND2X2_4594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7574_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7575_));
AND2X2 AND2X2_4595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7576_));
AND2X2 AND2X2_4596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7573_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7550_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7577_));
AND2X2 AND2X2_4597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7577_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7578_));
AND2X2 AND2X2_4598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7579_));
AND2X2 AND2X2_4599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7566_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7573_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7581_));
AND2X2 AND2X2_46 ( .A(_abc_44694_new_n694_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n695_));
AND2X2 AND2X2_460 ( .A(_abc_44694_new_n1456_), .B(_abc_44694_new_n1458_), .Y(_0epc_q_31_0__3_));
AND2X2 AND2X2_4600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7581_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7582_));
AND2X2 AND2X2_4601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7583_));
AND2X2 AND2X2_4602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7573_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7584_));
AND2X2 AND2X2_4603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7585_));
AND2X2 AND2X2_4604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7589_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7572_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7590_));
AND2X2 AND2X2_4605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7590_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7591_));
AND2X2 AND2X2_4606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7591_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7592_));
AND2X2 AND2X2_4607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7593_));
AND2X2 AND2X2_4608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7590_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7556_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7594_));
AND2X2 AND2X2_4609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7594_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7595_));
AND2X2 AND2X2_461 ( .A(_abc_44694_new_n1348__bF_buf3), .B(_abc_44694_new_n1460_), .Y(_abc_44694_new_n1461_));
AND2X2 AND2X2_4610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7596_));
AND2X2 AND2X2_4611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7590_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7550_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7597_));
AND2X2 AND2X2_4612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7597_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7598_));
AND2X2 AND2X2_4613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7599_));
AND2X2 AND2X2_4614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7589_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7602_));
AND2X2 AND2X2_4615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7566_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7603_));
AND2X2 AND2X2_4616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7603_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7604_));
AND2X2 AND2X2_4617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7605_));
AND2X2 AND2X2_4618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7606_));
AND2X2 AND2X2_4619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7607_));
AND2X2 AND2X2_462 ( .A(_abc_44694_new_n1462_), .B(_abc_44694_new_n1463_), .Y(_abc_44694_new_n1464_));
AND2X2 AND2X2_4620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7602_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7550_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7609_));
AND2X2 AND2X2_4621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7609_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7610_));
AND2X2 AND2X2_4622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7611_));
AND2X2 AND2X2_4623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7612_));
AND2X2 AND2X2_4624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7612_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7613_));
AND2X2 AND2X2_4625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7614_));
AND2X2 AND2X2_4626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7552_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7619_));
AND2X2 AND2X2_4627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7620_));
AND2X2 AND2X2_4628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7557_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7621_));
AND2X2 AND2X2_4629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7622_));
AND2X2 AND2X2_463 ( .A(_abc_44694_new_n1436_), .B(_abc_44694_new_n1432_), .Y(_abc_44694_new_n1466_));
AND2X2 AND2X2_4630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7562_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7624_));
AND2X2 AND2X2_4631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7551_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7625_));
AND2X2 AND2X2_4632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7626_));
AND2X2 AND2X2_4633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7567_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7627_));
AND2X2 AND2X2_4634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7628_));
AND2X2 AND2X2_4635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7581_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7631_));
AND2X2 AND2X2_4636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7632_));
AND2X2 AND2X2_4637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7573_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7633_));
AND2X2 AND2X2_4638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7634_));
AND2X2 AND2X2_4639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7574_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7636_));
AND2X2 AND2X2_464 ( .A(alu_op_r_2_), .B(pc_q_4_), .Y(_abc_44694_new_n1468_));
AND2X2 AND2X2_4640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7637_));
AND2X2 AND2X2_4641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7577_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7638_));
AND2X2 AND2X2_4642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7639_));
AND2X2 AND2X2_4643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7591_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7643_));
AND2X2 AND2X2_4644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7644_));
AND2X2 AND2X2_4645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7590_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7645_));
AND2X2 AND2X2_4646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7646_));
AND2X2 AND2X2_4647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7594_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7648_));
AND2X2 AND2X2_4648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7649_));
AND2X2 AND2X2_4649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7597_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7650_));
AND2X2 AND2X2_465 ( .A(_abc_44694_new_n1469_), .B(_abc_44694_new_n1467_), .Y(_abc_44694_new_n1470_));
AND2X2 AND2X2_4650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7651_));
AND2X2 AND2X2_4651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7654_));
AND2X2 AND2X2_4652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7655_));
AND2X2 AND2X2_4653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7603_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7656_));
AND2X2 AND2X2_4654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7657_));
AND2X2 AND2X2_4655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7612_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7659_));
AND2X2 AND2X2_4656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7660_));
AND2X2 AND2X2_4657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7609_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7661_));
AND2X2 AND2X2_4658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7662_));
AND2X2 AND2X2_4659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7668_));
AND2X2 AND2X2_466 ( .A(_abc_44694_new_n1474_), .B(_abc_44694_new_n1472_), .Y(_abc_44694_new_n1475_));
AND2X2 AND2X2_4660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7669_));
AND2X2 AND2X2_4661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7671_));
AND2X2 AND2X2_4662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7672_));
AND2X2 AND2X2_4663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7675_));
AND2X2 AND2X2_4664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7676_));
AND2X2 AND2X2_4665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7678_));
AND2X2 AND2X2_4666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7679_));
AND2X2 AND2X2_4667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7683_));
AND2X2 AND2X2_4668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7684_));
AND2X2 AND2X2_4669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7685_));
AND2X2 AND2X2_467 ( .A(_abc_44694_new_n1475_), .B(_abc_44694_new_n1194__bF_buf3), .Y(_abc_44694_new_n1476_));
AND2X2 AND2X2_4670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7688_));
AND2X2 AND2X2_4671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7689_));
AND2X2 AND2X2_4672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7691_));
AND2X2 AND2X2_4673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7692_));
AND2X2 AND2X2_4674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7697_));
AND2X2 AND2X2_4675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7698_));
AND2X2 AND2X2_4676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7700_));
AND2X2 AND2X2_4677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7701_));
AND2X2 AND2X2_4678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7704_));
AND2X2 AND2X2_4679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7705_));
AND2X2 AND2X2_468 ( .A(_abc_44694_new_n1019__bF_buf1), .B(epc_q_4_), .Y(_abc_44694_new_n1477_));
AND2X2 AND2X2_4680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7707_));
AND2X2 AND2X2_4681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7708_));
AND2X2 AND2X2_4682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7712_));
AND2X2 AND2X2_4683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7713_));
AND2X2 AND2X2_4684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7715_));
AND2X2 AND2X2_4685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7716_));
AND2X2 AND2X2_4686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7719_));
AND2X2 AND2X2_4687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7720_));
AND2X2 AND2X2_4688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7722_));
AND2X2 AND2X2_4689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7723_));
AND2X2 AND2X2_469 ( .A(_abc_44694_new_n1479_), .B(_abc_44694_new_n1480_), .Y(_abc_44694_new_n1481_));
AND2X2 AND2X2_4690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7729_));
AND2X2 AND2X2_4691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7730_));
AND2X2 AND2X2_4692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7732_));
AND2X2 AND2X2_4693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7733_));
AND2X2 AND2X2_4694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7736_));
AND2X2 AND2X2_4695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7737_));
AND2X2 AND2X2_4696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7739_));
AND2X2 AND2X2_4697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7740_));
AND2X2 AND2X2_4698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7744_));
AND2X2 AND2X2_4699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7745_));
AND2X2 AND2X2_47 ( .A(_abc_44694_new_n696_), .B(state_q_1_bF_buf1_), .Y(_abc_44694_new_n697_));
AND2X2 AND2X2_470 ( .A(_abc_44694_new_n1399__bF_buf1), .B(_abc_44694_new_n1481_), .Y(_abc_44694_new_n1482_));
AND2X2 AND2X2_4700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7746_));
AND2X2 AND2X2_4701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7749_));
AND2X2 AND2X2_4702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7750_));
AND2X2 AND2X2_4703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7752_));
AND2X2 AND2X2_4704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7753_));
AND2X2 AND2X2_4705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7758_));
AND2X2 AND2X2_4706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7759_));
AND2X2 AND2X2_4707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7761_));
AND2X2 AND2X2_4708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7762_));
AND2X2 AND2X2_4709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7765_));
AND2X2 AND2X2_471 ( .A(_abc_44694_new_n1446_), .B(pc_q_4_), .Y(_abc_44694_new_n1484_));
AND2X2 AND2X2_4710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7766_));
AND2X2 AND2X2_4711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7768_));
AND2X2 AND2X2_4712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7769_));
AND2X2 AND2X2_4713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7773_));
AND2X2 AND2X2_4714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7774_));
AND2X2 AND2X2_4715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7776_));
AND2X2 AND2X2_4716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7777_));
AND2X2 AND2X2_4717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7780_));
AND2X2 AND2X2_4718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7781_));
AND2X2 AND2X2_4719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7783_));
AND2X2 AND2X2_472 ( .A(_abc_44694_new_n1485_), .B(_abc_44694_new_n1483_), .Y(_abc_44694_new_n1486_));
AND2X2 AND2X2_4720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7784_));
AND2X2 AND2X2_4721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7790_));
AND2X2 AND2X2_4722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7791_));
AND2X2 AND2X2_4723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7793_));
AND2X2 AND2X2_4724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7794_));
AND2X2 AND2X2_4725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7797_));
AND2X2 AND2X2_4726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7798_));
AND2X2 AND2X2_4727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7800_));
AND2X2 AND2X2_4728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7801_));
AND2X2 AND2X2_4729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7805_));
AND2X2 AND2X2_473 ( .A(_abc_44694_new_n1400__bF_buf2), .B(_abc_44694_new_n1486_), .Y(_abc_44694_new_n1487_));
AND2X2 AND2X2_4730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7806_));
AND2X2 AND2X2_4731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7807_));
AND2X2 AND2X2_4732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7810_));
AND2X2 AND2X2_4733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7811_));
AND2X2 AND2X2_4734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7813_));
AND2X2 AND2X2_4735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7814_));
AND2X2 AND2X2_4736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7819_));
AND2X2 AND2X2_4737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7820_));
AND2X2 AND2X2_4738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7822_));
AND2X2 AND2X2_4739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7823_));
AND2X2 AND2X2_474 ( .A(_abc_44694_new_n1465_), .B(_abc_44694_new_n1489_), .Y(_abc_44694_new_n1490_));
AND2X2 AND2X2_4740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7826_));
AND2X2 AND2X2_4741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7827_));
AND2X2 AND2X2_4742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7829_));
AND2X2 AND2X2_4743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7830_));
AND2X2 AND2X2_4744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7834_));
AND2X2 AND2X2_4745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7835_));
AND2X2 AND2X2_4746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7837_));
AND2X2 AND2X2_4747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7838_));
AND2X2 AND2X2_4748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7841_));
AND2X2 AND2X2_4749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7842_));
AND2X2 AND2X2_475 ( .A(_abc_44694_new_n1491_), .B(_abc_44694_new_n1492_), .Y(_abc_44694_new_n1493_));
AND2X2 AND2X2_4750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7844_));
AND2X2 AND2X2_4751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7845_));
AND2X2 AND2X2_4752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7851_));
AND2X2 AND2X2_4753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7852_));
AND2X2 AND2X2_4754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7854_));
AND2X2 AND2X2_4755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7855_));
AND2X2 AND2X2_4756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7858_));
AND2X2 AND2X2_4757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7859_));
AND2X2 AND2X2_4758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7861_));
AND2X2 AND2X2_4759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7862_));
AND2X2 AND2X2_476 ( .A(_abc_44694_new_n1495_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n1496_));
AND2X2 AND2X2_4760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7866_));
AND2X2 AND2X2_4761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7867_));
AND2X2 AND2X2_4762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7868_));
AND2X2 AND2X2_4763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7871_));
AND2X2 AND2X2_4764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7872_));
AND2X2 AND2X2_4765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7874_));
AND2X2 AND2X2_4766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7875_));
AND2X2 AND2X2_4767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7880_));
AND2X2 AND2X2_4768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7881_));
AND2X2 AND2X2_4769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7883_));
AND2X2 AND2X2_477 ( .A(_abc_44694_new_n1494_), .B(_abc_44694_new_n1496_), .Y(_0epc_q_31_0__4_));
AND2X2 AND2X2_4770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7884_));
AND2X2 AND2X2_4771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7887_));
AND2X2 AND2X2_4772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7888_));
AND2X2 AND2X2_4773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7890_));
AND2X2 AND2X2_4774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7891_));
AND2X2 AND2X2_4775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7895_));
AND2X2 AND2X2_4776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7896_));
AND2X2 AND2X2_4777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7898_));
AND2X2 AND2X2_4778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7899_));
AND2X2 AND2X2_4779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7902_));
AND2X2 AND2X2_478 ( .A(_abc_44694_new_n1484_), .B(pc_q_5_), .Y(_abc_44694_new_n1499_));
AND2X2 AND2X2_4780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7903_));
AND2X2 AND2X2_4781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7905_));
AND2X2 AND2X2_4782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7906_));
AND2X2 AND2X2_4783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7912_));
AND2X2 AND2X2_4784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7913_));
AND2X2 AND2X2_4785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7915_));
AND2X2 AND2X2_4786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7916_));
AND2X2 AND2X2_4787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7919_));
AND2X2 AND2X2_4788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7920_));
AND2X2 AND2X2_4789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7922_));
AND2X2 AND2X2_479 ( .A(_abc_44694_new_n1500_), .B(_abc_44694_new_n1498_), .Y(_abc_44694_new_n1501_));
AND2X2 AND2X2_4790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7923_));
AND2X2 AND2X2_4791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7927_));
AND2X2 AND2X2_4792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7928_));
AND2X2 AND2X2_4793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7929_));
AND2X2 AND2X2_4794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7932_));
AND2X2 AND2X2_4795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7933_));
AND2X2 AND2X2_4796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7935_));
AND2X2 AND2X2_4797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7936_));
AND2X2 AND2X2_4798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7941_));
AND2X2 AND2X2_4799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7942_));
AND2X2 AND2X2_48 ( .A(_abc_44694_new_n671_), .B(alu_p_o_1_), .Y(_abc_44694_new_n699_));
AND2X2 AND2X2_480 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_5_), .Y(_abc_44694_new_n1503_));
AND2X2 AND2X2_4800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7944_));
AND2X2 AND2X2_4801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7945_));
AND2X2 AND2X2_4802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7948_));
AND2X2 AND2X2_4803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7949_));
AND2X2 AND2X2_4804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7951_));
AND2X2 AND2X2_4805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7952_));
AND2X2 AND2X2_4806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7956_));
AND2X2 AND2X2_4807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7957_));
AND2X2 AND2X2_4808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7959_));
AND2X2 AND2X2_4809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7960_));
AND2X2 AND2X2_481 ( .A(alu_op_r_3_), .B(pc_q_5_), .Y(_abc_44694_new_n1505_));
AND2X2 AND2X2_4810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7963_));
AND2X2 AND2X2_4811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7964_));
AND2X2 AND2X2_4812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7966_));
AND2X2 AND2X2_4813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7967_));
AND2X2 AND2X2_4814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7973_));
AND2X2 AND2X2_4815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7974_));
AND2X2 AND2X2_4816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7976_));
AND2X2 AND2X2_4817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7977_));
AND2X2 AND2X2_4818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7980_));
AND2X2 AND2X2_4819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7981_));
AND2X2 AND2X2_482 ( .A(_abc_44694_new_n1506_), .B(_abc_44694_new_n1504_), .Y(_abc_44694_new_n1507_));
AND2X2 AND2X2_4820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7983_));
AND2X2 AND2X2_4821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7984_));
AND2X2 AND2X2_4822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7988_));
AND2X2 AND2X2_4823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7989_));
AND2X2 AND2X2_4824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7990_));
AND2X2 AND2X2_4825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7993_));
AND2X2 AND2X2_4826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7994_));
AND2X2 AND2X2_4827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7996_));
AND2X2 AND2X2_4828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7997_));
AND2X2 AND2X2_4829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8002_));
AND2X2 AND2X2_483 ( .A(_abc_44694_new_n1472_), .B(_abc_44694_new_n1469_), .Y(_abc_44694_new_n1509_));
AND2X2 AND2X2_4830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8003_));
AND2X2 AND2X2_4831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8005_));
AND2X2 AND2X2_4832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8006_));
AND2X2 AND2X2_4833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8009_));
AND2X2 AND2X2_4834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8010_));
AND2X2 AND2X2_4835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8012_));
AND2X2 AND2X2_4836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8013_));
AND2X2 AND2X2_4837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8017_));
AND2X2 AND2X2_4838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8018_));
AND2X2 AND2X2_4839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8020_));
AND2X2 AND2X2_484 ( .A(_abc_44694_new_n1510_), .B(_abc_44694_new_n1508_), .Y(_abc_44694_new_n1511_));
AND2X2 AND2X2_4840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8021_));
AND2X2 AND2X2_4841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8024_));
AND2X2 AND2X2_4842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8025_));
AND2X2 AND2X2_4843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8027_));
AND2X2 AND2X2_4844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8028_));
AND2X2 AND2X2_4845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8034_));
AND2X2 AND2X2_4846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8035_));
AND2X2 AND2X2_4847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8037_));
AND2X2 AND2X2_4848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8038_));
AND2X2 AND2X2_4849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8041_));
AND2X2 AND2X2_485 ( .A(_abc_44694_new_n1509_), .B(_abc_44694_new_n1507_), .Y(_abc_44694_new_n1512_));
AND2X2 AND2X2_4850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8042_));
AND2X2 AND2X2_4851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8044_));
AND2X2 AND2X2_4852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8045_));
AND2X2 AND2X2_4853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8049_));
AND2X2 AND2X2_4854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8050_));
AND2X2 AND2X2_4855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8051_));
AND2X2 AND2X2_4856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8054_));
AND2X2 AND2X2_4857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8055_));
AND2X2 AND2X2_4858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8057_));
AND2X2 AND2X2_4859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8058_));
AND2X2 AND2X2_486 ( .A(_abc_44694_new_n1513_), .B(_abc_44694_new_n1194__bF_buf2), .Y(_abc_44694_new_n1514_));
AND2X2 AND2X2_4860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8063_));
AND2X2 AND2X2_4861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8064_));
AND2X2 AND2X2_4862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8066_));
AND2X2 AND2X2_4863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8067_));
AND2X2 AND2X2_4864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8070_));
AND2X2 AND2X2_4865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8071_));
AND2X2 AND2X2_4866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8073_));
AND2X2 AND2X2_4867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8074_));
AND2X2 AND2X2_4868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8078_));
AND2X2 AND2X2_4869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8079_));
AND2X2 AND2X2_487 ( .A(_abc_44694_new_n1515_), .B(_abc_44694_new_n1340__bF_buf4), .Y(_abc_44694_new_n1516_));
AND2X2 AND2X2_4870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8081_));
AND2X2 AND2X2_4871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8082_));
AND2X2 AND2X2_4872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8085_));
AND2X2 AND2X2_4873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8086_));
AND2X2 AND2X2_4874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8088_));
AND2X2 AND2X2_4875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8089_));
AND2X2 AND2X2_4876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8095_));
AND2X2 AND2X2_4877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8096_));
AND2X2 AND2X2_4878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8098_));
AND2X2 AND2X2_4879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8099_));
AND2X2 AND2X2_488 ( .A(_abc_44694_new_n1337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n1517_));
AND2X2 AND2X2_4880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8102_));
AND2X2 AND2X2_4881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8103_));
AND2X2 AND2X2_4882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8105_));
AND2X2 AND2X2_4883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8106_));
AND2X2 AND2X2_4884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8110_));
AND2X2 AND2X2_4885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8111_));
AND2X2 AND2X2_4886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8112_));
AND2X2 AND2X2_4887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8115_));
AND2X2 AND2X2_4888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8116_));
AND2X2 AND2X2_4889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8118_));
AND2X2 AND2X2_489 ( .A(_abc_44694_new_n1519_), .B(_abc_44694_new_n1502_), .Y(_abc_44694_new_n1520_));
AND2X2 AND2X2_4890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8119_));
AND2X2 AND2X2_4891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8124_));
AND2X2 AND2X2_4892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8125_));
AND2X2 AND2X2_4893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8127_));
AND2X2 AND2X2_4894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8128_));
AND2X2 AND2X2_4895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8131_));
AND2X2 AND2X2_4896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8132_));
AND2X2 AND2X2_4897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8134_));
AND2X2 AND2X2_4898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8135_));
AND2X2 AND2X2_4899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8139_));
AND2X2 AND2X2_49 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[1] ), .Y(_abc_44694_new_n700_));
AND2X2 AND2X2_490 ( .A(_abc_44694_new_n1522__bF_buf4), .B(epc_q_5_), .Y(_abc_44694_new_n1523_));
AND2X2 AND2X2_4900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8140_));
AND2X2 AND2X2_4901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8142_));
AND2X2 AND2X2_4902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8143_));
AND2X2 AND2X2_4903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8146_));
AND2X2 AND2X2_4904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8147_));
AND2X2 AND2X2_4905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8149_));
AND2X2 AND2X2_4906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8150_));
AND2X2 AND2X2_4907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8156_));
AND2X2 AND2X2_4908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8157_));
AND2X2 AND2X2_4909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8159_));
AND2X2 AND2X2_491 ( .A(_abc_44694_new_n1348__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_5_), .Y(_abc_44694_new_n1524_));
AND2X2 AND2X2_4910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8160_));
AND2X2 AND2X2_4911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8163_));
AND2X2 AND2X2_4912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8164_));
AND2X2 AND2X2_4913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8166_));
AND2X2 AND2X2_4914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8167_));
AND2X2 AND2X2_4915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8171_));
AND2X2 AND2X2_4916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8172_));
AND2X2 AND2X2_4917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8173_));
AND2X2 AND2X2_4918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8176_));
AND2X2 AND2X2_4919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8177_));
AND2X2 AND2X2_492 ( .A(_abc_44694_new_n1521_), .B(_abc_44694_new_n1526_), .Y(_abc_44694_new_n1527_));
AND2X2 AND2X2_4920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8179_));
AND2X2 AND2X2_4921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8180_));
AND2X2 AND2X2_4922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8185_));
AND2X2 AND2X2_4923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8186_));
AND2X2 AND2X2_4924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8188_));
AND2X2 AND2X2_4925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8189_));
AND2X2 AND2X2_4926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8192_));
AND2X2 AND2X2_4927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8193_));
AND2X2 AND2X2_4928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8195_));
AND2X2 AND2X2_4929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8196_));
AND2X2 AND2X2_493 ( .A(_abc_44694_new_n1528_), .B(_abc_44694_new_n1529_), .Y(_abc_44694_new_n1530_));
AND2X2 AND2X2_4930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8200_));
AND2X2 AND2X2_4931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8201_));
AND2X2 AND2X2_4932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8203_));
AND2X2 AND2X2_4933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8204_));
AND2X2 AND2X2_4934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8207_));
AND2X2 AND2X2_4935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8208_));
AND2X2 AND2X2_4936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8210_));
AND2X2 AND2X2_4937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8211_));
AND2X2 AND2X2_4938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8217_));
AND2X2 AND2X2_4939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8218_));
AND2X2 AND2X2_494 ( .A(_abc_44694_new_n1532_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n1533_));
AND2X2 AND2X2_4940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8220_));
AND2X2 AND2X2_4941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8221_));
AND2X2 AND2X2_4942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8224_));
AND2X2 AND2X2_4943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8225_));
AND2X2 AND2X2_4944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8227_));
AND2X2 AND2X2_4945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8228_));
AND2X2 AND2X2_4946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8232_));
AND2X2 AND2X2_4947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8233_));
AND2X2 AND2X2_4948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8234_));
AND2X2 AND2X2_4949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8237_));
AND2X2 AND2X2_495 ( .A(_abc_44694_new_n1531_), .B(_abc_44694_new_n1533_), .Y(_0epc_q_31_0__5_));
AND2X2 AND2X2_4950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8238_));
AND2X2 AND2X2_4951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8240_));
AND2X2 AND2X2_4952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8241_));
AND2X2 AND2X2_4953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8246_));
AND2X2 AND2X2_4954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8247_));
AND2X2 AND2X2_4955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8249_));
AND2X2 AND2X2_4956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8250_));
AND2X2 AND2X2_4957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8253_));
AND2X2 AND2X2_4958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8254_));
AND2X2 AND2X2_4959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8256_));
AND2X2 AND2X2_496 ( .A(_abc_44694_new_n1499_), .B(pc_q_6_), .Y(_abc_44694_new_n1537_));
AND2X2 AND2X2_4960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8257_));
AND2X2 AND2X2_4961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8261_));
AND2X2 AND2X2_4962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8262_));
AND2X2 AND2X2_4963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8264_));
AND2X2 AND2X2_4964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8265_));
AND2X2 AND2X2_4965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8268_));
AND2X2 AND2X2_4966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8269_));
AND2X2 AND2X2_4967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8271_));
AND2X2 AND2X2_4968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8272_));
AND2X2 AND2X2_4969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8278_));
AND2X2 AND2X2_497 ( .A(_abc_44694_new_n1538_), .B(_abc_44694_new_n1536_), .Y(_abc_44694_new_n1539_));
AND2X2 AND2X2_4970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8279_));
AND2X2 AND2X2_4971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8281_));
AND2X2 AND2X2_4972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8282_));
AND2X2 AND2X2_4973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8285_));
AND2X2 AND2X2_4974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8286_));
AND2X2 AND2X2_4975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8288_));
AND2X2 AND2X2_4976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8289_));
AND2X2 AND2X2_4977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8293_));
AND2X2 AND2X2_4978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8294_));
AND2X2 AND2X2_4979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8295_));
AND2X2 AND2X2_498 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1540_), .Y(_abc_44694_new_n1541_));
AND2X2 AND2X2_4980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8298_));
AND2X2 AND2X2_4981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8299_));
AND2X2 AND2X2_4982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8301_));
AND2X2 AND2X2_4983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8302_));
AND2X2 AND2X2_4984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8307_));
AND2X2 AND2X2_4985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8308_));
AND2X2 AND2X2_4986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8310_));
AND2X2 AND2X2_4987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8311_));
AND2X2 AND2X2_4988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8314_));
AND2X2 AND2X2_4989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8315_));
AND2X2 AND2X2_499 ( .A(_abc_44694_new_n1019__bF_buf4), .B(epc_q_6_), .Y(_abc_44694_new_n1543_));
AND2X2 AND2X2_4990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8317_));
AND2X2 AND2X2_4991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8318_));
AND2X2 AND2X2_4992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8322_));
AND2X2 AND2X2_4993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8323_));
AND2X2 AND2X2_4994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8325_));
AND2X2 AND2X2_4995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8326_));
AND2X2 AND2X2_4996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8329_));
AND2X2 AND2X2_4997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8330_));
AND2X2 AND2X2_4998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8332_));
AND2X2 AND2X2_4999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8333_));
AND2X2 AND2X2_5 ( .A(_abc_44694_new_n626_), .B(_abc_44694_new_n623_), .Y(_abc_44694_new_n627_));
AND2X2 AND2X2_50 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[17] ), .Y(_abc_44694_new_n701_));
AND2X2 AND2X2_500 ( .A(_abc_44694_new_n1470_), .B(_abc_44694_new_n1507_), .Y(_abc_44694_new_n1544_));
AND2X2 AND2X2_5000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8339_));
AND2X2 AND2X2_5001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8340_));
AND2X2 AND2X2_5002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8342_));
AND2X2 AND2X2_5003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8343_));
AND2X2 AND2X2_5004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8346_));
AND2X2 AND2X2_5005 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8347_));
AND2X2 AND2X2_5006 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8349_));
AND2X2 AND2X2_5007 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8350_));
AND2X2 AND2X2_5008 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8354_));
AND2X2 AND2X2_5009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8355_));
AND2X2 AND2X2_501 ( .A(_abc_44694_new_n1473_), .B(_abc_44694_new_n1544_), .Y(_abc_44694_new_n1545_));
AND2X2 AND2X2_5010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8356_));
AND2X2 AND2X2_5011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8359_));
AND2X2 AND2X2_5012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8360_));
AND2X2 AND2X2_5013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8362_));
AND2X2 AND2X2_5014 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8363_));
AND2X2 AND2X2_5015 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8368_));
AND2X2 AND2X2_5016 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8369_));
AND2X2 AND2X2_5017 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8371_));
AND2X2 AND2X2_5018 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8372_));
AND2X2 AND2X2_5019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8375_));
AND2X2 AND2X2_502 ( .A(_abc_44694_new_n1507_), .B(_abc_44694_new_n1468_), .Y(_abc_44694_new_n1546_));
AND2X2 AND2X2_5020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8376_));
AND2X2 AND2X2_5021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8378_));
AND2X2 AND2X2_5022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8379_));
AND2X2 AND2X2_5023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8383_));
AND2X2 AND2X2_5024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8384_));
AND2X2 AND2X2_5025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8386_));
AND2X2 AND2X2_5026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8387_));
AND2X2 AND2X2_5027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8390_));
AND2X2 AND2X2_5028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8391_));
AND2X2 AND2X2_5029 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8393_));
AND2X2 AND2X2_503 ( .A(int32_r_4_), .B(pc_q_6_), .Y(_abc_44694_new_n1550_));
AND2X2 AND2X2_5030 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8394_));
AND2X2 AND2X2_5031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8400_));
AND2X2 AND2X2_5032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8401_));
AND2X2 AND2X2_5033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8403_));
AND2X2 AND2X2_5034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8404_));
AND2X2 AND2X2_5035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8407_));
AND2X2 AND2X2_5036 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8408_));
AND2X2 AND2X2_5037 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8410_));
AND2X2 AND2X2_5038 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8411_));
AND2X2 AND2X2_5039 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8415_));
AND2X2 AND2X2_504 ( .A(_abc_44694_new_n1551_), .B(_abc_44694_new_n1549_), .Y(_abc_44694_new_n1552_));
AND2X2 AND2X2_5040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8416_));
AND2X2 AND2X2_5041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8417_));
AND2X2 AND2X2_5042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8420_));
AND2X2 AND2X2_5043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8421_));
AND2X2 AND2X2_5044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8423_));
AND2X2 AND2X2_5045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8424_));
AND2X2 AND2X2_5046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8429_));
AND2X2 AND2X2_5047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8430_));
AND2X2 AND2X2_5048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8432_));
AND2X2 AND2X2_5049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8433_));
AND2X2 AND2X2_505 ( .A(_abc_44694_new_n1548_), .B(_abc_44694_new_n1552_), .Y(_abc_44694_new_n1554_));
AND2X2 AND2X2_5050 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8436_));
AND2X2 AND2X2_5051 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8437_));
AND2X2 AND2X2_5052 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8439_));
AND2X2 AND2X2_5053 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8440_));
AND2X2 AND2X2_5054 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8444_));
AND2X2 AND2X2_5055 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8445_));
AND2X2 AND2X2_5056 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8447_));
AND2X2 AND2X2_5057 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8448_));
AND2X2 AND2X2_5058 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8451_));
AND2X2 AND2X2_5059 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8452_));
AND2X2 AND2X2_506 ( .A(_abc_44694_new_n1555_), .B(_abc_44694_new_n1194__bF_buf1), .Y(_abc_44694_new_n1556_));
AND2X2 AND2X2_5060 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8454_));
AND2X2 AND2X2_5061 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8455_));
AND2X2 AND2X2_5062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8461_));
AND2X2 AND2X2_5063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8462_));
AND2X2 AND2X2_5064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8464_));
AND2X2 AND2X2_5065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8465_));
AND2X2 AND2X2_5066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8468_));
AND2X2 AND2X2_5067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8469_));
AND2X2 AND2X2_5068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8471_));
AND2X2 AND2X2_5069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8472_));
AND2X2 AND2X2_507 ( .A(_abc_44694_new_n1556_), .B(_abc_44694_new_n1553_), .Y(_abc_44694_new_n1557_));
AND2X2 AND2X2_5070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8476_));
AND2X2 AND2X2_5071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8477_));
AND2X2 AND2X2_5072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8478_));
AND2X2 AND2X2_5073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8481_));
AND2X2 AND2X2_5074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8482_));
AND2X2 AND2X2_5075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8484_));
AND2X2 AND2X2_5076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8485_));
AND2X2 AND2X2_5077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8490_));
AND2X2 AND2X2_5078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8491_));
AND2X2 AND2X2_5079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8493_));
AND2X2 AND2X2_508 ( .A(_abc_44694_new_n1558_), .B(_abc_44694_new_n1340__bF_buf3), .Y(_abc_44694_new_n1559_));
AND2X2 AND2X2_5080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8494_));
AND2X2 AND2X2_5081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8497_));
AND2X2 AND2X2_5082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8498_));
AND2X2 AND2X2_5083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8500_));
AND2X2 AND2X2_5084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8501_));
AND2X2 AND2X2_5085 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8505_));
AND2X2 AND2X2_5086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8506_));
AND2X2 AND2X2_5087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8508_));
AND2X2 AND2X2_5088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8509_));
AND2X2 AND2X2_5089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8512_));
AND2X2 AND2X2_509 ( .A(_abc_44694_new_n1337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n1560_));
AND2X2 AND2X2_5090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8513_));
AND2X2 AND2X2_5091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8515_));
AND2X2 AND2X2_5092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8516_));
AND2X2 AND2X2_5093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8522_));
AND2X2 AND2X2_5094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8523_));
AND2X2 AND2X2_5095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8525_));
AND2X2 AND2X2_5096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8526_));
AND2X2 AND2X2_5097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8529_));
AND2X2 AND2X2_5098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8530_));
AND2X2 AND2X2_5099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8532_));
AND2X2 AND2X2_51 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[17] ), .Y(_abc_44694_new_n704_));
AND2X2 AND2X2_510 ( .A(_abc_44694_new_n1562_), .B(_abc_44694_new_n1542_), .Y(_abc_44694_new_n1563_));
AND2X2 AND2X2_5100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8533_));
AND2X2 AND2X2_5101 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8537_));
AND2X2 AND2X2_5102 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8538_));
AND2X2 AND2X2_5103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8539_));
AND2X2 AND2X2_5104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8542_));
AND2X2 AND2X2_5105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8543_));
AND2X2 AND2X2_5106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8545_));
AND2X2 AND2X2_5107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8546_));
AND2X2 AND2X2_5108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8551_));
AND2X2 AND2X2_5109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8552_));
AND2X2 AND2X2_511 ( .A(_abc_44694_new_n1522__bF_buf3), .B(epc_q_6_), .Y(_abc_44694_new_n1565_));
AND2X2 AND2X2_5110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8554_));
AND2X2 AND2X2_5111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8555_));
AND2X2 AND2X2_5112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8558_));
AND2X2 AND2X2_5113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8559_));
AND2X2 AND2X2_5114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8561_));
AND2X2 AND2X2_5115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8562_));
AND2X2 AND2X2_5116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8566_));
AND2X2 AND2X2_5117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8567_));
AND2X2 AND2X2_5118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8569_));
AND2X2 AND2X2_5119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8570_));
AND2X2 AND2X2_512 ( .A(_abc_44694_new_n1348__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_6_), .Y(_abc_44694_new_n1566_));
AND2X2 AND2X2_5120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8573_));
AND2X2 AND2X2_5121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8574_));
AND2X2 AND2X2_5122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8576_));
AND2X2 AND2X2_5123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8577_));
AND2X2 AND2X2_5124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8583_));
AND2X2 AND2X2_5125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8584_));
AND2X2 AND2X2_5126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8586_));
AND2X2 AND2X2_5127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8587_));
AND2X2 AND2X2_5128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8590_));
AND2X2 AND2X2_5129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8591_));
AND2X2 AND2X2_513 ( .A(_abc_44694_new_n1207__bF_buf1), .B(_abc_44694_new_n1568_), .Y(_abc_44694_new_n1569_));
AND2X2 AND2X2_5130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8593_));
AND2X2 AND2X2_5131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8594_));
AND2X2 AND2X2_5132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8598_));
AND2X2 AND2X2_5133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8599_));
AND2X2 AND2X2_5134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8600_));
AND2X2 AND2X2_5135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8603_));
AND2X2 AND2X2_5136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8604_));
AND2X2 AND2X2_5137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8606_));
AND2X2 AND2X2_5138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8607_));
AND2X2 AND2X2_5139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8612_));
AND2X2 AND2X2_514 ( .A(_abc_44694_new_n1569_), .B(_abc_44694_new_n1564_), .Y(_abc_44694_new_n1570_));
AND2X2 AND2X2_5140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8613_));
AND2X2 AND2X2_5141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8615_));
AND2X2 AND2X2_5142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8616_));
AND2X2 AND2X2_5143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8619_));
AND2X2 AND2X2_5144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8620_));
AND2X2 AND2X2_5145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8622_));
AND2X2 AND2X2_5146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8623_));
AND2X2 AND2X2_5147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8627_));
AND2X2 AND2X2_5148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8628_));
AND2X2 AND2X2_5149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8630_));
AND2X2 AND2X2_515 ( .A(_abc_44694_new_n1572_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n1573_));
AND2X2 AND2X2_5150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8631_));
AND2X2 AND2X2_5151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8634_));
AND2X2 AND2X2_5152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8635_));
AND2X2 AND2X2_5153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8637_));
AND2X2 AND2X2_5154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8638_));
AND2X2 AND2X2_5155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8644_));
AND2X2 AND2X2_5156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8645_));
AND2X2 AND2X2_5157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8647_));
AND2X2 AND2X2_5158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8648_));
AND2X2 AND2X2_5159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8651_));
AND2X2 AND2X2_516 ( .A(_abc_44694_new_n1571_), .B(_abc_44694_new_n1573_), .Y(_0epc_q_31_0__6_));
AND2X2 AND2X2_5160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8652_));
AND2X2 AND2X2_5161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8654_));
AND2X2 AND2X2_5162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8655_));
AND2X2 AND2X2_5163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8659_));
AND2X2 AND2X2_5164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8660_));
AND2X2 AND2X2_5165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8661_));
AND2X2 AND2X2_5166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8664_));
AND2X2 AND2X2_5167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8665_));
AND2X2 AND2X2_5168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8667_));
AND2X2 AND2X2_5169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8668_));
AND2X2 AND2X2_517 ( .A(_abc_44694_new_n1537_), .B(pc_q_7_), .Y(_abc_44694_new_n1576_));
AND2X2 AND2X2_5170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8673_));
AND2X2 AND2X2_5171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8674_));
AND2X2 AND2X2_5172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8676_));
AND2X2 AND2X2_5173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8677_));
AND2X2 AND2X2_5174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8680_));
AND2X2 AND2X2_5175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8681_));
AND2X2 AND2X2_5176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8683_));
AND2X2 AND2X2_5177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8684_));
AND2X2 AND2X2_5178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8688_));
AND2X2 AND2X2_5179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8689_));
AND2X2 AND2X2_518 ( .A(_abc_44694_new_n1577_), .B(_abc_44694_new_n1575_), .Y(_abc_44694_new_n1578_));
AND2X2 AND2X2_5180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8691_));
AND2X2 AND2X2_5181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8692_));
AND2X2 AND2X2_5182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8695_));
AND2X2 AND2X2_5183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8696_));
AND2X2 AND2X2_5184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8698_));
AND2X2 AND2X2_5185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8699_));
AND2X2 AND2X2_5186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8705_));
AND2X2 AND2X2_5187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8706_));
AND2X2 AND2X2_5188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8708_));
AND2X2 AND2X2_5189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8709_));
AND2X2 AND2X2_519 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1579_), .Y(_abc_44694_new_n1580_));
AND2X2 AND2X2_5190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8712_));
AND2X2 AND2X2_5191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8713_));
AND2X2 AND2X2_5192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8715_));
AND2X2 AND2X2_5193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8716_));
AND2X2 AND2X2_5194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8720_));
AND2X2 AND2X2_5195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8721_));
AND2X2 AND2X2_5196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8722_));
AND2X2 AND2X2_5197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8725_));
AND2X2 AND2X2_5198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8726_));
AND2X2 AND2X2_5199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8728_));
AND2X2 AND2X2_52 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[9] ), .Y(_abc_44694_new_n705_));
AND2X2 AND2X2_520 ( .A(_abc_44694_new_n1019__bF_buf3), .B(epc_q_7_), .Y(_abc_44694_new_n1582_));
AND2X2 AND2X2_5200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8729_));
AND2X2 AND2X2_5201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8734_));
AND2X2 AND2X2_5202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8735_));
AND2X2 AND2X2_5203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8737_));
AND2X2 AND2X2_5204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8738_));
AND2X2 AND2X2_5205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8741_));
AND2X2 AND2X2_5206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8742_));
AND2X2 AND2X2_5207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8744_));
AND2X2 AND2X2_5208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8745_));
AND2X2 AND2X2_5209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8749_));
AND2X2 AND2X2_521 ( .A(int32_r_5_), .B(pc_q_7_), .Y(_abc_44694_new_n1584_));
AND2X2 AND2X2_5210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8750_));
AND2X2 AND2X2_5211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8752_));
AND2X2 AND2X2_5212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8753_));
AND2X2 AND2X2_5213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8756_));
AND2X2 AND2X2_5214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8757_));
AND2X2 AND2X2_5215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8759_));
AND2X2 AND2X2_5216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8760_));
AND2X2 AND2X2_5217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8766_));
AND2X2 AND2X2_5218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8767_));
AND2X2 AND2X2_5219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8769_));
AND2X2 AND2X2_522 ( .A(_abc_44694_new_n1585_), .B(_abc_44694_new_n1583_), .Y(_abc_44694_new_n1586_));
AND2X2 AND2X2_5220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8770_));
AND2X2 AND2X2_5221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8773_));
AND2X2 AND2X2_5222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8774_));
AND2X2 AND2X2_5223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8776_));
AND2X2 AND2X2_5224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8777_));
AND2X2 AND2X2_5225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8781_));
AND2X2 AND2X2_5226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8782_));
AND2X2 AND2X2_5227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8783_));
AND2X2 AND2X2_5228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8786_));
AND2X2 AND2X2_5229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8787_));
AND2X2 AND2X2_523 ( .A(_abc_44694_new_n1552_), .B(_abc_44694_new_n1586_), .Y(_abc_44694_new_n1589_));
AND2X2 AND2X2_5230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8789_));
AND2X2 AND2X2_5231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8790_));
AND2X2 AND2X2_5232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8795_));
AND2X2 AND2X2_5233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8796_));
AND2X2 AND2X2_5234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8798_));
AND2X2 AND2X2_5235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8799_));
AND2X2 AND2X2_5236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8802_));
AND2X2 AND2X2_5237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8803_));
AND2X2 AND2X2_5238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8805_));
AND2X2 AND2X2_5239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8806_));
AND2X2 AND2X2_524 ( .A(_abc_44694_new_n1548_), .B(_abc_44694_new_n1589_), .Y(_abc_44694_new_n1590_));
AND2X2 AND2X2_5240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8810_));
AND2X2 AND2X2_5241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8811_));
AND2X2 AND2X2_5242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8813_));
AND2X2 AND2X2_5243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8814_));
AND2X2 AND2X2_5244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8817_));
AND2X2 AND2X2_5245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8818_));
AND2X2 AND2X2_5246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8820_));
AND2X2 AND2X2_5247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8821_));
AND2X2 AND2X2_5248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8827_));
AND2X2 AND2X2_5249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8828_));
AND2X2 AND2X2_525 ( .A(_abc_44694_new_n1586_), .B(_abc_44694_new_n1550_), .Y(_abc_44694_new_n1592_));
AND2X2 AND2X2_5250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8830_));
AND2X2 AND2X2_5251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8831_));
AND2X2 AND2X2_5252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8834_));
AND2X2 AND2X2_5253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8835_));
AND2X2 AND2X2_5254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8837_));
AND2X2 AND2X2_5255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8838_));
AND2X2 AND2X2_5256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8842_));
AND2X2 AND2X2_5257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8843_));
AND2X2 AND2X2_5258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8844_));
AND2X2 AND2X2_5259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8847_));
AND2X2 AND2X2_526 ( .A(_abc_44694_new_n1194__bF_buf0), .B(_abc_44694_new_n1593_), .Y(_abc_44694_new_n1594_));
AND2X2 AND2X2_5260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8848_));
AND2X2 AND2X2_5261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8850_));
AND2X2 AND2X2_5262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8851_));
AND2X2 AND2X2_5263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8856_));
AND2X2 AND2X2_5264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8857_));
AND2X2 AND2X2_5265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8859_));
AND2X2 AND2X2_5266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8860_));
AND2X2 AND2X2_5267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8863_));
AND2X2 AND2X2_5268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8864_));
AND2X2 AND2X2_5269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8866_));
AND2X2 AND2X2_527 ( .A(_abc_44694_new_n1591_), .B(_abc_44694_new_n1594_), .Y(_abc_44694_new_n1595_));
AND2X2 AND2X2_5270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8867_));
AND2X2 AND2X2_5271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8871_));
AND2X2 AND2X2_5272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8872_));
AND2X2 AND2X2_5273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8874_));
AND2X2 AND2X2_5274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8875_));
AND2X2 AND2X2_5275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8878_));
AND2X2 AND2X2_5276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8879_));
AND2X2 AND2X2_5277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8881_));
AND2X2 AND2X2_5278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8882_));
AND2X2 AND2X2_5279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8888_));
AND2X2 AND2X2_528 ( .A(_abc_44694_new_n1595_), .B(_abc_44694_new_n1588_), .Y(_abc_44694_new_n1596_));
AND2X2 AND2X2_5280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8889_));
AND2X2 AND2X2_5281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8891_));
AND2X2 AND2X2_5282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8892_));
AND2X2 AND2X2_5283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8895_));
AND2X2 AND2X2_5284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8896_));
AND2X2 AND2X2_5285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8898_));
AND2X2 AND2X2_5286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8899_));
AND2X2 AND2X2_5287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8903_));
AND2X2 AND2X2_5288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8904_));
AND2X2 AND2X2_5289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8905_));
AND2X2 AND2X2_529 ( .A(_abc_44694_new_n1597_), .B(_abc_44694_new_n1340__bF_buf2), .Y(_abc_44694_new_n1598_));
AND2X2 AND2X2_5290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8908_));
AND2X2 AND2X2_5291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8909_));
AND2X2 AND2X2_5292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8911_));
AND2X2 AND2X2_5293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8912_));
AND2X2 AND2X2_5294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8917_));
AND2X2 AND2X2_5295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8918_));
AND2X2 AND2X2_5296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8920_));
AND2X2 AND2X2_5297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8921_));
AND2X2 AND2X2_5298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8924_));
AND2X2 AND2X2_5299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8925_));
AND2X2 AND2X2_53 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[25] ), .Y(_abc_44694_new_n707_));
AND2X2 AND2X2_530 ( .A(_abc_44694_new_n1337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n1599_));
AND2X2 AND2X2_5300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8927_));
AND2X2 AND2X2_5301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8928_));
AND2X2 AND2X2_5302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8932_));
AND2X2 AND2X2_5303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8933_));
AND2X2 AND2X2_5304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8935_));
AND2X2 AND2X2_5305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8936_));
AND2X2 AND2X2_5306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8939_));
AND2X2 AND2X2_5307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8940_));
AND2X2 AND2X2_5308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8942_));
AND2X2 AND2X2_5309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8943_));
AND2X2 AND2X2_531 ( .A(_abc_44694_new_n1601_), .B(_abc_44694_new_n1581_), .Y(_abc_44694_new_n1602_));
AND2X2 AND2X2_5310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8949_));
AND2X2 AND2X2_5311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8950_));
AND2X2 AND2X2_5312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8952_));
AND2X2 AND2X2_5313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8953_));
AND2X2 AND2X2_5314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8956_));
AND2X2 AND2X2_5315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8957_));
AND2X2 AND2X2_5316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8959_));
AND2X2 AND2X2_5317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8960_));
AND2X2 AND2X2_5318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8964_));
AND2X2 AND2X2_5319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8965_));
AND2X2 AND2X2_532 ( .A(_abc_44694_new_n1522__bF_buf2), .B(epc_q_7_), .Y(_abc_44694_new_n1604_));
AND2X2 AND2X2_5320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8966_));
AND2X2 AND2X2_5321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8969_));
AND2X2 AND2X2_5322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8970_));
AND2X2 AND2X2_5323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8972_));
AND2X2 AND2X2_5324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8973_));
AND2X2 AND2X2_5325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8978_));
AND2X2 AND2X2_5326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8979_));
AND2X2 AND2X2_5327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8981_));
AND2X2 AND2X2_5328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8982_));
AND2X2 AND2X2_5329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8985_));
AND2X2 AND2X2_533 ( .A(_abc_44694_new_n1348__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_7_), .Y(_abc_44694_new_n1605_));
AND2X2 AND2X2_5330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8986_));
AND2X2 AND2X2_5331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8988_));
AND2X2 AND2X2_5332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8989_));
AND2X2 AND2X2_5333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8993_));
AND2X2 AND2X2_5334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8994_));
AND2X2 AND2X2_5335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8996_));
AND2X2 AND2X2_5336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8997_));
AND2X2 AND2X2_5337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9000_));
AND2X2 AND2X2_5338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9001_));
AND2X2 AND2X2_5339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9003_));
AND2X2 AND2X2_534 ( .A(_abc_44694_new_n1207__bF_buf0), .B(_abc_44694_new_n1607_), .Y(_abc_44694_new_n1608_));
AND2X2 AND2X2_5340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9004_));
AND2X2 AND2X2_5341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9010_));
AND2X2 AND2X2_5342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9011_));
AND2X2 AND2X2_5343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9013_));
AND2X2 AND2X2_5344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9014_));
AND2X2 AND2X2_5345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9017_));
AND2X2 AND2X2_5346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9018_));
AND2X2 AND2X2_5347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9020_));
AND2X2 AND2X2_5348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9021_));
AND2X2 AND2X2_5349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9025_));
AND2X2 AND2X2_535 ( .A(_abc_44694_new_n1608_), .B(_abc_44694_new_n1603_), .Y(_abc_44694_new_n1609_));
AND2X2 AND2X2_5350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9026_));
AND2X2 AND2X2_5351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9027_));
AND2X2 AND2X2_5352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9030_));
AND2X2 AND2X2_5353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9031_));
AND2X2 AND2X2_5354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9033_));
AND2X2 AND2X2_5355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9034_));
AND2X2 AND2X2_5356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9039_));
AND2X2 AND2X2_5357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9040_));
AND2X2 AND2X2_5358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9042_));
AND2X2 AND2X2_5359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9043_));
AND2X2 AND2X2_536 ( .A(_abc_44694_new_n1611_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n1612_));
AND2X2 AND2X2_5360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9046_));
AND2X2 AND2X2_5361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9047_));
AND2X2 AND2X2_5362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9049_));
AND2X2 AND2X2_5363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9050_));
AND2X2 AND2X2_5364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9054_));
AND2X2 AND2X2_5365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9055_));
AND2X2 AND2X2_5366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9057_));
AND2X2 AND2X2_5367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9058_));
AND2X2 AND2X2_5368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9061_));
AND2X2 AND2X2_5369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9062_));
AND2X2 AND2X2_537 ( .A(_abc_44694_new_n1610_), .B(_abc_44694_new_n1612_), .Y(_0epc_q_31_0__7_));
AND2X2 AND2X2_5370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9064_));
AND2X2 AND2X2_5371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9065_));
AND2X2 AND2X2_5372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9071_));
AND2X2 AND2X2_5373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9072_));
AND2X2 AND2X2_5374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9074_));
AND2X2 AND2X2_5375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9075_));
AND2X2 AND2X2_5376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9078_));
AND2X2 AND2X2_5377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9079_));
AND2X2 AND2X2_5378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9081_));
AND2X2 AND2X2_5379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9082_));
AND2X2 AND2X2_538 ( .A(_abc_44694_new_n1576_), .B(pc_q_8_), .Y(_abc_44694_new_n1615_));
AND2X2 AND2X2_5380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9086_));
AND2X2 AND2X2_5381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9087_));
AND2X2 AND2X2_5382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9088_));
AND2X2 AND2X2_5383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9091_));
AND2X2 AND2X2_5384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9092_));
AND2X2 AND2X2_5385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9094_));
AND2X2 AND2X2_5386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9095_));
AND2X2 AND2X2_5387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9100_));
AND2X2 AND2X2_5388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9101_));
AND2X2 AND2X2_5389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9103_));
AND2X2 AND2X2_539 ( .A(_abc_44694_new_n1616_), .B(_abc_44694_new_n1614_), .Y(_abc_44694_new_n1617_));
AND2X2 AND2X2_5390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9104_));
AND2X2 AND2X2_5391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9107_));
AND2X2 AND2X2_5392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9108_));
AND2X2 AND2X2_5393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9110_));
AND2X2 AND2X2_5394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9111_));
AND2X2 AND2X2_5395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9115_));
AND2X2 AND2X2_5396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9116_));
AND2X2 AND2X2_5397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9118_));
AND2X2 AND2X2_5398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9119_));
AND2X2 AND2X2_5399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9122_));
AND2X2 AND2X2_54 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[1] ), .Y(_abc_44694_new_n708_));
AND2X2 AND2X2_540 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1618_), .Y(_abc_44694_new_n1619_));
AND2X2 AND2X2_5400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9123_));
AND2X2 AND2X2_5401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9125_));
AND2X2 AND2X2_5402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9126_));
AND2X2 AND2X2_5403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9132_));
AND2X2 AND2X2_5404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9133_));
AND2X2 AND2X2_5405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9135_));
AND2X2 AND2X2_5406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9136_));
AND2X2 AND2X2_5407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9139_));
AND2X2 AND2X2_5408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9140_));
AND2X2 AND2X2_5409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9142_));
AND2X2 AND2X2_541 ( .A(_abc_44694_new_n1019__bF_buf2), .B(epc_q_8_), .Y(_abc_44694_new_n1621_));
AND2X2 AND2X2_5410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9143_));
AND2X2 AND2X2_5411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9147_));
AND2X2 AND2X2_5412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9148_));
AND2X2 AND2X2_5413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9149_));
AND2X2 AND2X2_5414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9152_));
AND2X2 AND2X2_5415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9153_));
AND2X2 AND2X2_5416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9155_));
AND2X2 AND2X2_5417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9156_));
AND2X2 AND2X2_5418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9161_));
AND2X2 AND2X2_5419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9162_));
AND2X2 AND2X2_542 ( .A(_abc_44694_new_n1593_), .B(_abc_44694_new_n1585_), .Y(_abc_44694_new_n1622_));
AND2X2 AND2X2_5420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9164_));
AND2X2 AND2X2_5421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9165_));
AND2X2 AND2X2_5422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9168_));
AND2X2 AND2X2_5423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9169_));
AND2X2 AND2X2_5424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9171_));
AND2X2 AND2X2_5425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9172_));
AND2X2 AND2X2_5426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9176_));
AND2X2 AND2X2_5427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9177_));
AND2X2 AND2X2_5428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9179_));
AND2X2 AND2X2_5429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9180_));
AND2X2 AND2X2_543 ( .A(alu_op_r_4_), .B(pc_q_8_), .Y(_abc_44694_new_n1626_));
AND2X2 AND2X2_5430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9183_));
AND2X2 AND2X2_5431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9184_));
AND2X2 AND2X2_5432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9186_));
AND2X2 AND2X2_5433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9187_));
AND2X2 AND2X2_5434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9193_));
AND2X2 AND2X2_5435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9194_));
AND2X2 AND2X2_5436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9196_));
AND2X2 AND2X2_5437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9197_));
AND2X2 AND2X2_5438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9200_));
AND2X2 AND2X2_5439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9201_));
AND2X2 AND2X2_544 ( .A(_abc_44694_new_n1627_), .B(_abc_44694_new_n1625_), .Y(_abc_44694_new_n1628_));
AND2X2 AND2X2_5440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9203_));
AND2X2 AND2X2_5441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9204_));
AND2X2 AND2X2_5442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9208_));
AND2X2 AND2X2_5443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9209_));
AND2X2 AND2X2_5444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9210_));
AND2X2 AND2X2_5445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9213_));
AND2X2 AND2X2_5446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9214_));
AND2X2 AND2X2_5447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9216_));
AND2X2 AND2X2_5448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9217_));
AND2X2 AND2X2_5449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9222_));
AND2X2 AND2X2_545 ( .A(_abc_44694_new_n1624_), .B(_abc_44694_new_n1628_), .Y(_abc_44694_new_n1630_));
AND2X2 AND2X2_5450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9223_));
AND2X2 AND2X2_5451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9225_));
AND2X2 AND2X2_5452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9226_));
AND2X2 AND2X2_5453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9229_));
AND2X2 AND2X2_5454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9230_));
AND2X2 AND2X2_5455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9232_));
AND2X2 AND2X2_5456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9233_));
AND2X2 AND2X2_5457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9237_));
AND2X2 AND2X2_5458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9238_));
AND2X2 AND2X2_5459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9240_));
AND2X2 AND2X2_546 ( .A(_abc_44694_new_n1631_), .B(_abc_44694_new_n1194__bF_buf4), .Y(_abc_44694_new_n1632_));
AND2X2 AND2X2_5460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9241_));
AND2X2 AND2X2_5461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9244_));
AND2X2 AND2X2_5462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9245_));
AND2X2 AND2X2_5463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9247_));
AND2X2 AND2X2_5464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9248_));
AND2X2 AND2X2_5465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9254_));
AND2X2 AND2X2_5466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9255_));
AND2X2 AND2X2_5467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9257_));
AND2X2 AND2X2_5468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9258_));
AND2X2 AND2X2_5469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9261_));
AND2X2 AND2X2_547 ( .A(_abc_44694_new_n1632_), .B(_abc_44694_new_n1629_), .Y(_abc_44694_new_n1633_));
AND2X2 AND2X2_5470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9262_));
AND2X2 AND2X2_5471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9264_));
AND2X2 AND2X2_5472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9265_));
AND2X2 AND2X2_5473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9269_));
AND2X2 AND2X2_5474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9270_));
AND2X2 AND2X2_5475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9271_));
AND2X2 AND2X2_5476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9274_));
AND2X2 AND2X2_5477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9275_));
AND2X2 AND2X2_5478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9277_));
AND2X2 AND2X2_5479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9278_));
AND2X2 AND2X2_548 ( .A(_abc_44694_new_n1634_), .B(_abc_44694_new_n1340__bF_buf1), .Y(_abc_44694_new_n1635_));
AND2X2 AND2X2_5480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9283_));
AND2X2 AND2X2_5481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9284_));
AND2X2 AND2X2_5482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9286_));
AND2X2 AND2X2_5483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9287_));
AND2X2 AND2X2_5484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9290_));
AND2X2 AND2X2_5485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9291_));
AND2X2 AND2X2_5486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9293_));
AND2X2 AND2X2_5487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9294_));
AND2X2 AND2X2_5488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9298_));
AND2X2 AND2X2_5489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9299_));
AND2X2 AND2X2_549 ( .A(_abc_44694_new_n1337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n1636_));
AND2X2 AND2X2_5490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9301_));
AND2X2 AND2X2_5491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9302_));
AND2X2 AND2X2_5492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9305_));
AND2X2 AND2X2_5493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9306_));
AND2X2 AND2X2_5494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9308_));
AND2X2 AND2X2_5495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9309_));
AND2X2 AND2X2_5496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9315_));
AND2X2 AND2X2_5497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9316_));
AND2X2 AND2X2_5498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9318_));
AND2X2 AND2X2_5499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9319_));
AND2X2 AND2X2_55 ( .A(_abc_44694_new_n711_), .B(state_q_1_bF_buf0_), .Y(_abc_44694_new_n712_));
AND2X2 AND2X2_550 ( .A(_abc_44694_new_n1638_), .B(_abc_44694_new_n1620_), .Y(_abc_44694_new_n1639_));
AND2X2 AND2X2_5500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9322_));
AND2X2 AND2X2_5501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9323_));
AND2X2 AND2X2_5502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9325_));
AND2X2 AND2X2_5503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9326_));
AND2X2 AND2X2_5504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9330_));
AND2X2 AND2X2_5505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9331_));
AND2X2 AND2X2_5506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9332_));
AND2X2 AND2X2_5507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9335_));
AND2X2 AND2X2_5508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9336_));
AND2X2 AND2X2_5509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9338_));
AND2X2 AND2X2_551 ( .A(_abc_44694_new_n1522__bF_buf1), .B(epc_q_8_), .Y(_abc_44694_new_n1641_));
AND2X2 AND2X2_5510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9339_));
AND2X2 AND2X2_5511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9344_));
AND2X2 AND2X2_5512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9345_));
AND2X2 AND2X2_5513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9347_));
AND2X2 AND2X2_5514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9348_));
AND2X2 AND2X2_5515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9351_));
AND2X2 AND2X2_5516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9352_));
AND2X2 AND2X2_5517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9354_));
AND2X2 AND2X2_5518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9355_));
AND2X2 AND2X2_5519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9359_));
AND2X2 AND2X2_552 ( .A(_abc_44694_new_n1348__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_8_), .Y(_abc_44694_new_n1642_));
AND2X2 AND2X2_5520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9360_));
AND2X2 AND2X2_5521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9362_));
AND2X2 AND2X2_5522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9363_));
AND2X2 AND2X2_5523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9366_));
AND2X2 AND2X2_5524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9367_));
AND2X2 AND2X2_5525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9369_));
AND2X2 AND2X2_5526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9370_));
AND2X2 AND2X2_5527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9376_));
AND2X2 AND2X2_5528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9377_));
AND2X2 AND2X2_5529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9379_));
AND2X2 AND2X2_553 ( .A(_abc_44694_new_n1207__bF_buf5), .B(_abc_44694_new_n1644_), .Y(_abc_44694_new_n1645_));
AND2X2 AND2X2_5530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9380_));
AND2X2 AND2X2_5531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9383_));
AND2X2 AND2X2_5532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9384_));
AND2X2 AND2X2_5533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9386_));
AND2X2 AND2X2_5534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9387_));
AND2X2 AND2X2_5535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9391_));
AND2X2 AND2X2_5536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9392_));
AND2X2 AND2X2_5537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9393_));
AND2X2 AND2X2_5538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9396_));
AND2X2 AND2X2_5539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9397_));
AND2X2 AND2X2_554 ( .A(_abc_44694_new_n1640_), .B(_abc_44694_new_n1645_), .Y(_abc_44694_new_n1646_));
AND2X2 AND2X2_5540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9399_));
AND2X2 AND2X2_5541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9400_));
AND2X2 AND2X2_5542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9405_));
AND2X2 AND2X2_5543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9406_));
AND2X2 AND2X2_5544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9408_));
AND2X2 AND2X2_5545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9409_));
AND2X2 AND2X2_5546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9412_));
AND2X2 AND2X2_5547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9413_));
AND2X2 AND2X2_5548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9415_));
AND2X2 AND2X2_5549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9416_));
AND2X2 AND2X2_555 ( .A(_abc_44694_new_n1648_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n1649_));
AND2X2 AND2X2_5550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9420_));
AND2X2 AND2X2_5551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9421_));
AND2X2 AND2X2_5552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9423_));
AND2X2 AND2X2_5553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9424_));
AND2X2 AND2X2_5554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9427_));
AND2X2 AND2X2_5555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9428_));
AND2X2 AND2X2_5556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9430_));
AND2X2 AND2X2_5557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9431_));
AND2X2 AND2X2_5558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9437_));
AND2X2 AND2X2_5559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9438_));
AND2X2 AND2X2_556 ( .A(_abc_44694_new_n1647_), .B(_abc_44694_new_n1649_), .Y(_0epc_q_31_0__8_));
AND2X2 AND2X2_5560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9440_));
AND2X2 AND2X2_5561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9441_));
AND2X2 AND2X2_5562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9444_));
AND2X2 AND2X2_5563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9445_));
AND2X2 AND2X2_5564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9447_));
AND2X2 AND2X2_5565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9448_));
AND2X2 AND2X2_5566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9452_));
AND2X2 AND2X2_5567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9453_));
AND2X2 AND2X2_5568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9454_));
AND2X2 AND2X2_5569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9457_));
AND2X2 AND2X2_557 ( .A(_abc_44694_new_n1615_), .B(pc_q_9_), .Y(_abc_44694_new_n1652_));
AND2X2 AND2X2_5570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9458_));
AND2X2 AND2X2_5571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9460_));
AND2X2 AND2X2_5572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9461_));
AND2X2 AND2X2_5573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9466_));
AND2X2 AND2X2_5574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9467_));
AND2X2 AND2X2_5575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9469_));
AND2X2 AND2X2_5576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9470_));
AND2X2 AND2X2_5577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9473_));
AND2X2 AND2X2_5578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9474_));
AND2X2 AND2X2_5579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9476_));
AND2X2 AND2X2_558 ( .A(_abc_44694_new_n1653_), .B(_abc_44694_new_n1651_), .Y(_abc_44694_new_n1654_));
AND2X2 AND2X2_5580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9477_));
AND2X2 AND2X2_5581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9481_));
AND2X2 AND2X2_5582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9482_));
AND2X2 AND2X2_5583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9484_));
AND2X2 AND2X2_5584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9485_));
AND2X2 AND2X2_5585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9488_));
AND2X2 AND2X2_5586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9489_));
AND2X2 AND2X2_5587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9491_));
AND2X2 AND2X2_5588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9492_));
AND2X2 AND2X2_5589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9498_));
AND2X2 AND2X2_559 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1655_), .Y(_abc_44694_new_n1656_));
AND2X2 AND2X2_5590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9499_));
AND2X2 AND2X2_5591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9501_));
AND2X2 AND2X2_5592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9502_));
AND2X2 AND2X2_5593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9505_));
AND2X2 AND2X2_5594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9506_));
AND2X2 AND2X2_5595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9508_));
AND2X2 AND2X2_5596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9509_));
AND2X2 AND2X2_5597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9513_));
AND2X2 AND2X2_5598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9514_));
AND2X2 AND2X2_5599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9515_));
AND2X2 AND2X2_56 ( .A(_abc_44694_new_n703_), .B(_abc_44694_new_n712_), .Y(_abc_44694_new_n713_));
AND2X2 AND2X2_560 ( .A(_abc_44694_new_n1019__bF_buf1), .B(epc_q_9_), .Y(_abc_44694_new_n1658_));
AND2X2 AND2X2_5600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9518_));
AND2X2 AND2X2_5601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9519_));
AND2X2 AND2X2_5602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9521_));
AND2X2 AND2X2_5603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9522_));
AND2X2 AND2X2_5604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9527_));
AND2X2 AND2X2_5605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9528_));
AND2X2 AND2X2_5606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9530_));
AND2X2 AND2X2_5607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9531_));
AND2X2 AND2X2_5608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9534_));
AND2X2 AND2X2_5609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9535_));
AND2X2 AND2X2_561 ( .A(_abc_44694_new_n1659_), .B(_abc_44694_new_n1021_), .Y(_abc_44694_new_n1660_));
AND2X2 AND2X2_5610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9537_));
AND2X2 AND2X2_5611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9538_));
AND2X2 AND2X2_5612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9542_));
AND2X2 AND2X2_5613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9543_));
AND2X2 AND2X2_5614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9545_));
AND2X2 AND2X2_5615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9546_));
AND2X2 AND2X2_5616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9549_));
AND2X2 AND2X2_5617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9550_));
AND2X2 AND2X2_5618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9552_));
AND2X2 AND2X2_5619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9553_));
AND2X2 AND2X2_562 ( .A(alu_op_r_5_), .B(pc_q_9_), .Y(_abc_44694_new_n1662_));
AND2X2 AND2X2_5620 ( .A(alu_b_i_20_), .B(alu_a_i_20_), .Y(alu__abc_42281_new_n110_));
AND2X2 AND2X2_5621 ( .A(alu__abc_42281_new_n112_), .B(alu__abc_42281_new_n113_), .Y(alu__abc_42281_new_n114_));
AND2X2 AND2X2_5622 ( .A(alu__abc_42281_new_n115_), .B(alu__abc_42281_new_n111_), .Y(alu__abc_42281_new_n116_));
AND2X2 AND2X2_5623 ( .A(alu_b_i_21_), .B(alu_a_i_21_), .Y(alu__abc_42281_new_n118_));
AND2X2 AND2X2_5624 ( .A(alu__abc_42281_new_n120_), .B(alu__abc_42281_new_n121_), .Y(alu__abc_42281_new_n122_));
AND2X2 AND2X2_5625 ( .A(alu__abc_42281_new_n123_), .B(alu__abc_42281_new_n119_), .Y(alu__abc_42281_new_n124_));
AND2X2 AND2X2_5626 ( .A(alu__abc_42281_new_n117_), .B(alu__abc_42281_new_n125_), .Y(alu__abc_42281_new_n126_));
AND2X2 AND2X2_5627 ( .A(alu_b_i_22_), .B(alu_a_i_22_), .Y(alu__abc_42281_new_n127_));
AND2X2 AND2X2_5628 ( .A(alu__abc_42281_new_n129_), .B(alu__abc_42281_new_n130_), .Y(alu__abc_42281_new_n131_));
AND2X2 AND2X2_5629 ( .A(alu__abc_42281_new_n132_), .B(alu__abc_42281_new_n128_), .Y(alu__abc_42281_new_n133_));
AND2X2 AND2X2_563 ( .A(_abc_44694_new_n1663_), .B(_abc_44694_new_n1661_), .Y(_abc_44694_new_n1664_));
AND2X2 AND2X2_5630 ( .A(alu_b_i_23_), .B(alu_a_i_23_), .Y(alu__abc_42281_new_n135_));
AND2X2 AND2X2_5631 ( .A(alu__abc_42281_new_n137_), .B(alu__abc_42281_new_n138_), .Y(alu__abc_42281_new_n139_));
AND2X2 AND2X2_5632 ( .A(alu__abc_42281_new_n140_), .B(alu__abc_42281_new_n136_), .Y(alu__abc_42281_new_n141_));
AND2X2 AND2X2_5633 ( .A(alu__abc_42281_new_n134_), .B(alu__abc_42281_new_n142_), .Y(alu__abc_42281_new_n143_));
AND2X2 AND2X2_5634 ( .A(alu__abc_42281_new_n126_), .B(alu__abc_42281_new_n143_), .Y(alu__abc_42281_new_n144_));
AND2X2 AND2X2_5635 ( .A(alu_b_i_18_), .B(alu_a_i_18_), .Y(alu__abc_42281_new_n145_));
AND2X2 AND2X2_5636 ( .A(alu__abc_42281_new_n147_), .B(alu__abc_42281_new_n148_), .Y(alu__abc_42281_new_n149_));
AND2X2 AND2X2_5637 ( .A(alu__abc_42281_new_n150_), .B(alu__abc_42281_new_n146_), .Y(alu__abc_42281_new_n151_));
AND2X2 AND2X2_5638 ( .A(alu_b_i_19_), .B(alu_a_i_19_), .Y(alu__abc_42281_new_n153_));
AND2X2 AND2X2_5639 ( .A(alu__abc_42281_new_n155_), .B(alu__abc_42281_new_n156_), .Y(alu__abc_42281_new_n157_));
AND2X2 AND2X2_564 ( .A(_abc_44694_new_n1664_), .B(_abc_44694_new_n1626_), .Y(_abc_44694_new_n1667_));
AND2X2 AND2X2_5640 ( .A(alu__abc_42281_new_n158_), .B(alu__abc_42281_new_n154_), .Y(alu__abc_42281_new_n159_));
AND2X2 AND2X2_5641 ( .A(alu__abc_42281_new_n152_), .B(alu__abc_42281_new_n160_), .Y(alu__abc_42281_new_n161_));
AND2X2 AND2X2_5642 ( .A(alu_b_i_16_), .B(alu_a_i_16_), .Y(alu__abc_42281_new_n162_));
AND2X2 AND2X2_5643 ( .A(alu__abc_42281_new_n164_), .B(alu__abc_42281_new_n165_), .Y(alu__abc_42281_new_n166_));
AND2X2 AND2X2_5644 ( .A(alu__abc_42281_new_n167_), .B(alu__abc_42281_new_n163_), .Y(alu__abc_42281_new_n168_));
AND2X2 AND2X2_5645 ( .A(alu_b_i_17_), .B(alu_a_i_17_), .Y(alu__abc_42281_new_n170_));
AND2X2 AND2X2_5646 ( .A(alu__abc_42281_new_n172_), .B(alu__abc_42281_new_n173_), .Y(alu__abc_42281_new_n174_));
AND2X2 AND2X2_5647 ( .A(alu__abc_42281_new_n175_), .B(alu__abc_42281_new_n171_), .Y(alu__abc_42281_new_n176_));
AND2X2 AND2X2_5648 ( .A(alu__abc_42281_new_n169_), .B(alu__abc_42281_new_n177_), .Y(alu__abc_42281_new_n178_));
AND2X2 AND2X2_5649 ( .A(alu__abc_42281_new_n161_), .B(alu__abc_42281_new_n178_), .Y(alu__abc_42281_new_n179_));
AND2X2 AND2X2_565 ( .A(_abc_44694_new_n1628_), .B(_abc_44694_new_n1664_), .Y(_abc_44694_new_n1669_));
AND2X2 AND2X2_5650 ( .A(alu__abc_42281_new_n144_), .B(alu__abc_42281_new_n179_), .Y(alu__abc_42281_new_n180_));
AND2X2 AND2X2_5651 ( .A(alu_b_i_25_), .B(alu_a_i_25_), .Y(alu__abc_42281_new_n181_));
AND2X2 AND2X2_5652 ( .A(alu__abc_42281_new_n183_), .B(alu__abc_42281_new_n184_), .Y(alu__abc_42281_new_n185_));
AND2X2 AND2X2_5653 ( .A(alu__abc_42281_new_n186_), .B(alu__abc_42281_new_n182_), .Y(alu__abc_42281_new_n187_));
AND2X2 AND2X2_5654 ( .A(alu_b_i_24_), .B(alu_a_i_24_), .Y(alu__abc_42281_new_n189_));
AND2X2 AND2X2_5655 ( .A(alu__abc_42281_new_n191_), .B(alu__abc_42281_new_n192_), .Y(alu__abc_42281_new_n193_));
AND2X2 AND2X2_5656 ( .A(alu__abc_42281_new_n194_), .B(alu__abc_42281_new_n190_), .Y(alu__abc_42281_new_n195_));
AND2X2 AND2X2_5657 ( .A(alu__abc_42281_new_n188_), .B(alu__abc_42281_new_n196_), .Y(alu__abc_42281_new_n197_));
AND2X2 AND2X2_5658 ( .A(alu_b_i_26_), .B(alu_a_i_26_), .Y(alu__abc_42281_new_n198_));
AND2X2 AND2X2_5659 ( .A(alu__abc_42281_new_n200_), .B(alu__abc_42281_new_n201_), .Y(alu__abc_42281_new_n202_));
AND2X2 AND2X2_566 ( .A(_abc_44694_new_n1624_), .B(_abc_44694_new_n1669_), .Y(_abc_44694_new_n1670_));
AND2X2 AND2X2_5660 ( .A(alu__abc_42281_new_n203_), .B(alu__abc_42281_new_n199_), .Y(alu__abc_42281_new_n204_));
AND2X2 AND2X2_5661 ( .A(alu_b_i_27_), .B(alu_a_i_27_), .Y(alu__abc_42281_new_n206_));
AND2X2 AND2X2_5662 ( .A(alu__abc_42281_new_n208_), .B(alu__abc_42281_new_n209_), .Y(alu__abc_42281_new_n210_));
AND2X2 AND2X2_5663 ( .A(alu__abc_42281_new_n211_), .B(alu__abc_42281_new_n207_), .Y(alu__abc_42281_new_n212_));
AND2X2 AND2X2_5664 ( .A(alu__abc_42281_new_n205_), .B(alu__abc_42281_new_n213_), .Y(alu__abc_42281_new_n214_));
AND2X2 AND2X2_5665 ( .A(alu__abc_42281_new_n197_), .B(alu__abc_42281_new_n214_), .Y(alu__abc_42281_new_n215_));
AND2X2 AND2X2_5666 ( .A(alu_b_i_28_), .B(alu_a_i_28_), .Y(alu__abc_42281_new_n216_));
AND2X2 AND2X2_5667 ( .A(alu__abc_42281_new_n218_), .B(alu__abc_42281_new_n219_), .Y(alu__abc_42281_new_n220_));
AND2X2 AND2X2_5668 ( .A(alu__abc_42281_new_n221_), .B(alu__abc_42281_new_n217_), .Y(alu__abc_42281_new_n222_));
AND2X2 AND2X2_5669 ( .A(alu_b_i_29_), .B(alu_a_i_29_), .Y(alu__abc_42281_new_n224_));
AND2X2 AND2X2_567 ( .A(_abc_44694_new_n1671_), .B(_abc_44694_new_n1668_), .Y(_abc_44694_new_n1672_));
AND2X2 AND2X2_5670 ( .A(alu__abc_42281_new_n226_), .B(alu__abc_42281_new_n227_), .Y(alu__abc_42281_new_n228_));
AND2X2 AND2X2_5671 ( .A(alu__abc_42281_new_n229_), .B(alu__abc_42281_new_n225_), .Y(alu__abc_42281_new_n230_));
AND2X2 AND2X2_5672 ( .A(alu__abc_42281_new_n223_), .B(alu__abc_42281_new_n231_), .Y(alu__abc_42281_new_n232_));
AND2X2 AND2X2_5673 ( .A(alu_b_i_30_), .B(alu_a_i_30_), .Y(alu__abc_42281_new_n233_));
AND2X2 AND2X2_5674 ( .A(alu__abc_42281_new_n235_), .B(alu__abc_42281_new_n236_), .Y(alu__abc_42281_new_n237_));
AND2X2 AND2X2_5675 ( .A(alu__abc_42281_new_n238_), .B(alu__abc_42281_new_n234_), .Y(alu__abc_42281_new_n239_));
AND2X2 AND2X2_5676 ( .A(alu_b_i_31_), .B(alu_a_i_31_), .Y(alu__abc_42281_new_n241_));
AND2X2 AND2X2_5677 ( .A(alu__abc_42281_new_n242_), .B(alu__abc_42281_new_n243_), .Y(alu__abc_42281_new_n244_));
AND2X2 AND2X2_5678 ( .A(alu__abc_42281_new_n240_), .B(alu__abc_42281_new_n245_), .Y(alu__abc_42281_new_n246_));
AND2X2 AND2X2_5679 ( .A(alu__abc_42281_new_n232_), .B(alu__abc_42281_new_n246_), .Y(alu__abc_42281_new_n247_));
AND2X2 AND2X2_568 ( .A(_abc_44694_new_n1672_), .B(_abc_44694_new_n1666_), .Y(_abc_44694_new_n1673_));
AND2X2 AND2X2_5680 ( .A(alu__abc_42281_new_n215_), .B(alu__abc_42281_new_n247_), .Y(alu__abc_42281_new_n248_));
AND2X2 AND2X2_5681 ( .A(alu__abc_42281_new_n180_), .B(alu__abc_42281_new_n248_), .Y(alu__abc_42281_new_n249_));
AND2X2 AND2X2_5682 ( .A(alu_b_i_6_), .B(alu_a_i_6_), .Y(alu__abc_42281_new_n250_));
AND2X2 AND2X2_5683 ( .A(alu__abc_42281_new_n252_), .B(alu__abc_42281_new_n253_), .Y(alu__abc_42281_new_n254_));
AND2X2 AND2X2_5684 ( .A(alu__abc_42281_new_n255_), .B(alu__abc_42281_new_n251_), .Y(alu__abc_42281_new_n256_));
AND2X2 AND2X2_5685 ( .A(alu_b_i_7_), .B(alu_a_i_7_), .Y(alu__abc_42281_new_n258_));
AND2X2 AND2X2_5686 ( .A(alu__abc_42281_new_n259_), .B(alu__abc_42281_new_n260_), .Y(alu__abc_42281_new_n261_));
AND2X2 AND2X2_5687 ( .A(alu__abc_42281_new_n257_), .B(alu__abc_42281_new_n262_), .Y(alu__abc_42281_new_n263_));
AND2X2 AND2X2_5688 ( .A(alu_b_i_5_), .B(alu_a_i_5_), .Y(alu__abc_42281_new_n264_));
AND2X2 AND2X2_5689 ( .A(alu__abc_42281_new_n265_), .B(alu__abc_42281_new_n266_), .Y(alu__abc_42281_new_n267_));
AND2X2 AND2X2_569 ( .A(_abc_44694_new_n1674_), .B(_abc_44694_new_n1660_), .Y(_abc_44694_new_n1675_));
AND2X2 AND2X2_5690 ( .A(alu_b_i_4_bF_buf5_), .B(alu_a_i_4_), .Y(alu__abc_42281_new_n269_));
AND2X2 AND2X2_5691 ( .A(alu__abc_42281_new_n271__bF_buf4), .B(alu__abc_42281_new_n272_), .Y(alu__abc_42281_new_n273_));
AND2X2 AND2X2_5692 ( .A(alu__abc_42281_new_n274_), .B(alu__abc_42281_new_n270_), .Y(alu__abc_42281_new_n275_));
AND2X2 AND2X2_5693 ( .A(alu__abc_42281_new_n276_), .B(alu__abc_42281_new_n268_), .Y(alu__abc_42281_new_n277_));
AND2X2 AND2X2_5694 ( .A(alu__abc_42281_new_n263_), .B(alu__abc_42281_new_n277_), .Y(alu__abc_42281_new_n278_));
AND2X2 AND2X2_5695 ( .A(alu_a_i_1_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n279_));
AND2X2 AND2X2_5696 ( .A(alu__abc_42281_new_n280_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n282_));
AND2X2 AND2X2_5697 ( .A(alu__abc_42281_new_n284_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n285_));
AND2X2 AND2X2_5698 ( .A(alu__abc_42281_new_n283_), .B(alu__abc_42281_new_n286_), .Y(alu__abc_42281_new_n287_));
AND2X2 AND2X2_5699 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_0_), .Y(alu__abc_42281_new_n289_));
AND2X2 AND2X2_57 ( .A(_abc_44694_new_n671_), .B(alu_p_o_2_), .Y(_abc_44694_new_n715_));
AND2X2 AND2X2_570 ( .A(_abc_44694_new_n1676_), .B(_abc_44694_new_n1340__bF_buf0), .Y(_abc_44694_new_n1677_));
AND2X2 AND2X2_5700 ( .A(alu__abc_42281_new_n287_), .B(alu__abc_42281_new_n290_), .Y(alu__abc_42281_new_n291_));
AND2X2 AND2X2_5701 ( .A(alu_a_i_2_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n292_));
AND2X2 AND2X2_5702 ( .A(alu__abc_42281_new_n293_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n295_));
AND2X2 AND2X2_5703 ( .A(alu_a_i_3_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n297_));
AND2X2 AND2X2_5704 ( .A(alu__abc_42281_new_n298_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n300_));
AND2X2 AND2X2_5705 ( .A(alu__abc_42281_new_n296_), .B(alu__abc_42281_new_n301_), .Y(alu__abc_42281_new_n302_));
AND2X2 AND2X2_5706 ( .A(alu__abc_42281_new_n291_), .B(alu__abc_42281_new_n302_), .Y(alu__abc_42281_new_n303_));
AND2X2 AND2X2_5707 ( .A(alu__abc_42281_new_n278_), .B(alu__abc_42281_new_n303_), .Y(alu__abc_42281_new_n304_));
AND2X2 AND2X2_5708 ( .A(alu_b_i_12_), .B(alu_a_i_12_), .Y(alu__abc_42281_new_n305_));
AND2X2 AND2X2_5709 ( .A(alu__abc_42281_new_n307_), .B(alu__abc_42281_new_n308_), .Y(alu__abc_42281_new_n309_));
AND2X2 AND2X2_571 ( .A(_abc_44694_new_n1337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n1678_));
AND2X2 AND2X2_5710 ( .A(alu__abc_42281_new_n310_), .B(alu__abc_42281_new_n306_), .Y(alu__abc_42281_new_n311_));
AND2X2 AND2X2_5711 ( .A(alu_b_i_13_), .B(alu_a_i_13_), .Y(alu__abc_42281_new_n313_));
AND2X2 AND2X2_5712 ( .A(alu__abc_42281_new_n315_), .B(alu__abc_42281_new_n316_), .Y(alu__abc_42281_new_n317_));
AND2X2 AND2X2_5713 ( .A(alu__abc_42281_new_n318_), .B(alu__abc_42281_new_n314_), .Y(alu__abc_42281_new_n319_));
AND2X2 AND2X2_5714 ( .A(alu__abc_42281_new_n312_), .B(alu__abc_42281_new_n320_), .Y(alu__abc_42281_new_n321_));
AND2X2 AND2X2_5715 ( .A(alu_b_i_14_), .B(alu_a_i_14_), .Y(alu__abc_42281_new_n322_));
AND2X2 AND2X2_5716 ( .A(alu__abc_42281_new_n324_), .B(alu__abc_42281_new_n325_), .Y(alu__abc_42281_new_n326_));
AND2X2 AND2X2_5717 ( .A(alu__abc_42281_new_n327_), .B(alu__abc_42281_new_n323_), .Y(alu__abc_42281_new_n328_));
AND2X2 AND2X2_5718 ( .A(alu_b_i_15_), .B(alu_a_i_15_), .Y(alu__abc_42281_new_n330_));
AND2X2 AND2X2_5719 ( .A(alu__abc_42281_new_n332_), .B(alu__abc_42281_new_n333_), .Y(alu__abc_42281_new_n334_));
AND2X2 AND2X2_572 ( .A(_abc_44694_new_n1680_), .B(_abc_44694_new_n1657_), .Y(_abc_44694_new_n1681_));
AND2X2 AND2X2_5720 ( .A(alu__abc_42281_new_n335_), .B(alu__abc_42281_new_n331_), .Y(alu__abc_42281_new_n336_));
AND2X2 AND2X2_5721 ( .A(alu__abc_42281_new_n329_), .B(alu__abc_42281_new_n337_), .Y(alu__abc_42281_new_n338_));
AND2X2 AND2X2_5722 ( .A(alu__abc_42281_new_n321_), .B(alu__abc_42281_new_n338_), .Y(alu__abc_42281_new_n339_));
AND2X2 AND2X2_5723 ( .A(alu_b_i_10_), .B(alu_a_i_10_), .Y(alu__abc_42281_new_n340_));
AND2X2 AND2X2_5724 ( .A(alu__abc_42281_new_n342_), .B(alu__abc_42281_new_n343_), .Y(alu__abc_42281_new_n344_));
AND2X2 AND2X2_5725 ( .A(alu__abc_42281_new_n345_), .B(alu__abc_42281_new_n341_), .Y(alu__abc_42281_new_n346_));
AND2X2 AND2X2_5726 ( .A(alu_b_i_11_), .B(alu_a_i_11_), .Y(alu__abc_42281_new_n348_));
AND2X2 AND2X2_5727 ( .A(alu__abc_42281_new_n350_), .B(alu__abc_42281_new_n351_), .Y(alu__abc_42281_new_n352_));
AND2X2 AND2X2_5728 ( .A(alu__abc_42281_new_n353_), .B(alu__abc_42281_new_n349_), .Y(alu__abc_42281_new_n354_));
AND2X2 AND2X2_5729 ( .A(alu__abc_42281_new_n347_), .B(alu__abc_42281_new_n355_), .Y(alu__abc_42281_new_n356_));
AND2X2 AND2X2_573 ( .A(_abc_44694_new_n1522__bF_buf0), .B(epc_q_9_), .Y(_abc_44694_new_n1683_));
AND2X2 AND2X2_5730 ( .A(alu_b_i_8_), .B(alu_a_i_8_), .Y(alu__abc_42281_new_n357_));
AND2X2 AND2X2_5731 ( .A(alu__abc_42281_new_n359_), .B(alu__abc_42281_new_n360_), .Y(alu__abc_42281_new_n361_));
AND2X2 AND2X2_5732 ( .A(alu__abc_42281_new_n362_), .B(alu__abc_42281_new_n358_), .Y(alu__abc_42281_new_n363_));
AND2X2 AND2X2_5733 ( .A(alu_b_i_9_), .B(alu_a_i_9_), .Y(alu__abc_42281_new_n365_));
AND2X2 AND2X2_5734 ( .A(alu__abc_42281_new_n367_), .B(alu__abc_42281_new_n368_), .Y(alu__abc_42281_new_n369_));
AND2X2 AND2X2_5735 ( .A(alu__abc_42281_new_n370_), .B(alu__abc_42281_new_n366_), .Y(alu__abc_42281_new_n371_));
AND2X2 AND2X2_5736 ( .A(alu__abc_42281_new_n364_), .B(alu__abc_42281_new_n372_), .Y(alu__abc_42281_new_n373_));
AND2X2 AND2X2_5737 ( .A(alu__abc_42281_new_n356_), .B(alu__abc_42281_new_n373_), .Y(alu__abc_42281_new_n374_));
AND2X2 AND2X2_5738 ( .A(alu__abc_42281_new_n339_), .B(alu__abc_42281_new_n374_), .Y(alu__abc_42281_new_n375_));
AND2X2 AND2X2_5739 ( .A(alu__abc_42281_new_n375_), .B(alu__abc_42281_new_n304_), .Y(alu__abc_42281_new_n376_));
AND2X2 AND2X2_574 ( .A(_abc_44694_new_n1348__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n1684_));
AND2X2 AND2X2_5740 ( .A(alu__abc_42281_new_n249_), .B(alu__abc_42281_new_n376_), .Y(alu_equal_o));
AND2X2 AND2X2_5741 ( .A(alu__abc_42281_new_n379_), .B(alu_op_i_2_), .Y(alu__abc_42281_new_n380_));
AND2X2 AND2X2_5742 ( .A(alu__abc_42281_new_n380_), .B(alu__abc_42281_new_n378_), .Y(alu_c_update_o));
AND2X2 AND2X2_5743 ( .A(alu__abc_42281_new_n382_), .B(alu_op_i_1_), .Y(alu__abc_42281_new_n383_));
AND2X2 AND2X2_5744 ( .A(alu__abc_42281_new_n384_), .B(alu_op_i_3_), .Y(alu__abc_42281_new_n385_));
AND2X2 AND2X2_5745 ( .A(alu__abc_42281_new_n383_), .B(alu__abc_42281_new_n385_), .Y(alu_flag_update_o));
AND2X2 AND2X2_5746 ( .A(alu__abc_42281_new_n242_), .B(alu_a_i_31_), .Y(alu__abc_42281_new_n387_));
AND2X2 AND2X2_5747 ( .A(alu__abc_42281_new_n259_), .B(alu_a_i_7_), .Y(alu__abc_42281_new_n388_));
AND2X2 AND2X2_5748 ( .A(alu__abc_42281_new_n260_), .B(alu_b_i_7_), .Y(alu__abc_42281_new_n389_));
AND2X2 AND2X2_5749 ( .A(alu__abc_42281_new_n252_), .B(alu_a_i_6_), .Y(alu__abc_42281_new_n391_));
AND2X2 AND2X2_575 ( .A(_abc_44694_new_n1207__bF_buf4), .B(_abc_44694_new_n1686_), .Y(_abc_44694_new_n1687_));
AND2X2 AND2X2_5750 ( .A(alu__abc_42281_new_n265_), .B(alu_a_i_5_), .Y(alu__abc_42281_new_n392_));
AND2X2 AND2X2_5751 ( .A(alu__abc_42281_new_n266_), .B(alu_b_i_5_), .Y(alu__abc_42281_new_n393_));
AND2X2 AND2X2_5752 ( .A(alu__abc_42281_new_n271__bF_buf3), .B(alu_a_i_4_), .Y(alu__abc_42281_new_n395_));
AND2X2 AND2X2_5753 ( .A(alu__abc_42281_new_n299__bF_buf5), .B(alu_a_i_3_), .Y(alu__abc_42281_new_n396_));
AND2X2 AND2X2_5754 ( .A(alu__abc_42281_new_n298_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n397_));
AND2X2 AND2X2_5755 ( .A(alu__abc_42281_new_n294__bF_buf5), .B(alu_a_i_2_), .Y(alu__abc_42281_new_n399_));
AND2X2 AND2X2_5756 ( .A(alu__abc_42281_new_n281__bF_buf5), .B(alu_a_i_1_), .Y(alu__abc_42281_new_n400_));
AND2X2 AND2X2_5757 ( .A(alu__abc_42281_new_n401_), .B(alu__abc_42281_new_n296_), .Y(alu__abc_42281_new_n402_));
AND2X2 AND2X2_5758 ( .A(alu__abc_42281_new_n403_), .B(alu__abc_42281_new_n398_), .Y(alu__abc_42281_new_n404_));
AND2X2 AND2X2_5759 ( .A(alu__abc_42281_new_n405_), .B(alu__abc_42281_new_n276_), .Y(alu__abc_42281_new_n406_));
AND2X2 AND2X2_576 ( .A(_abc_44694_new_n1682_), .B(_abc_44694_new_n1687_), .Y(_abc_44694_new_n1688_));
AND2X2 AND2X2_5760 ( .A(alu__abc_42281_new_n407_), .B(alu__abc_42281_new_n394_), .Y(alu__abc_42281_new_n408_));
AND2X2 AND2X2_5761 ( .A(alu__abc_42281_new_n409_), .B(alu__abc_42281_new_n257_), .Y(alu__abc_42281_new_n410_));
AND2X2 AND2X2_5762 ( .A(alu__abc_42281_new_n411_), .B(alu__abc_42281_new_n390_), .Y(alu__abc_42281_new_n412_));
AND2X2 AND2X2_5763 ( .A(alu__abc_42281_new_n413_), .B(alu__abc_42281_new_n375_), .Y(alu__abc_42281_new_n414_));
AND2X2 AND2X2_5764 ( .A(alu__abc_42281_new_n367_), .B(alu_a_i_9_), .Y(alu__abc_42281_new_n415_));
AND2X2 AND2X2_5765 ( .A(alu__abc_42281_new_n359_), .B(alu_a_i_8_), .Y(alu__abc_42281_new_n417_));
AND2X2 AND2X2_5766 ( .A(alu__abc_42281_new_n368_), .B(alu_b_i_9_), .Y(alu__abc_42281_new_n419_));
AND2X2 AND2X2_5767 ( .A(alu__abc_42281_new_n420_), .B(alu__abc_42281_new_n416_), .Y(alu__abc_42281_new_n421_));
AND2X2 AND2X2_5768 ( .A(alu__abc_42281_new_n422_), .B(alu__abc_42281_new_n356_), .Y(alu__abc_42281_new_n423_));
AND2X2 AND2X2_5769 ( .A(alu__abc_42281_new_n350_), .B(alu_a_i_11_), .Y(alu__abc_42281_new_n424_));
AND2X2 AND2X2_577 ( .A(_abc_44694_new_n1690_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n1691_));
AND2X2 AND2X2_5770 ( .A(alu__abc_42281_new_n342_), .B(alu_a_i_10_), .Y(alu__abc_42281_new_n425_));
AND2X2 AND2X2_5771 ( .A(alu__abc_42281_new_n355_), .B(alu__abc_42281_new_n425_), .Y(alu__abc_42281_new_n426_));
AND2X2 AND2X2_5772 ( .A(alu__abc_42281_new_n428_), .B(alu__abc_42281_new_n339_), .Y(alu__abc_42281_new_n429_));
AND2X2 AND2X2_5773 ( .A(alu__abc_42281_new_n315_), .B(alu_a_i_13_), .Y(alu__abc_42281_new_n430_));
AND2X2 AND2X2_5774 ( .A(alu__abc_42281_new_n307_), .B(alu_a_i_12_), .Y(alu__abc_42281_new_n432_));
AND2X2 AND2X2_5775 ( .A(alu__abc_42281_new_n316_), .B(alu_b_i_13_), .Y(alu__abc_42281_new_n434_));
AND2X2 AND2X2_5776 ( .A(alu__abc_42281_new_n435_), .B(alu__abc_42281_new_n431_), .Y(alu__abc_42281_new_n436_));
AND2X2 AND2X2_5777 ( .A(alu__abc_42281_new_n437_), .B(alu__abc_42281_new_n338_), .Y(alu__abc_42281_new_n438_));
AND2X2 AND2X2_5778 ( .A(alu__abc_42281_new_n332_), .B(alu_a_i_15_), .Y(alu__abc_42281_new_n439_));
AND2X2 AND2X2_5779 ( .A(alu__abc_42281_new_n324_), .B(alu_a_i_14_), .Y(alu__abc_42281_new_n440_));
AND2X2 AND2X2_578 ( .A(_abc_44694_new_n1689_), .B(_abc_44694_new_n1691_), .Y(_0epc_q_31_0__9_));
AND2X2 AND2X2_5780 ( .A(alu__abc_42281_new_n337_), .B(alu__abc_42281_new_n440_), .Y(alu__abc_42281_new_n441_));
AND2X2 AND2X2_5781 ( .A(alu__abc_42281_new_n445_), .B(alu__abc_42281_new_n180_), .Y(alu__abc_42281_new_n446_));
AND2X2 AND2X2_5782 ( .A(alu__abc_42281_new_n172_), .B(alu_a_i_17_), .Y(alu__abc_42281_new_n447_));
AND2X2 AND2X2_5783 ( .A(alu__abc_42281_new_n164_), .B(alu_a_i_16_), .Y(alu__abc_42281_new_n449_));
AND2X2 AND2X2_5784 ( .A(alu__abc_42281_new_n173_), .B(alu_b_i_17_), .Y(alu__abc_42281_new_n451_));
AND2X2 AND2X2_5785 ( .A(alu__abc_42281_new_n452_), .B(alu__abc_42281_new_n448_), .Y(alu__abc_42281_new_n453_));
AND2X2 AND2X2_5786 ( .A(alu__abc_42281_new_n454_), .B(alu__abc_42281_new_n161_), .Y(alu__abc_42281_new_n455_));
AND2X2 AND2X2_5787 ( .A(alu__abc_42281_new_n155_), .B(alu_a_i_19_), .Y(alu__abc_42281_new_n456_));
AND2X2 AND2X2_5788 ( .A(alu__abc_42281_new_n147_), .B(alu_a_i_18_), .Y(alu__abc_42281_new_n457_));
AND2X2 AND2X2_5789 ( .A(alu__abc_42281_new_n160_), .B(alu__abc_42281_new_n457_), .Y(alu__abc_42281_new_n458_));
AND2X2 AND2X2_579 ( .A(_abc_44694_new_n1652_), .B(pc_q_10_), .Y(_abc_44694_new_n1694_));
AND2X2 AND2X2_5790 ( .A(alu__abc_42281_new_n460_), .B(alu__abc_42281_new_n144_), .Y(alu__abc_42281_new_n461_));
AND2X2 AND2X2_5791 ( .A(alu__abc_42281_new_n120_), .B(alu_a_i_21_), .Y(alu__abc_42281_new_n462_));
AND2X2 AND2X2_5792 ( .A(alu__abc_42281_new_n112_), .B(alu_a_i_20_), .Y(alu__abc_42281_new_n464_));
AND2X2 AND2X2_5793 ( .A(alu__abc_42281_new_n121_), .B(alu_b_i_21_), .Y(alu__abc_42281_new_n466_));
AND2X2 AND2X2_5794 ( .A(alu__abc_42281_new_n467_), .B(alu__abc_42281_new_n463_), .Y(alu__abc_42281_new_n468_));
AND2X2 AND2X2_5795 ( .A(alu__abc_42281_new_n469_), .B(alu__abc_42281_new_n143_), .Y(alu__abc_42281_new_n470_));
AND2X2 AND2X2_5796 ( .A(alu__abc_42281_new_n137_), .B(alu_a_i_23_), .Y(alu__abc_42281_new_n471_));
AND2X2 AND2X2_5797 ( .A(alu__abc_42281_new_n129_), .B(alu_a_i_22_), .Y(alu__abc_42281_new_n472_));
AND2X2 AND2X2_5798 ( .A(alu__abc_42281_new_n142_), .B(alu__abc_42281_new_n472_), .Y(alu__abc_42281_new_n473_));
AND2X2 AND2X2_5799 ( .A(alu__abc_42281_new_n477_), .B(alu__abc_42281_new_n215_), .Y(alu__abc_42281_new_n478_));
AND2X2 AND2X2_58 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[2] ), .Y(_abc_44694_new_n716_));
AND2X2 AND2X2_580 ( .A(_abc_44694_new_n1695_), .B(_abc_44694_new_n1693_), .Y(_abc_44694_new_n1696_));
AND2X2 AND2X2_5800 ( .A(alu__abc_42281_new_n208_), .B(alu_a_i_27_), .Y(alu__abc_42281_new_n479_));
AND2X2 AND2X2_5801 ( .A(alu__abc_42281_new_n200_), .B(alu_a_i_26_), .Y(alu__abc_42281_new_n480_));
AND2X2 AND2X2_5802 ( .A(alu__abc_42281_new_n213_), .B(alu__abc_42281_new_n480_), .Y(alu__abc_42281_new_n481_));
AND2X2 AND2X2_5803 ( .A(alu__abc_42281_new_n184_), .B(alu_b_i_25_), .Y(alu__abc_42281_new_n485_));
AND2X2 AND2X2_5804 ( .A(alu__abc_42281_new_n183_), .B(alu_a_i_25_), .Y(alu__abc_42281_new_n486_));
AND2X2 AND2X2_5805 ( .A(alu__abc_42281_new_n191_), .B(alu_a_i_24_), .Y(alu__abc_42281_new_n488_));
AND2X2 AND2X2_5806 ( .A(alu__abc_42281_new_n487_), .B(alu__abc_42281_new_n489_), .Y(alu__abc_42281_new_n490_));
AND2X2 AND2X2_5807 ( .A(alu__abc_42281_new_n492_), .B(alu__abc_42281_new_n483_), .Y(alu__abc_42281_new_n493_));
AND2X2 AND2X2_5808 ( .A(alu__abc_42281_new_n495_), .B(alu__abc_42281_new_n232_), .Y(alu__abc_42281_new_n496_));
AND2X2 AND2X2_5809 ( .A(alu__abc_42281_new_n227_), .B(alu_b_i_29_), .Y(alu__abc_42281_new_n497_));
AND2X2 AND2X2_581 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1697_), .Y(_abc_44694_new_n1698_));
AND2X2 AND2X2_5810 ( .A(alu__abc_42281_new_n226_), .B(alu_a_i_29_), .Y(alu__abc_42281_new_n498_));
AND2X2 AND2X2_5811 ( .A(alu__abc_42281_new_n218_), .B(alu_a_i_28_), .Y(alu__abc_42281_new_n500_));
AND2X2 AND2X2_5812 ( .A(alu__abc_42281_new_n499_), .B(alu__abc_42281_new_n501_), .Y(alu__abc_42281_new_n502_));
AND2X2 AND2X2_5813 ( .A(alu__abc_42281_new_n505_), .B(alu__abc_42281_new_n240_), .Y(alu__abc_42281_new_n506_));
AND2X2 AND2X2_5814 ( .A(alu__abc_42281_new_n235_), .B(alu_a_i_30_), .Y(alu__abc_42281_new_n507_));
AND2X2 AND2X2_5815 ( .A(alu__abc_42281_new_n509_), .B(alu__abc_42281_new_n245_), .Y(alu__abc_42281_new_n510_));
AND2X2 AND2X2_5816 ( .A(alu__abc_42281_new_n512_), .B(alu__abc_42281_new_n239_), .Y(alu__abc_42281_new_n513_));
AND2X2 AND2X2_5817 ( .A(alu__abc_42281_new_n222_), .B(alu__abc_42281_new_n230_), .Y(alu__abc_42281_new_n514_));
AND2X2 AND2X2_5818 ( .A(alu__abc_42281_new_n513_), .B(alu__abc_42281_new_n514_), .Y(alu__abc_42281_new_n515_));
AND2X2 AND2X2_5819 ( .A(alu__abc_42281_new_n199_), .B(alu__abc_42281_new_n207_), .Y(alu__abc_42281_new_n516_));
AND2X2 AND2X2_582 ( .A(_abc_44694_new_n1671_), .B(_abc_44694_new_n1700_), .Y(_abc_44694_new_n1701_));
AND2X2 AND2X2_5820 ( .A(alu__abc_42281_new_n204_), .B(alu__abc_42281_new_n212_), .Y(alu__abc_42281_new_n519_));
AND2X2 AND2X2_5821 ( .A(alu__abc_42281_new_n182_), .B(alu__abc_42281_new_n190_), .Y(alu__abc_42281_new_n520_));
AND2X2 AND2X2_5822 ( .A(alu__abc_42281_new_n522_), .B(alu__abc_42281_new_n519_), .Y(alu__abc_42281_new_n523_));
AND2X2 AND2X2_5823 ( .A(alu__abc_42281_new_n524_), .B(alu__abc_42281_new_n515_), .Y(alu__abc_42281_new_n525_));
AND2X2 AND2X2_5824 ( .A(alu__abc_42281_new_n217_), .B(alu__abc_42281_new_n225_), .Y(alu__abc_42281_new_n526_));
AND2X2 AND2X2_5825 ( .A(alu__abc_42281_new_n528_), .B(alu__abc_42281_new_n513_), .Y(alu__abc_42281_new_n529_));
AND2X2 AND2X2_5826 ( .A(alu__abc_42281_new_n530_), .B(alu__abc_42281_new_n233_), .Y(alu__abc_42281_new_n531_));
AND2X2 AND2X2_5827 ( .A(alu__abc_42281_new_n133_), .B(alu__abc_42281_new_n141_), .Y(alu__abc_42281_new_n535_));
AND2X2 AND2X2_5828 ( .A(alu__abc_42281_new_n116_), .B(alu__abc_42281_new_n124_), .Y(alu__abc_42281_new_n536_));
AND2X2 AND2X2_5829 ( .A(alu__abc_42281_new_n535_), .B(alu__abc_42281_new_n536_), .Y(alu__abc_42281_new_n537_));
AND2X2 AND2X2_583 ( .A(alu_op_r_6_), .B(pc_q_10_), .Y(_abc_44694_new_n1704_));
AND2X2 AND2X2_5830 ( .A(alu__abc_42281_new_n151_), .B(alu__abc_42281_new_n159_), .Y(alu__abc_42281_new_n538_));
AND2X2 AND2X2_5831 ( .A(alu__abc_42281_new_n163_), .B(alu__abc_42281_new_n171_), .Y(alu__abc_42281_new_n539_));
AND2X2 AND2X2_5832 ( .A(alu__abc_42281_new_n541_), .B(alu__abc_42281_new_n538_), .Y(alu__abc_42281_new_n542_));
AND2X2 AND2X2_5833 ( .A(alu__abc_42281_new_n158_), .B(alu__abc_42281_new_n145_), .Y(alu__abc_42281_new_n543_));
AND2X2 AND2X2_5834 ( .A(alu__abc_42281_new_n545_), .B(alu__abc_42281_new_n537_), .Y(alu__abc_42281_new_n546_));
AND2X2 AND2X2_5835 ( .A(alu__abc_42281_new_n111_), .B(alu__abc_42281_new_n119_), .Y(alu__abc_42281_new_n547_));
AND2X2 AND2X2_5836 ( .A(alu__abc_42281_new_n549_), .B(alu__abc_42281_new_n535_), .Y(alu__abc_42281_new_n550_));
AND2X2 AND2X2_5837 ( .A(alu__abc_42281_new_n140_), .B(alu__abc_42281_new_n127_), .Y(alu__abc_42281_new_n551_));
AND2X2 AND2X2_5838 ( .A(alu__abc_42281_new_n336_), .B(alu__abc_42281_new_n322_), .Y(alu__abc_42281_new_n555_));
AND2X2 AND2X2_5839 ( .A(alu__abc_42281_new_n318_), .B(alu__abc_42281_new_n305_), .Y(alu__abc_42281_new_n557_));
AND2X2 AND2X2_584 ( .A(_abc_44694_new_n1705_), .B(_abc_44694_new_n1703_), .Y(_abc_44694_new_n1706_));
AND2X2 AND2X2_5840 ( .A(alu__abc_42281_new_n328_), .B(alu__abc_42281_new_n336_), .Y(alu__abc_42281_new_n559_));
AND2X2 AND2X2_5841 ( .A(alu__abc_42281_new_n558_), .B(alu__abc_42281_new_n559_), .Y(alu__abc_42281_new_n560_));
AND2X2 AND2X2_5842 ( .A(alu__abc_42281_new_n346_), .B(alu__abc_42281_new_n354_), .Y(alu__abc_42281_new_n562_));
AND2X2 AND2X2_5843 ( .A(alu__abc_42281_new_n358_), .B(alu__abc_42281_new_n366_), .Y(alu__abc_42281_new_n563_));
AND2X2 AND2X2_5844 ( .A(alu__abc_42281_new_n565_), .B(alu__abc_42281_new_n562_), .Y(alu__abc_42281_new_n566_));
AND2X2 AND2X2_5845 ( .A(alu__abc_42281_new_n353_), .B(alu__abc_42281_new_n340_), .Y(alu__abc_42281_new_n567_));
AND2X2 AND2X2_5846 ( .A(alu__abc_42281_new_n311_), .B(alu__abc_42281_new_n319_), .Y(alu__abc_42281_new_n570_));
AND2X2 AND2X2_5847 ( .A(alu__abc_42281_new_n570_), .B(alu__abc_42281_new_n559_), .Y(alu__abc_42281_new_n571_));
AND2X2 AND2X2_5848 ( .A(alu__abc_42281_new_n569_), .B(alu__abc_42281_new_n571_), .Y(alu__abc_42281_new_n572_));
AND2X2 AND2X2_5849 ( .A(alu__abc_42281_new_n574_), .B(alu__abc_42281_new_n575_), .Y(alu__abc_42281_new_n576_));
AND2X2 AND2X2_585 ( .A(_abc_44694_new_n1702_), .B(_abc_44694_new_n1706_), .Y(_abc_44694_new_n1707_));
AND2X2 AND2X2_5850 ( .A(alu_b_i_0_bF_buf2_), .B(alu_a_i_0_), .Y(alu__abc_42281_new_n577_));
AND2X2 AND2X2_5851 ( .A(alu__abc_42281_new_n576_), .B(alu__abc_42281_new_n577_), .Y(alu__abc_42281_new_n578_));
AND2X2 AND2X2_5852 ( .A(alu__abc_42281_new_n579_), .B(alu__abc_42281_new_n581_), .Y(alu__abc_42281_new_n582_));
AND2X2 AND2X2_5853 ( .A(alu__abc_42281_new_n583_), .B(alu__abc_42281_new_n292_), .Y(alu__abc_42281_new_n584_));
AND2X2 AND2X2_5854 ( .A(alu__abc_42281_new_n587_), .B(alu__abc_42281_new_n256_), .Y(alu__abc_42281_new_n588_));
AND2X2 AND2X2_5855 ( .A(alu__abc_42281_new_n589_), .B(alu__abc_42281_new_n275_), .Y(alu__abc_42281_new_n590_));
AND2X2 AND2X2_5856 ( .A(alu__abc_42281_new_n588_), .B(alu__abc_42281_new_n590_), .Y(alu__abc_42281_new_n591_));
AND2X2 AND2X2_5857 ( .A(alu__abc_42281_new_n586_), .B(alu__abc_42281_new_n591_), .Y(alu__abc_42281_new_n592_));
AND2X2 AND2X2_5858 ( .A(alu__abc_42281_new_n594_), .B(alu__abc_42281_new_n593_), .Y(alu__abc_42281_new_n595_));
AND2X2 AND2X2_5859 ( .A(alu__abc_42281_new_n588_), .B(alu__abc_42281_new_n595_), .Y(alu__abc_42281_new_n596_));
AND2X2 AND2X2_586 ( .A(_abc_44694_new_n1708_), .B(_abc_44694_new_n1709_), .Y(_abc_44694_new_n1710_));
AND2X2 AND2X2_5860 ( .A(alu__abc_42281_new_n597_), .B(alu__abc_42281_new_n250_), .Y(alu__abc_42281_new_n598_));
AND2X2 AND2X2_5861 ( .A(alu__abc_42281_new_n363_), .B(alu__abc_42281_new_n371_), .Y(alu__abc_42281_new_n602_));
AND2X2 AND2X2_5862 ( .A(alu__abc_42281_new_n562_), .B(alu__abc_42281_new_n602_), .Y(alu__abc_42281_new_n603_));
AND2X2 AND2X2_5863 ( .A(alu__abc_42281_new_n603_), .B(alu__abc_42281_new_n571_), .Y(alu__abc_42281_new_n604_));
AND2X2 AND2X2_5864 ( .A(alu__abc_42281_new_n601_), .B(alu__abc_42281_new_n604_), .Y(alu__abc_42281_new_n605_));
AND2X2 AND2X2_5865 ( .A(alu__abc_42281_new_n168_), .B(alu__abc_42281_new_n176_), .Y(alu__abc_42281_new_n607_));
AND2X2 AND2X2_5866 ( .A(alu__abc_42281_new_n606_), .B(alu__abc_42281_new_n607_), .Y(alu__abc_42281_new_n608_));
AND2X2 AND2X2_5867 ( .A(alu__abc_42281_new_n608_), .B(alu__abc_42281_new_n538_), .Y(alu__abc_42281_new_n609_));
AND2X2 AND2X2_5868 ( .A(alu__abc_42281_new_n609_), .B(alu__abc_42281_new_n537_), .Y(alu__abc_42281_new_n610_));
AND2X2 AND2X2_5869 ( .A(alu__abc_42281_new_n611_), .B(alu__abc_42281_new_n195_), .Y(alu__abc_42281_new_n612_));
AND2X2 AND2X2_587 ( .A(_abc_44694_new_n1340__bF_buf4), .B(_abc_44694_new_n1712_), .Y(_abc_44694_new_n1713_));
AND2X2 AND2X2_5870 ( .A(alu__abc_42281_new_n612_), .B(alu__abc_42281_new_n187_), .Y(alu__abc_42281_new_n613_));
AND2X2 AND2X2_5871 ( .A(alu__abc_42281_new_n515_), .B(alu__abc_42281_new_n519_), .Y(alu__abc_42281_new_n614_));
AND2X2 AND2X2_5872 ( .A(alu__abc_42281_new_n613_), .B(alu__abc_42281_new_n614_), .Y(alu__abc_42281_new_n615_));
AND2X2 AND2X2_5873 ( .A(alu__abc_42281_new_n617_), .B(alu__abc_42281_new_n519_), .Y(alu__abc_42281_new_n618_));
AND2X2 AND2X2_5874 ( .A(alu__abc_42281_new_n619_), .B(alu__abc_42281_new_n514_), .Y(alu__abc_42281_new_n620_));
AND2X2 AND2X2_5875 ( .A(alu__abc_42281_new_n621_), .B(alu__abc_42281_new_n239_), .Y(alu__abc_42281_new_n622_));
AND2X2 AND2X2_5876 ( .A(alu__abc_42281_new_n623_), .B(alu__abc_42281_new_n234_), .Y(alu__abc_42281_new_n624_));
AND2X2 AND2X2_5877 ( .A(alu__abc_42281_new_n626_), .B(alu__abc_42281_new_n627_), .Y(alu__abc_42281_new_n628_));
AND2X2 AND2X2_5878 ( .A(alu__abc_42281_new_n623_), .B(alu__abc_42281_new_n629_), .Y(alu__abc_42281_new_n630_));
AND2X2 AND2X2_5879 ( .A(alu__abc_42281_new_n619_), .B(alu__abc_42281_new_n222_), .Y(alu__abc_42281_new_n631_));
AND2X2 AND2X2_588 ( .A(_abc_44694_new_n1711_), .B(_abc_44694_new_n1713_), .Y(_abc_44694_new_n1714_));
AND2X2 AND2X2_5880 ( .A(alu__abc_42281_new_n632_), .B(alu__abc_42281_new_n217_), .Y(alu__abc_42281_new_n633_));
AND2X2 AND2X2_5881 ( .A(alu__abc_42281_new_n635_), .B(alu__abc_42281_new_n636_), .Y(alu__abc_42281_new_n637_));
AND2X2 AND2X2_5882 ( .A(alu__abc_42281_new_n632_), .B(alu__abc_42281_new_n638_), .Y(alu__abc_42281_new_n639_));
AND2X2 AND2X2_5883 ( .A(alu__abc_42281_new_n617_), .B(alu__abc_42281_new_n204_), .Y(alu__abc_42281_new_n640_));
AND2X2 AND2X2_5884 ( .A(alu__abc_42281_new_n641_), .B(alu__abc_42281_new_n199_), .Y(alu__abc_42281_new_n642_));
AND2X2 AND2X2_5885 ( .A(alu__abc_42281_new_n644_), .B(alu__abc_42281_new_n645_), .Y(alu__abc_42281_new_n646_));
AND2X2 AND2X2_5886 ( .A(alu__abc_42281_new_n646_), .B(alu__abc_42281_new_n639_), .Y(alu__abc_42281_new_n647_));
AND2X2 AND2X2_5887 ( .A(alu__abc_42281_new_n648_), .B(alu__abc_42281_new_n649_), .Y(alu__abc_42281_new_n650_));
AND2X2 AND2X2_5888 ( .A(alu__abc_42281_new_n651_), .B(alu__abc_42281_new_n116_), .Y(alu__abc_42281_new_n652_));
AND2X2 AND2X2_5889 ( .A(alu__abc_42281_new_n653_), .B(alu__abc_42281_new_n111_), .Y(alu__abc_42281_new_n654_));
AND2X2 AND2X2_589 ( .A(_abc_44694_new_n1337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n1715_));
AND2X2 AND2X2_5890 ( .A(alu__abc_42281_new_n656_), .B(alu__abc_42281_new_n657_), .Y(alu__abc_42281_new_n658_));
AND2X2 AND2X2_5891 ( .A(alu__abc_42281_new_n651_), .B(alu__abc_42281_new_n536_), .Y(alu__abc_42281_new_n659_));
AND2X2 AND2X2_5892 ( .A(alu__abc_42281_new_n660_), .B(alu__abc_42281_new_n133_), .Y(alu__abc_42281_new_n661_));
AND2X2 AND2X2_5893 ( .A(alu__abc_42281_new_n662_), .B(alu__abc_42281_new_n663_), .Y(alu__abc_42281_new_n664_));
AND2X2 AND2X2_5894 ( .A(alu__abc_42281_new_n658_), .B(alu__abc_42281_new_n664_), .Y(alu__abc_42281_new_n665_));
AND2X2 AND2X2_5895 ( .A(alu__abc_42281_new_n665_), .B(alu__abc_42281_new_n650_), .Y(alu__abc_42281_new_n666_));
AND2X2 AND2X2_5896 ( .A(alu__abc_42281_new_n648_), .B(alu__abc_42281_new_n190_), .Y(alu__abc_42281_new_n667_));
AND2X2 AND2X2_5897 ( .A(alu__abc_42281_new_n669_), .B(alu__abc_42281_new_n670_), .Y(alu__abc_42281_new_n671_));
AND2X2 AND2X2_5898 ( .A(alu__abc_42281_new_n653_), .B(alu__abc_42281_new_n672_), .Y(alu__abc_42281_new_n673_));
AND2X2 AND2X2_5899 ( .A(alu__abc_42281_new_n674_), .B(alu__abc_42281_new_n151_), .Y(alu__abc_42281_new_n675_));
AND2X2 AND2X2_59 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[18] ), .Y(_abc_44694_new_n717_));
AND2X2 AND2X2_590 ( .A(_abc_44694_new_n1716_), .B(_abc_44694_new_n1399__bF_buf0), .Y(_abc_44694_new_n1717_));
AND2X2 AND2X2_5900 ( .A(alu__abc_42281_new_n676_), .B(alu__abc_42281_new_n146_), .Y(alu__abc_42281_new_n677_));
AND2X2 AND2X2_5901 ( .A(alu__abc_42281_new_n679_), .B(alu__abc_42281_new_n680_), .Y(alu__abc_42281_new_n681_));
AND2X2 AND2X2_5902 ( .A(alu__abc_42281_new_n676_), .B(alu__abc_42281_new_n682_), .Y(alu__abc_42281_new_n683_));
AND2X2 AND2X2_5903 ( .A(alu__abc_42281_new_n606_), .B(alu__abc_42281_new_n168_), .Y(alu__abc_42281_new_n684_));
AND2X2 AND2X2_5904 ( .A(alu__abc_42281_new_n685_), .B(alu__abc_42281_new_n163_), .Y(alu__abc_42281_new_n686_));
AND2X2 AND2X2_5905 ( .A(alu__abc_42281_new_n686_), .B(alu__abc_42281_new_n177_), .Y(alu__abc_42281_new_n687_));
AND2X2 AND2X2_5906 ( .A(alu__abc_42281_new_n688_), .B(alu__abc_42281_new_n689_), .Y(alu__abc_42281_new_n690_));
AND2X2 AND2X2_5907 ( .A(alu__abc_42281_new_n685_), .B(alu__abc_42281_new_n691_), .Y(alu__abc_42281_new_n692_));
AND2X2 AND2X2_5908 ( .A(alu__abc_42281_new_n697_), .B(alu__abc_42281_new_n574_), .Y(alu__abc_42281_new_n698_));
AND2X2 AND2X2_5909 ( .A(alu__abc_42281_new_n699_), .B(alu__abc_42281_new_n700_), .Y(alu__abc_42281_new_n701_));
AND2X2 AND2X2_591 ( .A(_abc_44694_new_n1400__bF_buf1), .B(_abc_44694_new_n1696_), .Y(_abc_44694_new_n1718_));
AND2X2 AND2X2_5910 ( .A(alu__abc_42281_new_n703_), .B(alu__abc_42281_new_n704_), .Y(alu__abc_42281_new_n705_));
AND2X2 AND2X2_5911 ( .A(alu__abc_42281_new_n707_), .B(alu__abc_42281_new_n695_), .Y(alu__abc_42281_new_n708_));
AND2X2 AND2X2_5912 ( .A(alu__abc_42281_new_n709_), .B(alu__abc_42281_new_n693_), .Y(alu__abc_42281_new_n710_));
AND2X2 AND2X2_5913 ( .A(alu__abc_42281_new_n711_), .B(alu__abc_42281_new_n323_), .Y(alu__abc_42281_new_n712_));
AND2X2 AND2X2_5914 ( .A(alu__abc_42281_new_n601_), .B(alu__abc_42281_new_n603_), .Y(alu__abc_42281_new_n714_));
AND2X2 AND2X2_5915 ( .A(alu__abc_42281_new_n715_), .B(alu__abc_42281_new_n570_), .Y(alu__abc_42281_new_n716_));
AND2X2 AND2X2_5916 ( .A(alu__abc_42281_new_n717_), .B(alu__abc_42281_new_n328_), .Y(alu__abc_42281_new_n718_));
AND2X2 AND2X2_5917 ( .A(alu__abc_42281_new_n713_), .B(alu__abc_42281_new_n720_), .Y(alu__abc_42281_new_n721_));
AND2X2 AND2X2_5918 ( .A(alu__abc_42281_new_n601_), .B(alu__abc_42281_new_n363_), .Y(alu__abc_42281_new_n722_));
AND2X2 AND2X2_5919 ( .A(alu__abc_42281_new_n723_), .B(alu__abc_42281_new_n358_), .Y(alu__abc_42281_new_n724_));
AND2X2 AND2X2_592 ( .A(_abc_44694_new_n1522__bF_buf4), .B(epc_q_10_), .Y(_abc_44694_new_n1721_));
AND2X2 AND2X2_5920 ( .A(alu__abc_42281_new_n726_), .B(alu__abc_42281_new_n727_), .Y(alu__abc_42281_new_n728_));
AND2X2 AND2X2_5921 ( .A(alu__abc_42281_new_n705_), .B(alu__abc_42281_new_n364_), .Y(alu__abc_42281_new_n729_));
AND2X2 AND2X2_5922 ( .A(alu__abc_42281_new_n586_), .B(alu__abc_42281_new_n590_), .Y(alu__abc_42281_new_n732_));
AND2X2 AND2X2_5923 ( .A(alu__abc_42281_new_n733_), .B(alu__abc_42281_new_n256_), .Y(alu__abc_42281_new_n734_));
AND2X2 AND2X2_5924 ( .A(alu__abc_42281_new_n735_), .B(alu__abc_42281_new_n251_), .Y(alu__abc_42281_new_n736_));
AND2X2 AND2X2_5925 ( .A(alu__abc_42281_new_n738_), .B(alu__abc_42281_new_n739_), .Y(alu__abc_42281_new_n740_));
AND2X2 AND2X2_5926 ( .A(alu__abc_42281_new_n735_), .B(alu__abc_42281_new_n741_), .Y(alu__abc_42281_new_n742_));
AND2X2 AND2X2_5927 ( .A(alu__abc_42281_new_n586_), .B(alu__abc_42281_new_n275_), .Y(alu__abc_42281_new_n743_));
AND2X2 AND2X2_5928 ( .A(alu__abc_42281_new_n744_), .B(alu__abc_42281_new_n270_), .Y(alu__abc_42281_new_n745_));
AND2X2 AND2X2_5929 ( .A(alu__abc_42281_new_n747_), .B(alu__abc_42281_new_n748_), .Y(alu__abc_42281_new_n749_));
AND2X2 AND2X2_593 ( .A(_abc_44694_new_n1348__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n1722_));
AND2X2 AND2X2_5930 ( .A(alu__abc_42281_new_n579_), .B(alu__abc_42281_new_n751_), .Y(alu__abc_42281_new_n752_));
AND2X2 AND2X2_5931 ( .A(alu__abc_42281_new_n756_), .B(alu__abc_42281_new_n754_), .Y(alu__abc_42281_new_n757_));
AND2X2 AND2X2_5932 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu__abc_42281_new_n284_), .Y(alu__abc_42281_new_n758_));
AND2X2 AND2X2_5933 ( .A(alu__abc_42281_new_n759_), .B(alu__abc_42281_new_n696_), .Y(alu__abc_42281_new_n760_));
AND2X2 AND2X2_5934 ( .A(alu__abc_42281_new_n760_), .B(alu_c_i), .Y(alu__abc_42281_new_n761_));
AND2X2 AND2X2_5935 ( .A(alu__abc_42281_new_n761_), .B(alu__abc_42281_new_n576_), .Y(alu__abc_42281_new_n762_));
AND2X2 AND2X2_5936 ( .A(alu__abc_42281_new_n698_), .B(alu__abc_42281_new_n296_), .Y(alu__abc_42281_new_n763_));
AND2X2 AND2X2_5937 ( .A(alu__abc_42281_new_n765_), .B(alu__abc_42281_new_n762_), .Y(alu__abc_42281_new_n766_));
AND2X2 AND2X2_5938 ( .A(alu__abc_42281_new_n757_), .B(alu__abc_42281_new_n766_), .Y(alu__abc_42281_new_n767_));
AND2X2 AND2X2_5939 ( .A(alu__abc_42281_new_n744_), .B(alu__abc_42281_new_n768_), .Y(alu__abc_42281_new_n769_));
AND2X2 AND2X2_594 ( .A(_abc_44694_new_n1207__bF_buf3), .B(_abc_44694_new_n1724_), .Y(_abc_44694_new_n1725_));
AND2X2 AND2X2_5940 ( .A(alu__abc_42281_new_n767_), .B(alu__abc_42281_new_n769_), .Y(alu__abc_42281_new_n770_));
AND2X2 AND2X2_5941 ( .A(alu__abc_42281_new_n749_), .B(alu__abc_42281_new_n770_), .Y(alu__abc_42281_new_n771_));
AND2X2 AND2X2_5942 ( .A(alu__abc_42281_new_n771_), .B(alu__abc_42281_new_n742_), .Y(alu__abc_42281_new_n772_));
AND2X2 AND2X2_5943 ( .A(alu__abc_42281_new_n740_), .B(alu__abc_42281_new_n772_), .Y(alu__abc_42281_new_n773_));
AND2X2 AND2X2_5944 ( .A(alu__abc_42281_new_n773_), .B(alu__abc_42281_new_n731_), .Y(alu__abc_42281_new_n774_));
AND2X2 AND2X2_5945 ( .A(alu__abc_42281_new_n774_), .B(alu__abc_42281_new_n728_), .Y(alu__abc_42281_new_n775_));
AND2X2 AND2X2_5946 ( .A(alu__abc_42281_new_n715_), .B(alu__abc_42281_new_n311_), .Y(alu__abc_42281_new_n776_));
AND2X2 AND2X2_5947 ( .A(alu__abc_42281_new_n779_), .B(alu__abc_42281_new_n306_), .Y(alu__abc_42281_new_n780_));
AND2X2 AND2X2_5948 ( .A(alu__abc_42281_new_n781_), .B(alu__abc_42281_new_n778_), .Y(alu__abc_42281_new_n782_));
AND2X2 AND2X2_5949 ( .A(alu__abc_42281_new_n784_), .B(alu__abc_42281_new_n564_), .Y(alu__abc_42281_new_n785_));
AND2X2 AND2X2_595 ( .A(_abc_44694_new_n1720_), .B(_abc_44694_new_n1725_), .Y(_abc_44694_new_n1726_));
AND2X2 AND2X2_5950 ( .A(alu__abc_42281_new_n601_), .B(alu__abc_42281_new_n602_), .Y(alu__abc_42281_new_n787_));
AND2X2 AND2X2_5951 ( .A(alu__abc_42281_new_n786_), .B(alu__abc_42281_new_n789_), .Y(alu__abc_42281_new_n790_));
AND2X2 AND2X2_5952 ( .A(alu__abc_42281_new_n779_), .B(alu__abc_42281_new_n791_), .Y(alu__abc_42281_new_n792_));
AND2X2 AND2X2_5953 ( .A(alu__abc_42281_new_n790_), .B(alu__abc_42281_new_n792_), .Y(alu__abc_42281_new_n793_));
AND2X2 AND2X2_5954 ( .A(alu__abc_42281_new_n782_), .B(alu__abc_42281_new_n793_), .Y(alu__abc_42281_new_n794_));
AND2X2 AND2X2_5955 ( .A(alu__abc_42281_new_n788_), .B(alu__abc_42281_new_n346_), .Y(alu__abc_42281_new_n795_));
AND2X2 AND2X2_5956 ( .A(alu__abc_42281_new_n786_), .B(alu__abc_42281_new_n341_), .Y(alu__abc_42281_new_n798_));
AND2X2 AND2X2_5957 ( .A(alu__abc_42281_new_n799_), .B(alu__abc_42281_new_n797_), .Y(alu__abc_42281_new_n800_));
AND2X2 AND2X2_5958 ( .A(alu__abc_42281_new_n711_), .B(alu__abc_42281_new_n801_), .Y(alu__abc_42281_new_n802_));
AND2X2 AND2X2_5959 ( .A(alu__abc_42281_new_n800_), .B(alu__abc_42281_new_n802_), .Y(alu__abc_42281_new_n803_));
AND2X2 AND2X2_596 ( .A(_abc_44694_new_n1728_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n1729_));
AND2X2 AND2X2_5960 ( .A(alu__abc_42281_new_n803_), .B(alu__abc_42281_new_n794_), .Y(alu__abc_42281_new_n804_));
AND2X2 AND2X2_5961 ( .A(alu__abc_42281_new_n804_), .B(alu__abc_42281_new_n775_), .Y(alu__abc_42281_new_n805_));
AND2X2 AND2X2_5962 ( .A(alu__abc_42281_new_n805_), .B(alu__abc_42281_new_n721_), .Y(alu__abc_42281_new_n806_));
AND2X2 AND2X2_5963 ( .A(alu__abc_42281_new_n806_), .B(alu__abc_42281_new_n692_), .Y(alu__abc_42281_new_n807_));
AND2X2 AND2X2_5964 ( .A(alu__abc_42281_new_n807_), .B(alu__abc_42281_new_n690_), .Y(alu__abc_42281_new_n808_));
AND2X2 AND2X2_5965 ( .A(alu__abc_42281_new_n808_), .B(alu__abc_42281_new_n683_), .Y(alu__abc_42281_new_n809_));
AND2X2 AND2X2_5966 ( .A(alu__abc_42281_new_n809_), .B(alu__abc_42281_new_n681_), .Y(alu__abc_42281_new_n810_));
AND2X2 AND2X2_5967 ( .A(alu__abc_42281_new_n810_), .B(alu__abc_42281_new_n673_), .Y(alu__abc_42281_new_n811_));
AND2X2 AND2X2_5968 ( .A(alu__abc_42281_new_n811_), .B(alu__abc_42281_new_n671_), .Y(alu__abc_42281_new_n812_));
AND2X2 AND2X2_5969 ( .A(alu__abc_42281_new_n812_), .B(alu__abc_42281_new_n666_), .Y(alu__abc_42281_new_n813_));
AND2X2 AND2X2_597 ( .A(_abc_44694_new_n1727_), .B(_abc_44694_new_n1729_), .Y(_0epc_q_31_0__10_));
AND2X2 AND2X2_5970 ( .A(alu__abc_42281_new_n641_), .B(alu__abc_42281_new_n814_), .Y(alu__abc_42281_new_n815_));
AND2X2 AND2X2_5971 ( .A(alu__abc_42281_new_n662_), .B(alu__abc_42281_new_n128_), .Y(alu__abc_42281_new_n816_));
AND2X2 AND2X2_5972 ( .A(alu__abc_42281_new_n818_), .B(alu__abc_42281_new_n819_), .Y(alu__abc_42281_new_n820_));
AND2X2 AND2X2_5973 ( .A(alu__abc_42281_new_n820_), .B(alu__abc_42281_new_n815_), .Y(alu__abc_42281_new_n821_));
AND2X2 AND2X2_5974 ( .A(alu__abc_42281_new_n813_), .B(alu__abc_42281_new_n821_), .Y(alu__abc_42281_new_n822_));
AND2X2 AND2X2_5975 ( .A(alu__abc_42281_new_n822_), .B(alu__abc_42281_new_n647_), .Y(alu__abc_42281_new_n823_));
AND2X2 AND2X2_5976 ( .A(alu__abc_42281_new_n823_), .B(alu__abc_42281_new_n637_), .Y(alu__abc_42281_new_n824_));
AND2X2 AND2X2_5977 ( .A(alu__abc_42281_new_n824_), .B(alu__abc_42281_new_n630_), .Y(alu__abc_42281_new_n825_));
AND2X2 AND2X2_5978 ( .A(alu__abc_42281_new_n825_), .B(alu__abc_42281_new_n628_), .Y(alu__abc_42281_new_n826_));
AND2X2 AND2X2_5979 ( .A(alu__abc_42281_new_n826_), .B(alu_op_i_0_), .Y(alu__abc_42281_new_n827_));
AND2X2 AND2X2_598 ( .A(_abc_44694_new_n1694_), .B(pc_q_11_), .Y(_abc_44694_new_n1732_));
AND2X2 AND2X2_5980 ( .A(alu__abc_42281_new_n828_), .B(alu_c_update_o), .Y(alu_c_o));
AND2X2 AND2X2_5981 ( .A(alu__abc_42281_new_n831_), .B(alu__abc_42281_new_n830_), .Y(alu__abc_42281_new_n832_));
AND2X2 AND2X2_5982 ( .A(alu__abc_42281_new_n835_), .B(alu__abc_42281_new_n834_), .Y(alu__abc_42281_new_n836_));
AND2X2 AND2X2_5983 ( .A(alu__abc_42281_new_n833_), .B(alu__abc_42281_new_n837_), .Y(alu__abc_42281_new_n838_));
AND2X2 AND2X2_5984 ( .A(alu__abc_42281_new_n841_), .B(alu__abc_42281_new_n840_), .Y(alu__abc_42281_new_n842_));
AND2X2 AND2X2_5985 ( .A(alu__abc_42281_new_n845_), .B(alu__abc_42281_new_n844_), .Y(alu__abc_42281_new_n846_));
AND2X2 AND2X2_5986 ( .A(alu__abc_42281_new_n843_), .B(alu__abc_42281_new_n847_), .Y(alu__abc_42281_new_n848_));
AND2X2 AND2X2_5987 ( .A(alu__abc_42281_new_n839_), .B(alu__abc_42281_new_n849_), .Y(alu__abc_42281_new_n850_));
AND2X2 AND2X2_5988 ( .A(alu__abc_42281_new_n853_), .B(alu__abc_42281_new_n852_), .Y(alu__abc_42281_new_n854_));
AND2X2 AND2X2_5989 ( .A(alu__abc_42281_new_n857_), .B(alu__abc_42281_new_n856_), .Y(alu__abc_42281_new_n858_));
AND2X2 AND2X2_599 ( .A(_abc_44694_new_n1733_), .B(_abc_44694_new_n1731_), .Y(_abc_44694_new_n1734_));
AND2X2 AND2X2_5990 ( .A(alu__abc_42281_new_n855_), .B(alu__abc_42281_new_n859_), .Y(alu__abc_42281_new_n860_));
AND2X2 AND2X2_5991 ( .A(alu__abc_42281_new_n860_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n861_));
AND2X2 AND2X2_5992 ( .A(alu__abc_42281_new_n863_), .B(alu__abc_42281_new_n862_), .Y(alu__abc_42281_new_n864_));
AND2X2 AND2X2_5993 ( .A(alu__abc_42281_new_n864_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n865_));
AND2X2 AND2X2_5994 ( .A(alu__abc_42281_new_n759_), .B(alu__abc_42281_new_n866_), .Y(alu__abc_42281_new_n867_));
AND2X2 AND2X2_5995 ( .A(alu__abc_42281_new_n867_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n868_));
AND2X2 AND2X2_5996 ( .A(alu__abc_42281_new_n869_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n870_));
AND2X2 AND2X2_5997 ( .A(alu__abc_42281_new_n872_), .B(alu__abc_42281_new_n851_), .Y(alu__abc_42281_new_n873_));
AND2X2 AND2X2_5998 ( .A(alu__abc_42281_new_n379_), .B(alu__abc_42281_new_n384_), .Y(alu__abc_42281_new_n875_));
AND2X2 AND2X2_5999 ( .A(alu__abc_42281_new_n875_), .B(alu_op_i_1_), .Y(alu__abc_42281_new_n876_));
AND2X2 AND2X2_6 ( .A(_abc_44694_new_n627_), .B(opcode_q_24_), .Y(_abc_44694_new_n628_));
AND2X2 AND2X2_60 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[18] ), .Y(_abc_44694_new_n720_));
AND2X2 AND2X2_600 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1735_), .Y(_abc_44694_new_n1736_));
AND2X2 AND2X2_6000 ( .A(alu__abc_42281_new_n878_), .B(alu__abc_42281_new_n877_), .Y(alu__abc_42281_new_n879_));
AND2X2 AND2X2_6001 ( .A(alu__abc_42281_new_n882_), .B(alu__abc_42281_new_n881_), .Y(alu__abc_42281_new_n883_));
AND2X2 AND2X2_6002 ( .A(alu__abc_42281_new_n880_), .B(alu__abc_42281_new_n884_), .Y(alu__abc_42281_new_n885_));
AND2X2 AND2X2_6003 ( .A(alu__abc_42281_new_n888_), .B(alu__abc_42281_new_n887_), .Y(alu__abc_42281_new_n889_));
AND2X2 AND2X2_6004 ( .A(alu__abc_42281_new_n892_), .B(alu__abc_42281_new_n891_), .Y(alu__abc_42281_new_n893_));
AND2X2 AND2X2_6005 ( .A(alu__abc_42281_new_n890_), .B(alu__abc_42281_new_n894_), .Y(alu__abc_42281_new_n895_));
AND2X2 AND2X2_6006 ( .A(alu__abc_42281_new_n886_), .B(alu__abc_42281_new_n896_), .Y(alu__abc_42281_new_n897_));
AND2X2 AND2X2_6007 ( .A(alu__abc_42281_new_n900_), .B(alu__abc_42281_new_n899_), .Y(alu__abc_42281_new_n901_));
AND2X2 AND2X2_6008 ( .A(alu__abc_42281_new_n904_), .B(alu__abc_42281_new_n903_), .Y(alu__abc_42281_new_n905_));
AND2X2 AND2X2_6009 ( .A(alu__abc_42281_new_n902_), .B(alu__abc_42281_new_n906_), .Y(alu__abc_42281_new_n907_));
AND2X2 AND2X2_601 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_11_), .Y(_abc_44694_new_n1738_));
AND2X2 AND2X2_6010 ( .A(alu__abc_42281_new_n910_), .B(alu__abc_42281_new_n909_), .Y(alu__abc_42281_new_n911_));
AND2X2 AND2X2_6011 ( .A(alu__abc_42281_new_n914_), .B(alu__abc_42281_new_n913_), .Y(alu__abc_42281_new_n915_));
AND2X2 AND2X2_6012 ( .A(alu__abc_42281_new_n912_), .B(alu__abc_42281_new_n916_), .Y(alu__abc_42281_new_n917_));
AND2X2 AND2X2_6013 ( .A(alu__abc_42281_new_n908_), .B(alu__abc_42281_new_n918_), .Y(alu__abc_42281_new_n919_));
AND2X2 AND2X2_6014 ( .A(alu__abc_42281_new_n898_), .B(alu__abc_42281_new_n920_), .Y(alu__abc_42281_new_n921_));
AND2X2 AND2X2_6015 ( .A(alu__abc_42281_new_n922_), .B(alu__abc_42281_new_n876__bF_buf3), .Y(alu__abc_42281_new_n923_));
AND2X2 AND2X2_6016 ( .A(alu__abc_42281_new_n923_), .B(alu__abc_42281_new_n874_), .Y(alu__abc_42281_new_n924_));
AND2X2 AND2X2_6017 ( .A(alu__abc_42281_new_n378_), .B(alu__abc_42281_new_n382_), .Y(alu__abc_42281_new_n925_));
AND2X2 AND2X2_6018 ( .A(alu__abc_42281_new_n925_), .B(alu__abc_42281_new_n380_), .Y(alu__abc_42281_new_n926_));
AND2X2 AND2X2_6019 ( .A(alu__abc_42281_new_n760_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n927_));
AND2X2 AND2X2_602 ( .A(_abc_44694_new_n1708_), .B(_abc_44694_new_n1705_), .Y(_abc_44694_new_n1739_));
AND2X2 AND2X2_6020 ( .A(alu__abc_42281_new_n925_), .B(alu__abc_42281_new_n385_), .Y(alu__abc_42281_new_n928_));
AND2X2 AND2X2_6021 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n759_), .Y(alu__abc_42281_new_n929_));
AND2X2 AND2X2_6022 ( .A(alu__abc_42281_new_n289_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n931_));
AND2X2 AND2X2_6023 ( .A(alu__abc_42281_new_n931_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n932_));
AND2X2 AND2X2_6024 ( .A(alu__abc_42281_new_n932_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n933_));
AND2X2 AND2X2_6025 ( .A(alu__abc_42281_new_n378_), .B(alu_op_i_0_), .Y(alu__abc_42281_new_n934_));
AND2X2 AND2X2_6026 ( .A(alu__abc_42281_new_n875_), .B(alu__abc_42281_new_n934_), .Y(alu__abc_42281_new_n935_));
AND2X2 AND2X2_6027 ( .A(alu__abc_42281_new_n935_), .B(alu__abc_42281_new_n271__bF_buf1), .Y(alu__abc_42281_new_n936_));
AND2X2 AND2X2_6028 ( .A(alu__abc_42281_new_n933_), .B(alu__abc_42281_new_n936__bF_buf4), .Y(alu__abc_42281_new_n937_));
AND2X2 AND2X2_6029 ( .A(alu_op_i_1_), .B(alu_op_i_0_), .Y(alu__abc_42281_new_n938_));
AND2X2 AND2X2_603 ( .A(alu_op_r_7_), .B(pc_q_11_), .Y(_abc_44694_new_n1741_));
AND2X2 AND2X2_6030 ( .A(alu__abc_42281_new_n380_), .B(alu__abc_42281_new_n938_), .Y(alu__abc_42281_new_n939_));
AND2X2 AND2X2_6031 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n577_), .Y(alu__abc_42281_new_n940_));
AND2X2 AND2X2_6032 ( .A(alu__abc_42281_new_n934_), .B(alu__abc_42281_new_n385_), .Y(alu__abc_42281_new_n941_));
AND2X2 AND2X2_6033 ( .A(alu__abc_42281_new_n380_), .B(alu__abc_42281_new_n383_), .Y(alu__abc_42281_new_n942_));
AND2X2 AND2X2_6034 ( .A(alu__abc_42281_new_n943_), .B(alu__abc_42281_new_n760_), .Y(alu__abc_42281_new_n944_));
AND2X2 AND2X2_6035 ( .A(alu__abc_42281_new_n947_), .B(alu_op_i_3_), .Y(alu__abc_42281_new_n948_));
AND2X2 AND2X2_6036 ( .A(alu__abc_42281_new_n925_), .B(alu__abc_42281_new_n875_), .Y(alu__abc_42281_new_n949_));
AND2X2 AND2X2_6037 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_0_), .Y(alu__abc_42281_new_n951_));
AND2X2 AND2X2_6038 ( .A(alu__abc_42281_new_n380_), .B(alu__abc_42281_new_n934_), .Y(alu__abc_42281_new_n952_));
AND2X2 AND2X2_6039 ( .A(alu__abc_42281_new_n953_), .B(alu__abc_42281_new_n954_), .Y(alu__abc_42281_new_n955_));
AND2X2 AND2X2_604 ( .A(_abc_44694_new_n1742_), .B(_abc_44694_new_n1740_), .Y(_abc_44694_new_n1743_));
AND2X2 AND2X2_6040 ( .A(alu__abc_42281_new_n955_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n956_));
AND2X2 AND2X2_6041 ( .A(alu__abc_42281_new_n938_), .B(alu_a_i_31_), .Y(alu__abc_42281_new_n961_));
AND2X2 AND2X2_6042 ( .A(alu__abc_42281_new_n961_), .B(alu__abc_42281_new_n875_), .Y(alu__abc_42281_new_n962_));
AND2X2 AND2X2_6043 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_31_), .Y(alu__abc_42281_new_n963_));
AND2X2 AND2X2_6044 ( .A(alu__abc_42281_new_n964_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n965_));
AND2X2 AND2X2_6045 ( .A(alu_a_i_30_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n966_));
AND2X2 AND2X2_6046 ( .A(alu__abc_42281_new_n288__bF_buf0), .B(alu_a_i_29_), .Y(alu__abc_42281_new_n967_));
AND2X2 AND2X2_6047 ( .A(alu__abc_42281_new_n968_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n969_));
AND2X2 AND2X2_6048 ( .A(alu__abc_42281_new_n970_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n971_));
AND2X2 AND2X2_6049 ( .A(alu__abc_42281_new_n973_), .B(alu__abc_42281_new_n972_), .Y(alu__abc_42281_new_n974_));
AND2X2 AND2X2_605 ( .A(_abc_44694_new_n1739_), .B(_abc_44694_new_n1743_), .Y(_abc_44694_new_n1744_));
AND2X2 AND2X2_6050 ( .A(alu__abc_42281_new_n977_), .B(alu__abc_42281_new_n976_), .Y(alu__abc_42281_new_n978_));
AND2X2 AND2X2_6051 ( .A(alu__abc_42281_new_n975_), .B(alu__abc_42281_new_n979_), .Y(alu__abc_42281_new_n980_));
AND2X2 AND2X2_6052 ( .A(alu__abc_42281_new_n980_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n981_));
AND2X2 AND2X2_6053 ( .A(alu__abc_42281_new_n982_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n983_));
AND2X2 AND2X2_6054 ( .A(alu__abc_42281_new_n985_), .B(alu__abc_42281_new_n984_), .Y(alu__abc_42281_new_n986_));
AND2X2 AND2X2_6055 ( .A(alu__abc_42281_new_n989_), .B(alu__abc_42281_new_n988_), .Y(alu__abc_42281_new_n990_));
AND2X2 AND2X2_6056 ( .A(alu__abc_42281_new_n987_), .B(alu__abc_42281_new_n991_), .Y(alu__abc_42281_new_n992_));
AND2X2 AND2X2_6057 ( .A(alu__abc_42281_new_n995_), .B(alu__abc_42281_new_n994_), .Y(alu__abc_42281_new_n996_));
AND2X2 AND2X2_6058 ( .A(alu__abc_42281_new_n999_), .B(alu__abc_42281_new_n998_), .Y(alu__abc_42281_new_n1000_));
AND2X2 AND2X2_6059 ( .A(alu__abc_42281_new_n997_), .B(alu__abc_42281_new_n1001_), .Y(alu__abc_42281_new_n1002_));
AND2X2 AND2X2_606 ( .A(_abc_44694_new_n1745_), .B(_abc_44694_new_n1746_), .Y(_abc_44694_new_n1747_));
AND2X2 AND2X2_6060 ( .A(alu__abc_42281_new_n993_), .B(alu__abc_42281_new_n1003_), .Y(alu__abc_42281_new_n1004_));
AND2X2 AND2X2_6061 ( .A(alu__abc_42281_new_n1004_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1005_));
AND2X2 AND2X2_6062 ( .A(alu__abc_42281_new_n1009_), .B(alu__abc_42281_new_n1008_), .Y(alu__abc_42281_new_n1010_));
AND2X2 AND2X2_6063 ( .A(alu__abc_42281_new_n1010_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n1011_));
AND2X2 AND2X2_6064 ( .A(alu__abc_42281_new_n1013_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n1014_));
AND2X2 AND2X2_6065 ( .A(alu__abc_42281_new_n1014_), .B(alu__abc_42281_new_n1012_), .Y(alu__abc_42281_new_n1015_));
AND2X2 AND2X2_6066 ( .A(alu__abc_42281_new_n1019_), .B(alu__abc_42281_new_n1018_), .Y(alu__abc_42281_new_n1020_));
AND2X2 AND2X2_6067 ( .A(alu__abc_42281_new_n1023_), .B(alu__abc_42281_new_n1022_), .Y(alu__abc_42281_new_n1024_));
AND2X2 AND2X2_6068 ( .A(alu__abc_42281_new_n1021_), .B(alu__abc_42281_new_n1025_), .Y(alu__abc_42281_new_n1026_));
AND2X2 AND2X2_6069 ( .A(alu__abc_42281_new_n1027_), .B(alu__abc_42281_new_n1017_), .Y(alu__abc_42281_new_n1028_));
AND2X2 AND2X2_607 ( .A(_abc_44694_new_n1748_), .B(_abc_44694_new_n1194__bF_buf3), .Y(_abc_44694_new_n1749_));
AND2X2 AND2X2_6070 ( .A(alu__abc_42281_new_n1031_), .B(alu__abc_42281_new_n1030_), .Y(alu__abc_42281_new_n1032_));
AND2X2 AND2X2_6071 ( .A(alu__abc_42281_new_n1035_), .B(alu__abc_42281_new_n1034_), .Y(alu__abc_42281_new_n1036_));
AND2X2 AND2X2_6072 ( .A(alu__abc_42281_new_n1033_), .B(alu__abc_42281_new_n1037_), .Y(alu__abc_42281_new_n1038_));
AND2X2 AND2X2_6073 ( .A(alu__abc_42281_new_n1041_), .B(alu__abc_42281_new_n1040_), .Y(alu__abc_42281_new_n1042_));
AND2X2 AND2X2_6074 ( .A(alu__abc_42281_new_n1045_), .B(alu__abc_42281_new_n1044_), .Y(alu__abc_42281_new_n1046_));
AND2X2 AND2X2_6075 ( .A(alu__abc_42281_new_n1043_), .B(alu__abc_42281_new_n1047_), .Y(alu__abc_42281_new_n1048_));
AND2X2 AND2X2_6076 ( .A(alu__abc_42281_new_n1039_), .B(alu__abc_42281_new_n1049_), .Y(alu__abc_42281_new_n1050_));
AND2X2 AND2X2_6077 ( .A(alu__abc_42281_new_n1051_), .B(alu__abc_42281_new_n1029_), .Y(alu__abc_42281_new_n1052_));
AND2X2 AND2X2_6078 ( .A(alu__abc_42281_new_n1053_), .B(alu__abc_42281_new_n876__bF_buf2), .Y(alu__abc_42281_new_n1054_));
AND2X2 AND2X2_6079 ( .A(alu__abc_42281_new_n1007_), .B(alu__abc_42281_new_n1054_), .Y(alu__abc_42281_new_n1055_));
AND2X2 AND2X2_608 ( .A(_abc_44694_new_n1750_), .B(_abc_44694_new_n1340__bF_buf3), .Y(_abc_44694_new_n1751_));
AND2X2 AND2X2_6080 ( .A(alu__abc_42281_new_n1057_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n1058_));
AND2X2 AND2X2_6081 ( .A(alu__abc_42281_new_n1058_), .B(alu__abc_42281_new_n1056_), .Y(alu__abc_42281_new_n1059_));
AND2X2 AND2X2_6082 ( .A(alu__abc_42281_new_n697_), .B(alu__abc_42281_new_n1060_), .Y(alu__abc_42281_new_n1061_));
AND2X2 AND2X2_6083 ( .A(alu__abc_42281_new_n1061_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n1062_));
AND2X2 AND2X2_6084 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n575_), .Y(alu__abc_42281_new_n1063_));
AND2X2 AND2X2_6085 ( .A(alu__abc_42281_new_n576_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n1064_));
AND2X2 AND2X2_6086 ( .A(alu__abc_42281_new_n1069_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n1070_));
AND2X2 AND2X2_6087 ( .A(alu__abc_42281_new_n1070_), .B(alu__abc_42281_new_n1068_), .Y(alu__abc_42281_new_n1071_));
AND2X2 AND2X2_6088 ( .A(alu__abc_42281_new_n1014_), .B(alu__abc_42281_new_n286_), .Y(alu__abc_42281_new_n1072_));
AND2X2 AND2X2_6089 ( .A(alu__abc_42281_new_n1072_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n1073_));
AND2X2 AND2X2_609 ( .A(_abc_44694_new_n1337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n1752_));
AND2X2 AND2X2_6090 ( .A(alu__abc_42281_new_n1073_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n1074_));
AND2X2 AND2X2_6091 ( .A(alu__abc_42281_new_n1074_), .B(alu__abc_42281_new_n936__bF_buf3), .Y(alu__abc_42281_new_n1075_));
AND2X2 AND2X2_6092 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_1_), .Y(alu__abc_42281_new_n1076_));
AND2X2 AND2X2_6093 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n279_), .Y(alu__abc_42281_new_n1077_));
AND2X2 AND2X2_6094 ( .A(alu__abc_42281_new_n1084_), .B(alu__abc_42281_new_n1083_), .Y(alu__abc_42281_new_n1085_));
AND2X2 AND2X2_6095 ( .A(alu__abc_42281_new_n1085_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n1086_));
AND2X2 AND2X2_6096 ( .A(alu__abc_42281_new_n1087_), .B(alu__abc_42281_new_n1088_), .Y(alu__abc_42281_new_n1089_));
AND2X2 AND2X2_6097 ( .A(alu__abc_42281_new_n1089_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n1090_));
AND2X2 AND2X2_6098 ( .A(alu__abc_42281_new_n1091_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n1092_));
AND2X2 AND2X2_6099 ( .A(alu__abc_42281_new_n1093_), .B(alu__abc_42281_new_n1094_), .Y(alu__abc_42281_new_n1095_));
AND2X2 AND2X2_61 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[10] ), .Y(_abc_44694_new_n721_));
AND2X2 AND2X2_610 ( .A(_abc_44694_new_n1754_), .B(_abc_44694_new_n1737_), .Y(_abc_44694_new_n1755_));
AND2X2 AND2X2_6100 ( .A(alu__abc_42281_new_n1097_), .B(alu__abc_42281_new_n1098_), .Y(alu__abc_42281_new_n1099_));
AND2X2 AND2X2_6101 ( .A(alu__abc_42281_new_n1096_), .B(alu__abc_42281_new_n1100_), .Y(alu__abc_42281_new_n1101_));
AND2X2 AND2X2_6102 ( .A(alu__abc_42281_new_n1101_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n1102_));
AND2X2 AND2X2_6103 ( .A(alu__abc_42281_new_n864_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n1105_));
AND2X2 AND2X2_6104 ( .A(alu__abc_42281_new_n854_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n1106_));
AND2X2 AND2X2_6105 ( .A(alu__abc_42281_new_n1109_), .B(alu__abc_42281_new_n1110_), .Y(alu__abc_42281_new_n1111_));
AND2X2 AND2X2_6106 ( .A(alu__abc_42281_new_n1112_), .B(alu__abc_42281_new_n1108_), .Y(alu__abc_42281_new_n1113_));
AND2X2 AND2X2_6107 ( .A(alu__abc_42281_new_n1113_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n1114_));
AND2X2 AND2X2_6108 ( .A(alu__abc_42281_new_n1115_), .B(alu__abc_42281_new_n1116_), .Y(alu__abc_42281_new_n1117_));
AND2X2 AND2X2_6109 ( .A(alu__abc_42281_new_n1119_), .B(alu__abc_42281_new_n1120_), .Y(alu__abc_42281_new_n1121_));
AND2X2 AND2X2_611 ( .A(_abc_44694_new_n1522__bF_buf3), .B(epc_q_11_), .Y(_abc_44694_new_n1757_));
AND2X2 AND2X2_6110 ( .A(alu__abc_42281_new_n1118_), .B(alu__abc_42281_new_n1122_), .Y(alu__abc_42281_new_n1123_));
AND2X2 AND2X2_6111 ( .A(alu__abc_42281_new_n1123_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n1124_));
AND2X2 AND2X2_6112 ( .A(alu__abc_42281_new_n1126_), .B(alu__abc_42281_new_n876__bF_buf1), .Y(alu__abc_42281_new_n1127_));
AND2X2 AND2X2_6113 ( .A(alu__abc_42281_new_n1127_), .B(alu__abc_42281_new_n1104_), .Y(alu__abc_42281_new_n1128_));
AND2X2 AND2X2_6114 ( .A(alu__abc_42281_new_n1129_), .B(alu__abc_42281_new_n1130_), .Y(alu__abc_42281_new_n1131_));
AND2X2 AND2X2_6115 ( .A(alu__abc_42281_new_n1131_), .B(alu__abc_42281_new_n952__bF_buf2), .Y(alu__abc_42281_new_n1132_));
AND2X2 AND2X2_6116 ( .A(alu__abc_42281_new_n866_), .B(alu__abc_42281_new_n862_), .Y(alu__abc_42281_new_n1133_));
AND2X2 AND2X2_6117 ( .A(alu__abc_42281_new_n290_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n1135_));
AND2X2 AND2X2_6118 ( .A(alu__abc_42281_new_n1134_), .B(alu__abc_42281_new_n1136_), .Y(alu__abc_42281_new_n1137_));
AND2X2 AND2X2_6119 ( .A(alu__abc_42281_new_n1137_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1138_));
AND2X2 AND2X2_612 ( .A(_abc_44694_new_n1348__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_11_), .Y(_abc_44694_new_n1758_));
AND2X2 AND2X2_6120 ( .A(alu__abc_42281_new_n1138_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n1139_));
AND2X2 AND2X2_6121 ( .A(alu__abc_42281_new_n1139_), .B(alu__abc_42281_new_n936__bF_buf2), .Y(alu__abc_42281_new_n1140_));
AND2X2 AND2X2_6122 ( .A(alu__abc_42281_new_n950__bF_buf2), .B(alu_a_i_2_), .Y(alu__abc_42281_new_n1141_));
AND2X2 AND2X2_6123 ( .A(alu__abc_42281_new_n928__bF_buf2), .B(alu__abc_42281_new_n1142_), .Y(alu__abc_42281_new_n1143_));
AND2X2 AND2X2_6124 ( .A(alu__abc_42281_new_n751_), .B(alu__abc_42281_new_n941__bF_buf2), .Y(alu__abc_42281_new_n1144_));
AND2X2 AND2X2_6125 ( .A(alu__abc_42281_new_n939__bF_buf2), .B(alu__abc_42281_new_n292_), .Y(alu__abc_42281_new_n1145_));
AND2X2 AND2X2_6126 ( .A(alu__abc_42281_new_n765_), .B(alu__abc_42281_new_n926__bF_buf2), .Y(alu__abc_42281_new_n1150_));
AND2X2 AND2X2_6127 ( .A(alu__abc_42281_new_n1152_), .B(alu__abc_42281_new_n942__bF_buf2), .Y(alu__abc_42281_new_n1153_));
AND2X2 AND2X2_6128 ( .A(alu__abc_42281_new_n1153_), .B(alu__abc_42281_new_n1151_), .Y(alu__abc_42281_new_n1154_));
AND2X2 AND2X2_6129 ( .A(alu__abc_42281_new_n964_), .B(alu__abc_42281_new_n1084_), .Y(alu__abc_42281_new_n1159_));
AND2X2 AND2X2_613 ( .A(_abc_44694_new_n1207__bF_buf2), .B(_abc_44694_new_n1760_), .Y(_abc_44694_new_n1761_));
AND2X2 AND2X2_6130 ( .A(alu__abc_42281_new_n1159_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n1160_));
AND2X2 AND2X2_6131 ( .A(alu__abc_42281_new_n1161_), .B(alu__abc_42281_new_n1162_), .Y(alu__abc_42281_new_n1163_));
AND2X2 AND2X2_6132 ( .A(alu__abc_42281_new_n1163_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n1164_));
AND2X2 AND2X2_6133 ( .A(alu__abc_42281_new_n1165_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n1166_));
AND2X2 AND2X2_6134 ( .A(alu__abc_42281_new_n1167_), .B(alu__abc_42281_new_n1168_), .Y(alu__abc_42281_new_n1169_));
AND2X2 AND2X2_6135 ( .A(alu__abc_42281_new_n1171_), .B(alu__abc_42281_new_n1172_), .Y(alu__abc_42281_new_n1173_));
AND2X2 AND2X2_6136 ( .A(alu__abc_42281_new_n1170_), .B(alu__abc_42281_new_n1174_), .Y(alu__abc_42281_new_n1175_));
AND2X2 AND2X2_6137 ( .A(alu__abc_42281_new_n1175_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n1176_));
AND2X2 AND2X2_6138 ( .A(alu__abc_42281_new_n1010_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n1179_));
AND2X2 AND2X2_6139 ( .A(alu__abc_42281_new_n1020_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n1180_));
AND2X2 AND2X2_614 ( .A(_abc_44694_new_n1756_), .B(_abc_44694_new_n1761_), .Y(_abc_44694_new_n1762_));
AND2X2 AND2X2_6140 ( .A(alu__abc_42281_new_n1183_), .B(alu__abc_42281_new_n1184_), .Y(alu__abc_42281_new_n1185_));
AND2X2 AND2X2_6141 ( .A(alu__abc_42281_new_n1186_), .B(alu__abc_42281_new_n1182_), .Y(alu__abc_42281_new_n1187_));
AND2X2 AND2X2_6142 ( .A(alu__abc_42281_new_n1187_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1188_));
AND2X2 AND2X2_6143 ( .A(alu__abc_42281_new_n1189_), .B(alu__abc_42281_new_n1190_), .Y(alu__abc_42281_new_n1191_));
AND2X2 AND2X2_6144 ( .A(alu__abc_42281_new_n1193_), .B(alu__abc_42281_new_n1194_), .Y(alu__abc_42281_new_n1195_));
AND2X2 AND2X2_6145 ( .A(alu__abc_42281_new_n1192_), .B(alu__abc_42281_new_n1196_), .Y(alu__abc_42281_new_n1197_));
AND2X2 AND2X2_6146 ( .A(alu__abc_42281_new_n1197_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n1198_));
AND2X2 AND2X2_6147 ( .A(alu__abc_42281_new_n1200_), .B(alu__abc_42281_new_n876__bF_buf0), .Y(alu__abc_42281_new_n1201_));
AND2X2 AND2X2_6148 ( .A(alu__abc_42281_new_n1201_), .B(alu__abc_42281_new_n1178_), .Y(alu__abc_42281_new_n1202_));
AND2X2 AND2X2_6149 ( .A(alu__abc_42281_new_n1204_), .B(alu__abc_42281_new_n952__bF_buf1), .Y(alu__abc_42281_new_n1205_));
AND2X2 AND2X2_615 ( .A(_abc_44694_new_n1764_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n1765_));
AND2X2 AND2X2_6150 ( .A(alu__abc_42281_new_n1205_), .B(alu__abc_42281_new_n1203_), .Y(alu__abc_42281_new_n1206_));
AND2X2 AND2X2_6151 ( .A(alu__abc_42281_new_n757_), .B(alu__abc_42281_new_n926__bF_buf1), .Y(alu__abc_42281_new_n1207_));
AND2X2 AND2X2_6152 ( .A(alu__abc_42281_new_n286_), .B(alu__abc_42281_new_n1013_), .Y(alu__abc_42281_new_n1208_));
AND2X2 AND2X2_6153 ( .A(alu__abc_42281_new_n1012_), .B(alu__abc_42281_new_n1008_), .Y(alu__abc_42281_new_n1210_));
AND2X2 AND2X2_6154 ( .A(alu__abc_42281_new_n1209_), .B(alu__abc_42281_new_n1211_), .Y(alu__abc_42281_new_n1212_));
AND2X2 AND2X2_6155 ( .A(alu__abc_42281_new_n1212_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n1213_));
AND2X2 AND2X2_6156 ( .A(alu__abc_42281_new_n1213_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n1214_));
AND2X2 AND2X2_6157 ( .A(alu__abc_42281_new_n1214_), .B(alu__abc_42281_new_n936__bF_buf1), .Y(alu__abc_42281_new_n1215_));
AND2X2 AND2X2_6158 ( .A(alu__abc_42281_new_n950__bF_buf1), .B(alu_a_i_3_), .Y(alu__abc_42281_new_n1216_));
AND2X2 AND2X2_6159 ( .A(alu__abc_42281_new_n939__bF_buf1), .B(alu__abc_42281_new_n297_), .Y(alu__abc_42281_new_n1217_));
AND2X2 AND2X2_616 ( .A(_abc_44694_new_n1763_), .B(_abc_44694_new_n1765_), .Y(_0epc_q_31_0__11_));
AND2X2 AND2X2_6160 ( .A(alu__abc_42281_new_n750_), .B(alu__abc_42281_new_n941__bF_buf1), .Y(alu__abc_42281_new_n1218_));
AND2X2 AND2X2_6161 ( .A(alu__abc_42281_new_n928__bF_buf1), .B(alu__abc_42281_new_n583_), .Y(alu__abc_42281_new_n1223_));
AND2X2 AND2X2_6162 ( .A(alu__abc_42281_new_n1226_), .B(alu__abc_42281_new_n942__bF_buf1), .Y(alu__abc_42281_new_n1227_));
AND2X2 AND2X2_6163 ( .A(alu__abc_42281_new_n1227_), .B(alu__abc_42281_new_n1225_), .Y(alu__abc_42281_new_n1228_));
AND2X2 AND2X2_6164 ( .A(alu__abc_42281_new_n1234_), .B(alu__abc_42281_new_n952__bF_buf0), .Y(alu__abc_42281_new_n1235_));
AND2X2 AND2X2_6165 ( .A(alu__abc_42281_new_n1235_), .B(alu__abc_42281_new_n1233_), .Y(alu__abc_42281_new_n1236_));
AND2X2 AND2X2_6166 ( .A(alu__abc_42281_new_n1238_), .B(alu__abc_42281_new_n942__bF_buf0), .Y(alu__abc_42281_new_n1239_));
AND2X2 AND2X2_6167 ( .A(alu__abc_42281_new_n1239_), .B(alu__abc_42281_new_n1237_), .Y(alu__abc_42281_new_n1240_));
AND2X2 AND2X2_6168 ( .A(alu__abc_42281_new_n1241_), .B(alu__abc_42281_new_n1242_), .Y(alu__abc_42281_new_n1243_));
AND2X2 AND2X2_6169 ( .A(alu__abc_42281_new_n1243_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n1244_));
AND2X2 AND2X2_617 ( .A(_abc_44694_new_n1732_), .B(pc_q_12_), .Y(_abc_44694_new_n1768_));
AND2X2 AND2X2_6170 ( .A(alu__abc_42281_new_n1245_), .B(alu__abc_42281_new_n1246_), .Y(alu__abc_42281_new_n1247_));
AND2X2 AND2X2_6171 ( .A(alu__abc_42281_new_n1247_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n1248_));
AND2X2 AND2X2_6172 ( .A(alu__abc_42281_new_n1251_), .B(alu__abc_42281_new_n1252_), .Y(alu__abc_42281_new_n1253_));
AND2X2 AND2X2_6173 ( .A(alu__abc_42281_new_n1255_), .B(alu__abc_42281_new_n1256_), .Y(alu__abc_42281_new_n1257_));
AND2X2 AND2X2_6174 ( .A(alu__abc_42281_new_n1254_), .B(alu__abc_42281_new_n1258_), .Y(alu__abc_42281_new_n1259_));
AND2X2 AND2X2_6175 ( .A(alu__abc_42281_new_n1260_), .B(alu__abc_42281_new_n876__bF_buf3), .Y(alu__abc_42281_new_n1261_));
AND2X2 AND2X2_6176 ( .A(alu__abc_42281_new_n1261_), .B(alu__abc_42281_new_n1250_), .Y(alu__abc_42281_new_n1262_));
AND2X2 AND2X2_6177 ( .A(alu__abc_42281_new_n769_), .B(alu__abc_42281_new_n926__bF_buf0), .Y(alu__abc_42281_new_n1263_));
AND2X2 AND2X2_6178 ( .A(alu__abc_42281_new_n863_), .B(alu__abc_42281_new_n852_), .Y(alu__abc_42281_new_n1265_));
AND2X2 AND2X2_6179 ( .A(alu__abc_42281_new_n1266_), .B(alu__abc_42281_new_n1267_), .Y(alu__abc_42281_new_n1268_));
AND2X2 AND2X2_618 ( .A(_abc_44694_new_n1769_), .B(_abc_44694_new_n1767_), .Y(_abc_44694_new_n1770_));
AND2X2 AND2X2_6180 ( .A(alu__abc_42281_new_n1269_), .B(alu__abc_42281_new_n1264_), .Y(alu__abc_42281_new_n1270_));
AND2X2 AND2X2_6181 ( .A(alu__abc_42281_new_n1270_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n1271_));
AND2X2 AND2X2_6182 ( .A(alu__abc_42281_new_n1271_), .B(alu__abc_42281_new_n936__bF_buf0), .Y(alu__abc_42281_new_n1272_));
AND2X2 AND2X2_6183 ( .A(alu__abc_42281_new_n950__bF_buf0), .B(alu_a_i_4_), .Y(alu__abc_42281_new_n1273_));
AND2X2 AND2X2_6184 ( .A(alu__abc_42281_new_n275_), .B(alu__abc_42281_new_n941__bF_buf0), .Y(alu__abc_42281_new_n1274_));
AND2X2 AND2X2_6185 ( .A(alu__abc_42281_new_n928__bF_buf0), .B(alu__abc_42281_new_n274_), .Y(alu__abc_42281_new_n1275_));
AND2X2 AND2X2_6186 ( .A(alu__abc_42281_new_n939__bF_buf0), .B(alu__abc_42281_new_n269_), .Y(alu__abc_42281_new_n1276_));
AND2X2 AND2X2_6187 ( .A(alu__abc_42281_new_n749_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n1285_));
AND2X2 AND2X2_6188 ( .A(alu__abc_42281_new_n1287_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n1288_));
AND2X2 AND2X2_6189 ( .A(alu__abc_42281_new_n1288_), .B(alu__abc_42281_new_n1286_), .Y(alu__abc_42281_new_n1289_));
AND2X2 AND2X2_619 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1771_), .Y(_abc_44694_new_n1772_));
AND2X2 AND2X2_6190 ( .A(alu__abc_42281_new_n1293_), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n1294_));
AND2X2 AND2X2_6191 ( .A(alu__abc_42281_new_n1294_), .B(alu__abc_42281_new_n1292_), .Y(alu__abc_42281_new_n1295_));
AND2X2 AND2X2_6192 ( .A(alu__abc_42281_new_n1296_), .B(alu__abc_42281_new_n1256_), .Y(alu__abc_42281_new_n1297_));
AND2X2 AND2X2_6193 ( .A(alu__abc_42281_new_n1297_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n1298_));
AND2X2 AND2X2_6194 ( .A(alu__abc_42281_new_n1299_), .B(alu__abc_42281_new_n1300_), .Y(alu__abc_42281_new_n1301_));
AND2X2 AND2X2_6195 ( .A(alu__abc_42281_new_n1301_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n1302_));
AND2X2 AND2X2_6196 ( .A(alu__abc_42281_new_n1026_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n1305_));
AND2X2 AND2X2_6197 ( .A(alu__abc_42281_new_n1038_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n1306_));
AND2X2 AND2X2_6198 ( .A(alu__abc_42281_new_n1309_), .B(alu__abc_42281_new_n1310_), .Y(alu__abc_42281_new_n1311_));
AND2X2 AND2X2_6199 ( .A(alu__abc_42281_new_n1312_), .B(alu__abc_42281_new_n1308_), .Y(alu__abc_42281_new_n1313_));
AND2X2 AND2X2_62 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[26] ), .Y(_abc_44694_new_n723_));
AND2X2 AND2X2_620 ( .A(_abc_44694_new_n1019__bF_buf4), .B(epc_q_12_), .Y(_abc_44694_new_n1774_));
AND2X2 AND2X2_6200 ( .A(alu__abc_42281_new_n1314_), .B(alu__abc_42281_new_n876__bF_buf2), .Y(alu__abc_42281_new_n1315_));
AND2X2 AND2X2_6201 ( .A(alu__abc_42281_new_n1304_), .B(alu__abc_42281_new_n1315_), .Y(alu__abc_42281_new_n1316_));
AND2X2 AND2X2_6202 ( .A(alu__abc_42281_new_n1009_), .B(alu__abc_42281_new_n1018_), .Y(alu__abc_42281_new_n1318_));
AND2X2 AND2X2_6203 ( .A(alu__abc_42281_new_n1319_), .B(alu__abc_42281_new_n1320_), .Y(alu__abc_42281_new_n1321_));
AND2X2 AND2X2_6204 ( .A(alu__abc_42281_new_n1322_), .B(alu__abc_42281_new_n1317_), .Y(alu__abc_42281_new_n1323_));
AND2X2 AND2X2_6205 ( .A(alu__abc_42281_new_n1323_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1324_));
AND2X2 AND2X2_6206 ( .A(alu__abc_42281_new_n1324_), .B(alu__abc_42281_new_n936__bF_buf4), .Y(alu__abc_42281_new_n1325_));
AND2X2 AND2X2_6207 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_5_), .Y(alu__abc_42281_new_n1326_));
AND2X2 AND2X2_6208 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n593_), .Y(alu__abc_42281_new_n1327_));
AND2X2 AND2X2_6209 ( .A(alu__abc_42281_new_n589_), .B(alu__abc_42281_new_n941__bF_buf4), .Y(alu__abc_42281_new_n1328_));
AND2X2 AND2X2_621 ( .A(_abc_44694_new_n1706_), .B(_abc_44694_new_n1743_), .Y(_abc_44694_new_n1775_));
AND2X2 AND2X2_6210 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n264_), .Y(alu__abc_42281_new_n1330_));
AND2X2 AND2X2_6211 ( .A(alu__abc_42281_new_n1338_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n1339_));
AND2X2 AND2X2_6212 ( .A(alu__abc_42281_new_n1339_), .B(alu__abc_42281_new_n1337_), .Y(alu__abc_42281_new_n1340_));
AND2X2 AND2X2_6213 ( .A(alu__abc_42281_new_n1342_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n1343_));
AND2X2 AND2X2_6214 ( .A(alu__abc_42281_new_n1343_), .B(alu__abc_42281_new_n1341_), .Y(alu__abc_42281_new_n1344_));
AND2X2 AND2X2_6215 ( .A(alu__abc_42281_new_n742_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n1345_));
AND2X2 AND2X2_6216 ( .A(alu__abc_42281_new_n1346_), .B(alu__abc_42281_new_n1256_), .Y(alu__abc_42281_new_n1347_));
AND2X2 AND2X2_6217 ( .A(alu__abc_42281_new_n1347_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n1348_));
AND2X2 AND2X2_6218 ( .A(alu__abc_42281_new_n1349_), .B(alu__abc_42281_new_n1350_), .Y(alu__abc_42281_new_n1351_));
AND2X2 AND2X2_6219 ( .A(alu__abc_42281_new_n1351_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n1352_));
AND2X2 AND2X2_622 ( .A(_abc_44694_new_n1699_), .B(_abc_44694_new_n1775_), .Y(_abc_44694_new_n1776_));
AND2X2 AND2X2_6220 ( .A(alu__abc_42281_new_n1355_), .B(alu__abc_42281_new_n1356_), .Y(alu__abc_42281_new_n1357_));
AND2X2 AND2X2_6221 ( .A(alu__abc_42281_new_n1357_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n1358_));
AND2X2 AND2X2_6222 ( .A(alu__abc_42281_new_n1359_), .B(alu__abc_42281_new_n1360_), .Y(alu__abc_42281_new_n1361_));
AND2X2 AND2X2_6223 ( .A(alu__abc_42281_new_n1361_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n1362_));
AND2X2 AND2X2_6224 ( .A(alu__abc_42281_new_n1364_), .B(alu__abc_42281_new_n876__bF_buf1), .Y(alu__abc_42281_new_n1365_));
AND2X2 AND2X2_6225 ( .A(alu__abc_42281_new_n1365_), .B(alu__abc_42281_new_n1354_), .Y(alu__abc_42281_new_n1366_));
AND2X2 AND2X2_6226 ( .A(alu__abc_42281_new_n853_), .B(alu__abc_42281_new_n856_), .Y(alu__abc_42281_new_n1368_));
AND2X2 AND2X2_6227 ( .A(alu__abc_42281_new_n1369_), .B(alu__abc_42281_new_n1370_), .Y(alu__abc_42281_new_n1371_));
AND2X2 AND2X2_6228 ( .A(alu__abc_42281_new_n1372_), .B(alu__abc_42281_new_n1367_), .Y(alu__abc_42281_new_n1373_));
AND2X2 AND2X2_6229 ( .A(alu__abc_42281_new_n1373_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n1374_));
AND2X2 AND2X2_623 ( .A(_abc_44694_new_n1740_), .B(_abc_44694_new_n1704_), .Y(_abc_44694_new_n1777_));
AND2X2 AND2X2_6230 ( .A(alu__abc_42281_new_n1374_), .B(alu__abc_42281_new_n936__bF_buf3), .Y(alu__abc_42281_new_n1375_));
AND2X2 AND2X2_6231 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_6_), .Y(alu__abc_42281_new_n1376_));
AND2X2 AND2X2_6232 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n255_), .Y(alu__abc_42281_new_n1377_));
AND2X2 AND2X2_6233 ( .A(alu__abc_42281_new_n256_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n1378_));
AND2X2 AND2X2_6234 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n250_), .Y(alu__abc_42281_new_n1379_));
AND2X2 AND2X2_6235 ( .A(alu__abc_42281_new_n1390_), .B(alu__abc_42281_new_n942__bF_buf2), .Y(alu__abc_42281_new_n1391_));
AND2X2 AND2X2_6236 ( .A(alu__abc_42281_new_n1391_), .B(alu__abc_42281_new_n1388_), .Y(alu__abc_42281_new_n1392_));
AND2X2 AND2X2_6237 ( .A(alu__abc_42281_new_n1394_), .B(alu__abc_42281_new_n952__bF_buf2), .Y(alu__abc_42281_new_n1395_));
AND2X2 AND2X2_6238 ( .A(alu__abc_42281_new_n1395_), .B(alu__abc_42281_new_n1393_), .Y(alu__abc_42281_new_n1396_));
AND2X2 AND2X2_6239 ( .A(alu__abc_42281_new_n740_), .B(alu__abc_42281_new_n926__bF_buf2), .Y(alu__abc_42281_new_n1397_));
AND2X2 AND2X2_624 ( .A(_abc_44694_new_n1669_), .B(_abc_44694_new_n1775_), .Y(_abc_44694_new_n1780_));
AND2X2 AND2X2_6240 ( .A(alu__abc_42281_new_n1398_), .B(alu__abc_42281_new_n1256_), .Y(alu__abc_42281_new_n1399_));
AND2X2 AND2X2_6241 ( .A(alu__abc_42281_new_n1399_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n1400_));
AND2X2 AND2X2_6242 ( .A(alu__abc_42281_new_n1401_), .B(alu__abc_42281_new_n1402_), .Y(alu__abc_42281_new_n1403_));
AND2X2 AND2X2_6243 ( .A(alu__abc_42281_new_n1403_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n1404_));
AND2X2 AND2X2_6244 ( .A(alu__abc_42281_new_n1407_), .B(alu__abc_42281_new_n1408_), .Y(alu__abc_42281_new_n1409_));
AND2X2 AND2X2_6245 ( .A(alu__abc_42281_new_n1409_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n1410_));
AND2X2 AND2X2_6246 ( .A(alu__abc_42281_new_n1411_), .B(alu__abc_42281_new_n1412_), .Y(alu__abc_42281_new_n1413_));
AND2X2 AND2X2_6247 ( .A(alu__abc_42281_new_n1413_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n1414_));
AND2X2 AND2X2_6248 ( .A(alu__abc_42281_new_n1416_), .B(alu__abc_42281_new_n876__bF_buf0), .Y(alu__abc_42281_new_n1417_));
AND2X2 AND2X2_6249 ( .A(alu__abc_42281_new_n1417_), .B(alu__abc_42281_new_n1406_), .Y(alu__abc_42281_new_n1418_));
AND2X2 AND2X2_625 ( .A(_abc_44694_new_n1624_), .B(_abc_44694_new_n1780_), .Y(_abc_44694_new_n1781_));
AND2X2 AND2X2_6250 ( .A(alu__abc_42281_new_n1212_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n1419_));
AND2X2 AND2X2_6251 ( .A(alu__abc_42281_new_n1019_), .B(alu__abc_42281_new_n1022_), .Y(alu__abc_42281_new_n1420_));
AND2X2 AND2X2_6252 ( .A(alu__abc_42281_new_n1421_), .B(alu__abc_42281_new_n1422_), .Y(alu__abc_42281_new_n1423_));
AND2X2 AND2X2_6253 ( .A(alu__abc_42281_new_n1423_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n1424_));
AND2X2 AND2X2_6254 ( .A(alu__abc_42281_new_n1425_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n1426_));
AND2X2 AND2X2_6255 ( .A(alu__abc_42281_new_n1426_), .B(alu__abc_42281_new_n936__bF_buf2), .Y(alu__abc_42281_new_n1427_));
AND2X2 AND2X2_6256 ( .A(alu__abc_42281_new_n950__bF_buf2), .B(alu_a_i_7_), .Y(alu__abc_42281_new_n1428_));
AND2X2 AND2X2_6257 ( .A(alu__abc_42281_new_n587_), .B(alu__abc_42281_new_n941__bF_buf2), .Y(alu__abc_42281_new_n1429_));
AND2X2 AND2X2_6258 ( .A(alu__abc_42281_new_n928__bF_buf2), .B(alu__abc_42281_new_n597_), .Y(alu__abc_42281_new_n1430_));
AND2X2 AND2X2_6259 ( .A(alu__abc_42281_new_n939__bF_buf2), .B(alu__abc_42281_new_n258_), .Y(alu__abc_42281_new_n1431_));
AND2X2 AND2X2_626 ( .A(int32_r_10_), .B(pc_q_12_), .Y(_abc_44694_new_n1784_));
AND2X2 AND2X2_6260 ( .A(alu__abc_42281_new_n413_), .B(alu__abc_42281_new_n364_), .Y(alu__abc_42281_new_n1440_));
AND2X2 AND2X2_6261 ( .A(alu__abc_42281_new_n1442_), .B(alu__abc_42281_new_n942__bF_buf1), .Y(alu__abc_42281_new_n1443_));
AND2X2 AND2X2_6262 ( .A(alu__abc_42281_new_n1443_), .B(alu__abc_42281_new_n1441_), .Y(alu__abc_42281_new_n1444_));
AND2X2 AND2X2_6263 ( .A(alu__abc_42281_new_n1446_), .B(alu__abc_42281_new_n952__bF_buf1), .Y(alu__abc_42281_new_n1447_));
AND2X2 AND2X2_6264 ( .A(alu__abc_42281_new_n1447_), .B(alu__abc_42281_new_n1445_), .Y(alu__abc_42281_new_n1448_));
AND2X2 AND2X2_6265 ( .A(alu__abc_42281_new_n731_), .B(alu__abc_42281_new_n926__bF_buf1), .Y(alu__abc_42281_new_n1449_));
AND2X2 AND2X2_6266 ( .A(alu__abc_42281_new_n1450_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1452_));
AND2X2 AND2X2_6267 ( .A(alu__abc_42281_new_n1454_), .B(alu__abc_42281_new_n1455_), .Y(alu__abc_42281_new_n1456_));
AND2X2 AND2X2_6268 ( .A(alu__abc_42281_new_n1457_), .B(alu__abc_42281_new_n1453_), .Y(alu__abc_42281_new_n1458_));
AND2X2 AND2X2_6269 ( .A(alu__abc_42281_new_n1458_), .B(alu__abc_42281_new_n876__bF_buf3), .Y(alu__abc_42281_new_n1459_));
AND2X2 AND2X2_627 ( .A(_abc_44694_new_n1785_), .B(_abc_44694_new_n1783_), .Y(_abc_44694_new_n1786_));
AND2X2 AND2X2_6270 ( .A(alu__abc_42281_new_n857_), .B(alu__abc_42281_new_n830_), .Y(alu__abc_42281_new_n1462_));
AND2X2 AND2X2_6271 ( .A(alu__abc_42281_new_n1463_), .B(alu__abc_42281_new_n1464_), .Y(alu__abc_42281_new_n1465_));
AND2X2 AND2X2_6272 ( .A(alu__abc_42281_new_n1461_), .B(alu__abc_42281_new_n1466_), .Y(alu__abc_42281_new_n1467_));
AND2X2 AND2X2_6273 ( .A(alu__abc_42281_new_n1468_), .B(alu__abc_42281_new_n1460_), .Y(alu__abc_42281_new_n1469_));
AND2X2 AND2X2_6274 ( .A(alu__abc_42281_new_n1469_), .B(alu__abc_42281_new_n936__bF_buf1), .Y(alu__abc_42281_new_n1470_));
AND2X2 AND2X2_6275 ( .A(alu__abc_42281_new_n950__bF_buf1), .B(alu_a_i_8_), .Y(alu__abc_42281_new_n1471_));
AND2X2 AND2X2_6276 ( .A(alu__abc_42281_new_n363_), .B(alu__abc_42281_new_n941__bF_buf1), .Y(alu__abc_42281_new_n1472_));
AND2X2 AND2X2_6277 ( .A(alu__abc_42281_new_n928__bF_buf1), .B(alu__abc_42281_new_n362_), .Y(alu__abc_42281_new_n1473_));
AND2X2 AND2X2_6278 ( .A(alu__abc_42281_new_n939__bF_buf1), .B(alu__abc_42281_new_n357_), .Y(alu__abc_42281_new_n1475_));
AND2X2 AND2X2_6279 ( .A(alu__abc_42281_new_n1441_), .B(alu__abc_42281_new_n418_), .Y(alu__abc_42281_new_n1483_));
AND2X2 AND2X2_628 ( .A(_abc_44694_new_n1782_), .B(_abc_44694_new_n1786_), .Y(_abc_44694_new_n1788_));
AND2X2 AND2X2_6280 ( .A(alu__abc_42281_new_n1486_), .B(alu__abc_42281_new_n942__bF_buf0), .Y(alu__abc_42281_new_n1487_));
AND2X2 AND2X2_6281 ( .A(alu__abc_42281_new_n1487_), .B(alu__abc_42281_new_n1485_), .Y(alu__abc_42281_new_n1488_));
AND2X2 AND2X2_6282 ( .A(alu__abc_42281_new_n1490_), .B(alu__abc_42281_new_n952__bF_buf0), .Y(alu__abc_42281_new_n1491_));
AND2X2 AND2X2_6283 ( .A(alu__abc_42281_new_n1491_), .B(alu__abc_42281_new_n1489_), .Y(alu__abc_42281_new_n1492_));
AND2X2 AND2X2_6284 ( .A(alu__abc_42281_new_n728_), .B(alu__abc_42281_new_n926__bF_buf0), .Y(alu__abc_42281_new_n1493_));
AND2X2 AND2X2_6285 ( .A(alu__abc_42281_new_n1494_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1495_));
AND2X2 AND2X2_6286 ( .A(alu__abc_42281_new_n1004_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n1497_));
AND2X2 AND2X2_6287 ( .A(alu__abc_42281_new_n1050_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n1498_));
AND2X2 AND2X2_6288 ( .A(alu__abc_42281_new_n1500_), .B(alu__abc_42281_new_n876__bF_buf2), .Y(alu__abc_42281_new_n1501_));
AND2X2 AND2X2_6289 ( .A(alu__abc_42281_new_n1496_), .B(alu__abc_42281_new_n1501_), .Y(alu__abc_42281_new_n1502_));
AND2X2 AND2X2_629 ( .A(_abc_44694_new_n1789_), .B(_abc_44694_new_n1194__bF_buf2), .Y(_abc_44694_new_n1790_));
AND2X2 AND2X2_6290 ( .A(alu__abc_42281_new_n1073_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n1503_));
AND2X2 AND2X2_6291 ( .A(alu__abc_42281_new_n1023_), .B(alu__abc_42281_new_n1030_), .Y(alu__abc_42281_new_n1504_));
AND2X2 AND2X2_6292 ( .A(alu__abc_42281_new_n1505_), .B(alu__abc_42281_new_n1506_), .Y(alu__abc_42281_new_n1507_));
AND2X2 AND2X2_6293 ( .A(alu__abc_42281_new_n1508_), .B(alu__abc_42281_new_n1509_), .Y(alu__abc_42281_new_n1510_));
AND2X2 AND2X2_6294 ( .A(alu__abc_42281_new_n1510_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n1511_));
AND2X2 AND2X2_6295 ( .A(alu__abc_42281_new_n1512_), .B(alu__abc_42281_new_n936__bF_buf0), .Y(alu__abc_42281_new_n1513_));
AND2X2 AND2X2_6296 ( .A(alu__abc_42281_new_n950__bF_buf0), .B(alu_a_i_9_), .Y(alu__abc_42281_new_n1514_));
AND2X2 AND2X2_6297 ( .A(alu__abc_42281_new_n371_), .B(alu__abc_42281_new_n941__bF_buf0), .Y(alu__abc_42281_new_n1515_));
AND2X2 AND2X2_6298 ( .A(alu__abc_42281_new_n928__bF_buf0), .B(alu__abc_42281_new_n370_), .Y(alu__abc_42281_new_n1516_));
AND2X2 AND2X2_6299 ( .A(alu__abc_42281_new_n939__bF_buf0), .B(alu__abc_42281_new_n365_), .Y(alu__abc_42281_new_n1517_));
AND2X2 AND2X2_63 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[2] ), .Y(_abc_44694_new_n724_));
AND2X2 AND2X2_630 ( .A(_abc_44694_new_n1790_), .B(_abc_44694_new_n1787_), .Y(_abc_44694_new_n1791_));
AND2X2 AND2X2_6300 ( .A(alu__abc_42281_new_n413_), .B(alu__abc_42281_new_n373_), .Y(alu__abc_42281_new_n1526_));
AND2X2 AND2X2_6301 ( .A(alu__abc_42281_new_n1527_), .B(alu__abc_42281_new_n347_), .Y(alu__abc_42281_new_n1528_));
AND2X2 AND2X2_6302 ( .A(alu__abc_42281_new_n1530_), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n1531_));
AND2X2 AND2X2_6303 ( .A(alu__abc_42281_new_n1531_), .B(alu__abc_42281_new_n1529_), .Y(alu__abc_42281_new_n1532_));
AND2X2 AND2X2_6304 ( .A(alu__abc_42281_new_n775_), .B(alu__abc_42281_new_n790_), .Y(alu__abc_42281_new_n1534_));
AND2X2 AND2X2_6305 ( .A(alu__abc_42281_new_n1535_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n1536_));
AND2X2 AND2X2_6306 ( .A(alu__abc_42281_new_n1536_), .B(alu__abc_42281_new_n1533_), .Y(alu__abc_42281_new_n1537_));
AND2X2 AND2X2_6307 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n345_), .Y(alu__abc_42281_new_n1538_));
AND2X2 AND2X2_6308 ( .A(alu__abc_42281_new_n790_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n1539_));
AND2X2 AND2X2_6309 ( .A(alu__abc_42281_new_n1540_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1541_));
AND2X2 AND2X2_631 ( .A(_abc_44694_new_n1792_), .B(_abc_44694_new_n1340__bF_buf2), .Y(_abc_44694_new_n1793_));
AND2X2 AND2X2_6310 ( .A(alu__abc_42281_new_n1101_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n1543_));
AND2X2 AND2X2_6311 ( .A(alu__abc_42281_new_n1123_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n1544_));
AND2X2 AND2X2_6312 ( .A(alu__abc_42281_new_n1546_), .B(alu__abc_42281_new_n876__bF_buf1), .Y(alu__abc_42281_new_n1547_));
AND2X2 AND2X2_6313 ( .A(alu__abc_42281_new_n1547_), .B(alu__abc_42281_new_n1542_), .Y(alu__abc_42281_new_n1548_));
AND2X2 AND2X2_6314 ( .A(alu__abc_42281_new_n1138_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n1549_));
AND2X2 AND2X2_6315 ( .A(alu__abc_42281_new_n831_), .B(alu__abc_42281_new_n834_), .Y(alu__abc_42281_new_n1550_));
AND2X2 AND2X2_6316 ( .A(alu__abc_42281_new_n1551_), .B(alu__abc_42281_new_n1552_), .Y(alu__abc_42281_new_n1553_));
AND2X2 AND2X2_6317 ( .A(alu__abc_42281_new_n1554_), .B(alu__abc_42281_new_n1555_), .Y(alu__abc_42281_new_n1556_));
AND2X2 AND2X2_6318 ( .A(alu__abc_42281_new_n1556_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n1557_));
AND2X2 AND2X2_6319 ( .A(alu__abc_42281_new_n1558_), .B(alu__abc_42281_new_n936__bF_buf4), .Y(alu__abc_42281_new_n1559_));
AND2X2 AND2X2_632 ( .A(_abc_44694_new_n1337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n1794_));
AND2X2 AND2X2_6320 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_10_), .Y(alu__abc_42281_new_n1560_));
AND2X2 AND2X2_6321 ( .A(alu__abc_42281_new_n346_), .B(alu__abc_42281_new_n941__bF_buf4), .Y(alu__abc_42281_new_n1561_));
AND2X2 AND2X2_6322 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n340_), .Y(alu__abc_42281_new_n1562_));
AND2X2 AND2X2_6323 ( .A(alu__abc_42281_new_n1574_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n1575_));
AND2X2 AND2X2_6324 ( .A(alu__abc_42281_new_n1575_), .B(alu__abc_42281_new_n1572_), .Y(alu__abc_42281_new_n1576_));
AND2X2 AND2X2_6325 ( .A(alu__abc_42281_new_n1534_), .B(alu__abc_42281_new_n800_), .Y(alu__abc_42281_new_n1577_));
AND2X2 AND2X2_6326 ( .A(alu__abc_42281_new_n1579_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n1580_));
AND2X2 AND2X2_6327 ( .A(alu__abc_42281_new_n1580_), .B(alu__abc_42281_new_n1578_), .Y(alu__abc_42281_new_n1581_));
AND2X2 AND2X2_6328 ( .A(alu__abc_42281_new_n1582_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1583_));
AND2X2 AND2X2_6329 ( .A(alu__abc_42281_new_n1585_), .B(alu__abc_42281_new_n1586_), .Y(alu__abc_42281_new_n1587_));
AND2X2 AND2X2_633 ( .A(_abc_44694_new_n1796_), .B(_abc_44694_new_n1773_), .Y(_abc_44694_new_n1797_));
AND2X2 AND2X2_6330 ( .A(alu__abc_42281_new_n1588_), .B(alu__abc_42281_new_n876__bF_buf0), .Y(alu__abc_42281_new_n1589_));
AND2X2 AND2X2_6331 ( .A(alu__abc_42281_new_n1589_), .B(alu__abc_42281_new_n1584_), .Y(alu__abc_42281_new_n1590_));
AND2X2 AND2X2_6332 ( .A(alu__abc_42281_new_n800_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n1591_));
AND2X2 AND2X2_6333 ( .A(alu__abc_42281_new_n1213_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n1592_));
AND2X2 AND2X2_6334 ( .A(alu__abc_42281_new_n1031_), .B(alu__abc_42281_new_n1034_), .Y(alu__abc_42281_new_n1593_));
AND2X2 AND2X2_6335 ( .A(alu__abc_42281_new_n1594_), .B(alu__abc_42281_new_n1595_), .Y(alu__abc_42281_new_n1596_));
AND2X2 AND2X2_6336 ( .A(alu__abc_42281_new_n1597_), .B(alu__abc_42281_new_n1598_), .Y(alu__abc_42281_new_n1599_));
AND2X2 AND2X2_6337 ( .A(alu__abc_42281_new_n1599_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n1600_));
AND2X2 AND2X2_6338 ( .A(alu__abc_42281_new_n1601_), .B(alu__abc_42281_new_n936__bF_buf3), .Y(alu__abc_42281_new_n1602_));
AND2X2 AND2X2_6339 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_11_), .Y(alu__abc_42281_new_n1603_));
AND2X2 AND2X2_634 ( .A(_abc_44694_new_n1522__bF_buf2), .B(epc_q_12_), .Y(_abc_44694_new_n1799_));
AND2X2 AND2X2_6340 ( .A(alu__abc_42281_new_n354_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n1604_));
AND2X2 AND2X2_6341 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n353_), .Y(alu__abc_42281_new_n1605_));
AND2X2 AND2X2_6342 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n348_), .Y(alu__abc_42281_new_n1607_));
AND2X2 AND2X2_6343 ( .A(alu__abc_42281_new_n413_), .B(alu__abc_42281_new_n374_), .Y(alu__abc_42281_new_n1615_));
AND2X2 AND2X2_6344 ( .A(alu__abc_42281_new_n1616_), .B(alu__abc_42281_new_n312_), .Y(alu__abc_42281_new_n1618_));
AND2X2 AND2X2_6345 ( .A(alu__abc_42281_new_n1619_), .B(alu__abc_42281_new_n942__bF_buf2), .Y(alu__abc_42281_new_n1620_));
AND2X2 AND2X2_6346 ( .A(alu__abc_42281_new_n1620_), .B(alu__abc_42281_new_n1617_), .Y(alu__abc_42281_new_n1621_));
AND2X2 AND2X2_6347 ( .A(alu__abc_42281_new_n1577_), .B(alu__abc_42281_new_n792_), .Y(alu__abc_42281_new_n1623_));
AND2X2 AND2X2_6348 ( .A(alu__abc_42281_new_n1624_), .B(alu__abc_42281_new_n952__bF_buf2), .Y(alu__abc_42281_new_n1625_));
AND2X2 AND2X2_6349 ( .A(alu__abc_42281_new_n1625_), .B(alu__abc_42281_new_n1622_), .Y(alu__abc_42281_new_n1626_));
AND2X2 AND2X2_635 ( .A(_abc_44694_new_n1348__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_12_), .Y(_abc_44694_new_n1800_));
AND2X2 AND2X2_6350 ( .A(alu__abc_42281_new_n1253_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n1627_));
AND2X2 AND2X2_6351 ( .A(alu__abc_42281_new_n1247_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n1628_));
AND2X2 AND2X2_6352 ( .A(alu__abc_42281_new_n1631_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1632_));
AND2X2 AND2X2_6353 ( .A(alu__abc_42281_new_n1633_), .B(alu__abc_42281_new_n876__bF_buf3), .Y(alu__abc_42281_new_n1634_));
AND2X2 AND2X2_6354 ( .A(alu__abc_42281_new_n1634_), .B(alu__abc_42281_new_n1630_), .Y(alu__abc_42281_new_n1635_));
AND2X2 AND2X2_6355 ( .A(alu__abc_42281_new_n792_), .B(alu__abc_42281_new_n926__bF_buf2), .Y(alu__abc_42281_new_n1636_));
AND2X2 AND2X2_6356 ( .A(alu__abc_42281_new_n835_), .B(alu__abc_42281_new_n840_), .Y(alu__abc_42281_new_n1637_));
AND2X2 AND2X2_6357 ( .A(alu__abc_42281_new_n1638_), .B(alu__abc_42281_new_n1639_), .Y(alu__abc_42281_new_n1640_));
AND2X2 AND2X2_6358 ( .A(alu__abc_42281_new_n1641_), .B(alu__abc_42281_new_n1642_), .Y(alu__abc_42281_new_n1643_));
AND2X2 AND2X2_6359 ( .A(alu__abc_42281_new_n1644_), .B(alu__abc_42281_new_n1645_), .Y(alu__abc_42281_new_n1646_));
AND2X2 AND2X2_636 ( .A(_abc_44694_new_n1207__bF_buf1), .B(_abc_44694_new_n1802_), .Y(_abc_44694_new_n1803_));
AND2X2 AND2X2_6360 ( .A(alu__abc_42281_new_n1646_), .B(alu__abc_42281_new_n936__bF_buf2), .Y(alu__abc_42281_new_n1647_));
AND2X2 AND2X2_6361 ( .A(alu__abc_42281_new_n950__bF_buf2), .B(alu_a_i_12_), .Y(alu__abc_42281_new_n1648_));
AND2X2 AND2X2_6362 ( .A(alu__abc_42281_new_n311_), .B(alu__abc_42281_new_n941__bF_buf2), .Y(alu__abc_42281_new_n1649_));
AND2X2 AND2X2_6363 ( .A(alu__abc_42281_new_n928__bF_buf2), .B(alu__abc_42281_new_n310_), .Y(alu__abc_42281_new_n1650_));
AND2X2 AND2X2_6364 ( .A(alu__abc_42281_new_n939__bF_buf2), .B(alu__abc_42281_new_n305_), .Y(alu__abc_42281_new_n1651_));
AND2X2 AND2X2_6365 ( .A(alu__abc_42281_new_n1619_), .B(alu__abc_42281_new_n433_), .Y(alu__abc_42281_new_n1660_));
AND2X2 AND2X2_6366 ( .A(alu__abc_42281_new_n1663_), .B(alu__abc_42281_new_n942__bF_buf1), .Y(alu__abc_42281_new_n1664_));
AND2X2 AND2X2_6367 ( .A(alu__abc_42281_new_n1664_), .B(alu__abc_42281_new_n1662_), .Y(alu__abc_42281_new_n1665_));
AND2X2 AND2X2_6368 ( .A(alu__abc_42281_new_n1623_), .B(alu__abc_42281_new_n782_), .Y(alu__abc_42281_new_n1666_));
AND2X2 AND2X2_6369 ( .A(alu__abc_42281_new_n1668_), .B(alu__abc_42281_new_n952__bF_buf1), .Y(alu__abc_42281_new_n1669_));
AND2X2 AND2X2_637 ( .A(_abc_44694_new_n1798_), .B(_abc_44694_new_n1803_), .Y(_abc_44694_new_n1804_));
AND2X2 AND2X2_6370 ( .A(alu__abc_42281_new_n1669_), .B(alu__abc_42281_new_n1667_), .Y(alu__abc_42281_new_n1670_));
AND2X2 AND2X2_6371 ( .A(alu__abc_42281_new_n1671_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1672_));
AND2X2 AND2X2_6372 ( .A(alu__abc_42281_new_n1311_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n1674_));
AND2X2 AND2X2_6373 ( .A(alu__abc_42281_new_n1301_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n1675_));
AND2X2 AND2X2_6374 ( .A(alu__abc_42281_new_n1677_), .B(alu__abc_42281_new_n876__bF_buf2), .Y(alu__abc_42281_new_n1678_));
AND2X2 AND2X2_6375 ( .A(alu__abc_42281_new_n1673_), .B(alu__abc_42281_new_n1678_), .Y(alu__abc_42281_new_n1679_));
AND2X2 AND2X2_6376 ( .A(alu__abc_42281_new_n782_), .B(alu__abc_42281_new_n926__bF_buf1), .Y(alu__abc_42281_new_n1680_));
AND2X2 AND2X2_6377 ( .A(alu__abc_42281_new_n1035_), .B(alu__abc_42281_new_n1040_), .Y(alu__abc_42281_new_n1681_));
AND2X2 AND2X2_6378 ( .A(alu__abc_42281_new_n1682_), .B(alu__abc_42281_new_n1683_), .Y(alu__abc_42281_new_n1684_));
AND2X2 AND2X2_6379 ( .A(alu__abc_42281_new_n1685_), .B(alu__abc_42281_new_n1686_), .Y(alu__abc_42281_new_n1687_));
AND2X2 AND2X2_638 ( .A(_abc_44694_new_n1806_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n1807_));
AND2X2 AND2X2_6380 ( .A(alu__abc_42281_new_n1688_), .B(alu__abc_42281_new_n1689_), .Y(alu__abc_42281_new_n1690_));
AND2X2 AND2X2_6381 ( .A(alu__abc_42281_new_n1690_), .B(alu__abc_42281_new_n936__bF_buf1), .Y(alu__abc_42281_new_n1691_));
AND2X2 AND2X2_6382 ( .A(alu__abc_42281_new_n950__bF_buf1), .B(alu_a_i_13_), .Y(alu__abc_42281_new_n1692_));
AND2X2 AND2X2_6383 ( .A(alu__abc_42281_new_n319_), .B(alu__abc_42281_new_n941__bF_buf1), .Y(alu__abc_42281_new_n1693_));
AND2X2 AND2X2_6384 ( .A(alu__abc_42281_new_n928__bF_buf1), .B(alu__abc_42281_new_n318_), .Y(alu__abc_42281_new_n1694_));
AND2X2 AND2X2_6385 ( .A(alu__abc_42281_new_n939__bF_buf1), .B(alu__abc_42281_new_n313_), .Y(alu__abc_42281_new_n1696_));
AND2X2 AND2X2_6386 ( .A(alu__abc_42281_new_n1616_), .B(alu__abc_42281_new_n321_), .Y(alu__abc_42281_new_n1704_));
AND2X2 AND2X2_6387 ( .A(alu__abc_42281_new_n1705_), .B(alu__abc_42281_new_n329_), .Y(alu__abc_42281_new_n1707_));
AND2X2 AND2X2_6388 ( .A(alu__abc_42281_new_n1708_), .B(alu__abc_42281_new_n942__bF_buf0), .Y(alu__abc_42281_new_n1709_));
AND2X2 AND2X2_6389 ( .A(alu__abc_42281_new_n1709_), .B(alu__abc_42281_new_n1706_), .Y(alu__abc_42281_new_n1710_));
AND2X2 AND2X2_639 ( .A(_abc_44694_new_n1805_), .B(_abc_44694_new_n1807_), .Y(_0epc_q_31_0__12_));
AND2X2 AND2X2_6390 ( .A(alu__abc_42281_new_n1666_), .B(alu__abc_42281_new_n802_), .Y(alu__abc_42281_new_n1712_));
AND2X2 AND2X2_6391 ( .A(alu__abc_42281_new_n1713_), .B(alu__abc_42281_new_n952__bF_buf0), .Y(alu__abc_42281_new_n1714_));
AND2X2 AND2X2_6392 ( .A(alu__abc_42281_new_n1714_), .B(alu__abc_42281_new_n1711_), .Y(alu__abc_42281_new_n1715_));
AND2X2 AND2X2_6393 ( .A(alu__abc_42281_new_n802_), .B(alu__abc_42281_new_n926__bF_buf0), .Y(alu__abc_42281_new_n1716_));
AND2X2 AND2X2_6394 ( .A(alu__abc_42281_new_n1717_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1718_));
AND2X2 AND2X2_6395 ( .A(alu__abc_42281_new_n1351_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n1720_));
AND2X2 AND2X2_6396 ( .A(alu__abc_42281_new_n1361_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n1721_));
AND2X2 AND2X2_6397 ( .A(alu__abc_42281_new_n1723_), .B(alu__abc_42281_new_n876__bF_buf1), .Y(alu__abc_42281_new_n1724_));
AND2X2 AND2X2_6398 ( .A(alu__abc_42281_new_n1724_), .B(alu__abc_42281_new_n1719_), .Y(alu__abc_42281_new_n1725_));
AND2X2 AND2X2_6399 ( .A(alu__abc_42281_new_n841_), .B(alu__abc_42281_new_n844_), .Y(alu__abc_42281_new_n1726_));
AND2X2 AND2X2_64 ( .A(_abc_44694_new_n727_), .B(state_q_1_bF_buf4_), .Y(_abc_44694_new_n728_));
AND2X2 AND2X2_640 ( .A(_abc_44694_new_n1768_), .B(pc_q_13_), .Y(_abc_44694_new_n1810_));
AND2X2 AND2X2_6400 ( .A(alu__abc_42281_new_n1727_), .B(alu__abc_42281_new_n1728_), .Y(alu__abc_42281_new_n1729_));
AND2X2 AND2X2_6401 ( .A(alu__abc_42281_new_n1730_), .B(alu__abc_42281_new_n1731_), .Y(alu__abc_42281_new_n1732_));
AND2X2 AND2X2_6402 ( .A(alu__abc_42281_new_n1733_), .B(alu__abc_42281_new_n1734_), .Y(alu__abc_42281_new_n1735_));
AND2X2 AND2X2_6403 ( .A(alu__abc_42281_new_n1735_), .B(alu__abc_42281_new_n936__bF_buf0), .Y(alu__abc_42281_new_n1736_));
AND2X2 AND2X2_6404 ( .A(alu__abc_42281_new_n950__bF_buf0), .B(alu_a_i_14_), .Y(alu__abc_42281_new_n1737_));
AND2X2 AND2X2_6405 ( .A(alu__abc_42281_new_n928__bF_buf0), .B(alu__abc_42281_new_n327_), .Y(alu__abc_42281_new_n1738_));
AND2X2 AND2X2_6406 ( .A(alu__abc_42281_new_n328_), .B(alu__abc_42281_new_n941__bF_buf0), .Y(alu__abc_42281_new_n1739_));
AND2X2 AND2X2_6407 ( .A(alu__abc_42281_new_n939__bF_buf0), .B(alu__abc_42281_new_n322_), .Y(alu__abc_42281_new_n1741_));
AND2X2 AND2X2_6408 ( .A(alu__abc_42281_new_n1752_), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n1753_));
AND2X2 AND2X2_6409 ( .A(alu__abc_42281_new_n1753_), .B(alu__abc_42281_new_n1751_), .Y(alu__abc_42281_new_n1754_));
AND2X2 AND2X2_641 ( .A(_abc_44694_new_n1811_), .B(_abc_44694_new_n1809_), .Y(_abc_44694_new_n1812_));
AND2X2 AND2X2_6410 ( .A(alu__abc_42281_new_n721_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n1756_));
AND2X2 AND2X2_6411 ( .A(alu__abc_42281_new_n1757_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n1758_));
AND2X2 AND2X2_6412 ( .A(alu__abc_42281_new_n1755_), .B(alu__abc_42281_new_n1759_), .Y(alu__abc_42281_new_n1760_));
AND2X2 AND2X2_6413 ( .A(alu__abc_42281_new_n1761_), .B(alu__abc_42281_new_n1451_), .Y(alu__abc_42281_new_n1762_));
AND2X2 AND2X2_6414 ( .A(alu__abc_42281_new_n1409_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n1764_));
AND2X2 AND2X2_6415 ( .A(alu__abc_42281_new_n1403_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n1765_));
AND2X2 AND2X2_6416 ( .A(alu__abc_42281_new_n1767_), .B(alu__abc_42281_new_n876__bF_buf0), .Y(alu__abc_42281_new_n1768_));
AND2X2 AND2X2_6417 ( .A(alu__abc_42281_new_n1768_), .B(alu__abc_42281_new_n1763_), .Y(alu__abc_42281_new_n1769_));
AND2X2 AND2X2_6418 ( .A(alu__abc_42281_new_n1425_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n1770_));
AND2X2 AND2X2_6419 ( .A(alu__abc_42281_new_n1041_), .B(alu__abc_42281_new_n1044_), .Y(alu__abc_42281_new_n1771_));
AND2X2 AND2X2_642 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1813_), .Y(_abc_44694_new_n1814_));
AND2X2 AND2X2_6420 ( .A(alu__abc_42281_new_n1772_), .B(alu__abc_42281_new_n1773_), .Y(alu__abc_42281_new_n1774_));
AND2X2 AND2X2_6421 ( .A(alu__abc_42281_new_n1775_), .B(alu__abc_42281_new_n1776_), .Y(alu__abc_42281_new_n1777_));
AND2X2 AND2X2_6422 ( .A(alu__abc_42281_new_n1777_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n1778_));
AND2X2 AND2X2_6423 ( .A(alu__abc_42281_new_n1779_), .B(alu__abc_42281_new_n936__bF_buf4), .Y(alu__abc_42281_new_n1780_));
AND2X2 AND2X2_6424 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n335_), .Y(alu__abc_42281_new_n1781_));
AND2X2 AND2X2_6425 ( .A(alu__abc_42281_new_n336_), .B(alu__abc_42281_new_n941__bF_buf4), .Y(alu__abc_42281_new_n1782_));
AND2X2 AND2X2_6426 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_15_), .Y(alu__abc_42281_new_n1784_));
AND2X2 AND2X2_6427 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n330_), .Y(alu__abc_42281_new_n1785_));
AND2X2 AND2X2_6428 ( .A(alu__abc_42281_new_n1793_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n1794_));
AND2X2 AND2X2_6429 ( .A(alu__abc_42281_new_n1794_), .B(alu__abc_42281_new_n1792_), .Y(alu__abc_42281_new_n1795_));
AND2X2 AND2X2_643 ( .A(_abc_44694_new_n1019__bF_buf3), .B(epc_q_13_), .Y(_abc_44694_new_n1816_));
AND2X2 AND2X2_6430 ( .A(alu__abc_42281_new_n445_), .B(alu__abc_42281_new_n169_), .Y(alu__abc_42281_new_n1797_));
AND2X2 AND2X2_6431 ( .A(alu__abc_42281_new_n1798_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n1799_));
AND2X2 AND2X2_6432 ( .A(alu__abc_42281_new_n1799_), .B(alu__abc_42281_new_n1796_), .Y(alu__abc_42281_new_n1800_));
AND2X2 AND2X2_6433 ( .A(alu__abc_42281_new_n692_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n1801_));
AND2X2 AND2X2_6434 ( .A(alu__abc_42281_new_n1802_), .B(alu__abc_42281_new_n876__bF_buf3), .Y(alu__abc_42281_new_n1803_));
AND2X2 AND2X2_6435 ( .A(alu__abc_42281_new_n1804_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n1805_));
AND2X2 AND2X2_6436 ( .A(alu__abc_42281_new_n845_), .B(alu__abc_42281_new_n899_), .Y(alu__abc_42281_new_n1807_));
AND2X2 AND2X2_6437 ( .A(alu__abc_42281_new_n1808_), .B(alu__abc_42281_new_n1809_), .Y(alu__abc_42281_new_n1810_));
AND2X2 AND2X2_6438 ( .A(alu__abc_42281_new_n1806_), .B(alu__abc_42281_new_n1811_), .Y(alu__abc_42281_new_n1812_));
AND2X2 AND2X2_6439 ( .A(alu__abc_42281_new_n1812_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n1813_));
AND2X2 AND2X2_644 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_44694_new_n1818_));
AND2X2 AND2X2_6440 ( .A(alu__abc_42281_new_n1467_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n1814_));
AND2X2 AND2X2_6441 ( .A(alu__abc_42281_new_n1815_), .B(alu__abc_42281_new_n936__bF_buf3), .Y(alu__abc_42281_new_n1816_));
AND2X2 AND2X2_6442 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n162_), .Y(alu__abc_42281_new_n1817_));
AND2X2 AND2X2_6443 ( .A(alu__abc_42281_new_n935_), .B(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n1818_));
AND2X2 AND2X2_6444 ( .A(alu__abc_42281_new_n933_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n1819_));
AND2X2 AND2X2_6445 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_16_), .Y(alu__abc_42281_new_n1821_));
AND2X2 AND2X2_6446 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n167_), .Y(alu__abc_42281_new_n1822_));
AND2X2 AND2X2_6447 ( .A(alu__abc_42281_new_n168_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n1823_));
AND2X2 AND2X2_6448 ( .A(alu__abc_42281_new_n775_), .B(alu__abc_42281_new_n794_), .Y(alu__abc_42281_new_n1832_));
AND2X2 AND2X2_6449 ( .A(alu__abc_42281_new_n721_), .B(alu__abc_42281_new_n803_), .Y(alu__abc_42281_new_n1833_));
AND2X2 AND2X2_645 ( .A(_abc_44694_new_n1819_), .B(_abc_44694_new_n1817_), .Y(_abc_44694_new_n1820_));
AND2X2 AND2X2_6450 ( .A(alu__abc_42281_new_n1833_), .B(alu__abc_42281_new_n1832_), .Y(alu__abc_42281_new_n1834_));
AND2X2 AND2X2_6451 ( .A(alu__abc_42281_new_n1834_), .B(alu__abc_42281_new_n692_), .Y(alu__abc_42281_new_n1835_));
AND2X2 AND2X2_6452 ( .A(alu__abc_42281_new_n1835_), .B(alu__abc_42281_new_n690_), .Y(alu__abc_42281_new_n1836_));
AND2X2 AND2X2_6453 ( .A(alu__abc_42281_new_n1837_), .B(alu__abc_42281_new_n1838_), .Y(alu__abc_42281_new_n1839_));
AND2X2 AND2X2_6454 ( .A(alu__abc_42281_new_n1839_), .B(alu__abc_42281_new_n952__bF_buf2), .Y(alu__abc_42281_new_n1840_));
AND2X2 AND2X2_6455 ( .A(alu__abc_42281_new_n1798_), .B(alu__abc_42281_new_n450_), .Y(alu__abc_42281_new_n1841_));
AND2X2 AND2X2_6456 ( .A(alu__abc_42281_new_n1844_), .B(alu__abc_42281_new_n942__bF_buf2), .Y(alu__abc_42281_new_n1845_));
AND2X2 AND2X2_6457 ( .A(alu__abc_42281_new_n1845_), .B(alu__abc_42281_new_n1842_), .Y(alu__abc_42281_new_n1846_));
AND2X2 AND2X2_6458 ( .A(alu__abc_42281_new_n690_), .B(alu__abc_42281_new_n926__bF_buf2), .Y(alu__abc_42281_new_n1847_));
AND2X2 AND2X2_6459 ( .A(alu__abc_42281_new_n1848_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n1849_));
AND2X2 AND2X2_646 ( .A(_abc_44694_new_n1786_), .B(_abc_44694_new_n1820_), .Y(_abc_44694_new_n1823_));
AND2X2 AND2X2_6460 ( .A(alu__abc_42281_new_n950__bF_buf2), .B(alu_a_i_17_), .Y(alu__abc_42281_new_n1850_));
AND2X2 AND2X2_6461 ( .A(alu__abc_42281_new_n176_), .B(alu__abc_42281_new_n941__bF_buf2), .Y(alu__abc_42281_new_n1851_));
AND2X2 AND2X2_6462 ( .A(alu__abc_42281_new_n928__bF_buf2), .B(alu__abc_42281_new_n175_), .Y(alu__abc_42281_new_n1852_));
AND2X2 AND2X2_6463 ( .A(alu__abc_42281_new_n939__bF_buf2), .B(alu__abc_42281_new_n170_), .Y(alu__abc_42281_new_n1854_));
AND2X2 AND2X2_6464 ( .A(alu__abc_42281_new_n1045_), .B(alu__abc_42281_new_n984_), .Y(alu__abc_42281_new_n1857_));
AND2X2 AND2X2_6465 ( .A(alu__abc_42281_new_n1858_), .B(alu__abc_42281_new_n1859_), .Y(alu__abc_42281_new_n1860_));
AND2X2 AND2X2_6466 ( .A(alu__abc_42281_new_n1861_), .B(alu__abc_42281_new_n1862_), .Y(alu__abc_42281_new_n1863_));
AND2X2 AND2X2_6467 ( .A(alu__abc_42281_new_n1863_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n1864_));
AND2X2 AND2X2_6468 ( .A(alu__abc_42281_new_n1510_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n1865_));
AND2X2 AND2X2_6469 ( .A(alu__abc_42281_new_n1868_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n1869_));
AND2X2 AND2X2_647 ( .A(_abc_44694_new_n1782_), .B(_abc_44694_new_n1823_), .Y(_abc_44694_new_n1824_));
AND2X2 AND2X2_6470 ( .A(alu__abc_42281_new_n1867_), .B(alu__abc_42281_new_n1869_), .Y(alu__abc_42281_new_n1870_));
AND2X2 AND2X2_6471 ( .A(alu__abc_42281_new_n1836_), .B(alu__abc_42281_new_n683_), .Y(alu__abc_42281_new_n1876_));
AND2X2 AND2X2_6472 ( .A(alu__abc_42281_new_n1878_), .B(alu__abc_42281_new_n952__bF_buf1), .Y(alu__abc_42281_new_n1879_));
AND2X2 AND2X2_6473 ( .A(alu__abc_42281_new_n1879_), .B(alu__abc_42281_new_n1877_), .Y(alu__abc_42281_new_n1880_));
AND2X2 AND2X2_6474 ( .A(alu__abc_42281_new_n445_), .B(alu__abc_42281_new_n178_), .Y(alu__abc_42281_new_n1881_));
AND2X2 AND2X2_6475 ( .A(alu__abc_42281_new_n1882_), .B(alu__abc_42281_new_n152_), .Y(alu__abc_42281_new_n1884_));
AND2X2 AND2X2_6476 ( .A(alu__abc_42281_new_n1885_), .B(alu__abc_42281_new_n942__bF_buf1), .Y(alu__abc_42281_new_n1886_));
AND2X2 AND2X2_6477 ( .A(alu__abc_42281_new_n1886_), .B(alu__abc_42281_new_n1883_), .Y(alu__abc_42281_new_n1887_));
AND2X2 AND2X2_6478 ( .A(alu__abc_42281_new_n683_), .B(alu__abc_42281_new_n926__bF_buf1), .Y(alu__abc_42281_new_n1888_));
AND2X2 AND2X2_6479 ( .A(alu__abc_42281_new_n1889_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n1890_));
AND2X2 AND2X2_648 ( .A(_abc_44694_new_n1820_), .B(_abc_44694_new_n1784_), .Y(_abc_44694_new_n1826_));
AND2X2 AND2X2_6480 ( .A(alu__abc_42281_new_n900_), .B(alu__abc_42281_new_n903_), .Y(alu__abc_42281_new_n1891_));
AND2X2 AND2X2_6481 ( .A(alu__abc_42281_new_n1892_), .B(alu__abc_42281_new_n1893_), .Y(alu__abc_42281_new_n1894_));
AND2X2 AND2X2_6482 ( .A(alu__abc_42281_new_n1895_), .B(alu__abc_42281_new_n1896_), .Y(alu__abc_42281_new_n1897_));
AND2X2 AND2X2_6483 ( .A(alu__abc_42281_new_n1897_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n1898_));
AND2X2 AND2X2_6484 ( .A(alu__abc_42281_new_n1556_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n1899_));
AND2X2 AND2X2_6485 ( .A(alu__abc_42281_new_n1902_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n1903_));
AND2X2 AND2X2_6486 ( .A(alu__abc_42281_new_n1901_), .B(alu__abc_42281_new_n1903_), .Y(alu__abc_42281_new_n1904_));
AND2X2 AND2X2_6487 ( .A(alu__abc_42281_new_n950__bF_buf1), .B(alu_a_i_18_), .Y(alu__abc_42281_new_n1905_));
AND2X2 AND2X2_6488 ( .A(alu__abc_42281_new_n151_), .B(alu__abc_42281_new_n941__bF_buf1), .Y(alu__abc_42281_new_n1906_));
AND2X2 AND2X2_6489 ( .A(alu__abc_42281_new_n939__bF_buf1), .B(alu__abc_42281_new_n145_), .Y(alu__abc_42281_new_n1907_));
AND2X2 AND2X2_649 ( .A(_abc_44694_new_n1194__bF_buf1), .B(_abc_44694_new_n1827_), .Y(_abc_44694_new_n1828_));
AND2X2 AND2X2_6490 ( .A(alu__abc_42281_new_n928__bF_buf1), .B(alu__abc_42281_new_n150_), .Y(alu__abc_42281_new_n1908_));
AND2X2 AND2X2_6491 ( .A(alu__abc_42281_new_n1876_), .B(alu__abc_42281_new_n681_), .Y(alu__abc_42281_new_n1918_));
AND2X2 AND2X2_6492 ( .A(alu__abc_42281_new_n1919_), .B(alu__abc_42281_new_n1917_), .Y(alu__abc_42281_new_n1920_));
AND2X2 AND2X2_6493 ( .A(alu__abc_42281_new_n1920_), .B(alu__abc_42281_new_n952__bF_buf0), .Y(alu__abc_42281_new_n1921_));
AND2X2 AND2X2_6494 ( .A(alu__abc_42281_new_n1925_), .B(alu__abc_42281_new_n942__bF_buf0), .Y(alu__abc_42281_new_n1926_));
AND2X2 AND2X2_6495 ( .A(alu__abc_42281_new_n1926_), .B(alu__abc_42281_new_n1923_), .Y(alu__abc_42281_new_n1927_));
AND2X2 AND2X2_6496 ( .A(alu__abc_42281_new_n681_), .B(alu__abc_42281_new_n926__bF_buf0), .Y(alu__abc_42281_new_n1928_));
AND2X2 AND2X2_6497 ( .A(alu__abc_42281_new_n985_), .B(alu__abc_42281_new_n988_), .Y(alu__abc_42281_new_n1929_));
AND2X2 AND2X2_6498 ( .A(alu__abc_42281_new_n1930_), .B(alu__abc_42281_new_n1931_), .Y(alu__abc_42281_new_n1932_));
AND2X2 AND2X2_6499 ( .A(alu__abc_42281_new_n1933_), .B(alu__abc_42281_new_n1934_), .Y(alu__abc_42281_new_n1935_));
AND2X2 AND2X2_65 ( .A(_abc_44694_new_n719_), .B(_abc_44694_new_n728_), .Y(_abc_44694_new_n729_));
AND2X2 AND2X2_650 ( .A(_abc_44694_new_n1825_), .B(_abc_44694_new_n1828_), .Y(_abc_44694_new_n1829_));
AND2X2 AND2X2_6500 ( .A(alu__abc_42281_new_n1935_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n1936_));
AND2X2 AND2X2_6501 ( .A(alu__abc_42281_new_n1599_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n1937_));
AND2X2 AND2X2_6502 ( .A(alu__abc_42281_new_n1940_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n1941_));
AND2X2 AND2X2_6503 ( .A(alu__abc_42281_new_n1939_), .B(alu__abc_42281_new_n1941_), .Y(alu__abc_42281_new_n1942_));
AND2X2 AND2X2_6504 ( .A(alu__abc_42281_new_n1943_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n1944_));
AND2X2 AND2X2_6505 ( .A(alu__abc_42281_new_n950__bF_buf0), .B(alu_a_i_19_), .Y(alu__abc_42281_new_n1945_));
AND2X2 AND2X2_6506 ( .A(alu__abc_42281_new_n159_), .B(alu__abc_42281_new_n941__bF_buf0), .Y(alu__abc_42281_new_n1946_));
AND2X2 AND2X2_6507 ( .A(alu__abc_42281_new_n939__bF_buf0), .B(alu__abc_42281_new_n153_), .Y(alu__abc_42281_new_n1947_));
AND2X2 AND2X2_6508 ( .A(alu__abc_42281_new_n928__bF_buf0), .B(alu__abc_42281_new_n158_), .Y(alu__abc_42281_new_n1948_));
AND2X2 AND2X2_6509 ( .A(alu__abc_42281_new_n1958_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n1959_));
AND2X2 AND2X2_651 ( .A(_abc_44694_new_n1829_), .B(_abc_44694_new_n1822_), .Y(_abc_44694_new_n1830_));
AND2X2 AND2X2_6510 ( .A(alu__abc_42281_new_n1959_), .B(alu__abc_42281_new_n1957_), .Y(alu__abc_42281_new_n1960_));
AND2X2 AND2X2_6511 ( .A(alu__abc_42281_new_n445_), .B(alu__abc_42281_new_n179_), .Y(alu__abc_42281_new_n1961_));
AND2X2 AND2X2_6512 ( .A(alu__abc_42281_new_n1962_), .B(alu__abc_42281_new_n117_), .Y(alu__abc_42281_new_n1963_));
AND2X2 AND2X2_6513 ( .A(alu__abc_42281_new_n1965_), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n1966_));
AND2X2 AND2X2_6514 ( .A(alu__abc_42281_new_n1966_), .B(alu__abc_42281_new_n1964_), .Y(alu__abc_42281_new_n1967_));
AND2X2 AND2X2_6515 ( .A(alu__abc_42281_new_n673_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n1968_));
AND2X2 AND2X2_6516 ( .A(alu__abc_42281_new_n904_), .B(alu__abc_42281_new_n909_), .Y(alu__abc_42281_new_n1969_));
AND2X2 AND2X2_6517 ( .A(alu__abc_42281_new_n1970_), .B(alu__abc_42281_new_n1971_), .Y(alu__abc_42281_new_n1972_));
AND2X2 AND2X2_6518 ( .A(alu__abc_42281_new_n1973_), .B(alu__abc_42281_new_n1974_), .Y(alu__abc_42281_new_n1975_));
AND2X2 AND2X2_6519 ( .A(alu__abc_42281_new_n1975_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1976_));
AND2X2 AND2X2_652 ( .A(_abc_44694_new_n1831_), .B(_abc_44694_new_n1340__bF_buf1), .Y(_abc_44694_new_n1832_));
AND2X2 AND2X2_6520 ( .A(alu__abc_42281_new_n1643_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n1977_));
AND2X2 AND2X2_6521 ( .A(alu__abc_42281_new_n1980_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n1981_));
AND2X2 AND2X2_6522 ( .A(alu__abc_42281_new_n1979_), .B(alu__abc_42281_new_n1981_), .Y(alu__abc_42281_new_n1982_));
AND2X2 AND2X2_6523 ( .A(alu__abc_42281_new_n1983_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n1984_));
AND2X2 AND2X2_6524 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n115_), .Y(alu__abc_42281_new_n1985_));
AND2X2 AND2X2_6525 ( .A(alu__abc_42281_new_n116_), .B(alu__abc_42281_new_n941__bF_buf4), .Y(alu__abc_42281_new_n1986_));
AND2X2 AND2X2_6526 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_20_), .Y(alu__abc_42281_new_n1988_));
AND2X2 AND2X2_6527 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n110_), .Y(alu__abc_42281_new_n1989_));
AND2X2 AND2X2_6528 ( .A(alu__abc_42281_new_n1918_), .B(alu__abc_42281_new_n673_), .Y(alu__abc_42281_new_n1998_));
AND2X2 AND2X2_6529 ( .A(alu__abc_42281_new_n1998_), .B(alu__abc_42281_new_n658_), .Y(alu__abc_42281_new_n1999_));
AND2X2 AND2X2_653 ( .A(_abc_44694_new_n1337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n1833_));
AND2X2 AND2X2_6530 ( .A(alu__abc_42281_new_n2000_), .B(alu__abc_42281_new_n1997_), .Y(alu__abc_42281_new_n2001_));
AND2X2 AND2X2_6531 ( .A(alu__abc_42281_new_n2001_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n2002_));
AND2X2 AND2X2_6532 ( .A(alu__abc_42281_new_n1964_), .B(alu__abc_42281_new_n465_), .Y(alu__abc_42281_new_n2003_));
AND2X2 AND2X2_6533 ( .A(alu__abc_42281_new_n2006_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n2007_));
AND2X2 AND2X2_6534 ( .A(alu__abc_42281_new_n2007_), .B(alu__abc_42281_new_n2005_), .Y(alu__abc_42281_new_n2008_));
AND2X2 AND2X2_6535 ( .A(alu__abc_42281_new_n658_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n2009_));
AND2X2 AND2X2_6536 ( .A(alu__abc_42281_new_n2010_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2011_));
AND2X2 AND2X2_6537 ( .A(alu__abc_42281_new_n989_), .B(alu__abc_42281_new_n994_), .Y(alu__abc_42281_new_n2012_));
AND2X2 AND2X2_6538 ( .A(alu__abc_42281_new_n2013_), .B(alu__abc_42281_new_n2014_), .Y(alu__abc_42281_new_n2015_));
AND2X2 AND2X2_6539 ( .A(alu__abc_42281_new_n2016_), .B(alu__abc_42281_new_n2017_), .Y(alu__abc_42281_new_n2018_));
AND2X2 AND2X2_654 ( .A(_abc_44694_new_n1835_), .B(_abc_44694_new_n1815_), .Y(_abc_44694_new_n1836_));
AND2X2 AND2X2_6540 ( .A(alu__abc_42281_new_n2018_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n2019_));
AND2X2 AND2X2_6541 ( .A(alu__abc_42281_new_n1687_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n2020_));
AND2X2 AND2X2_6542 ( .A(alu__abc_42281_new_n2023_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n2024_));
AND2X2 AND2X2_6543 ( .A(alu__abc_42281_new_n2022_), .B(alu__abc_42281_new_n2024_), .Y(alu__abc_42281_new_n2025_));
AND2X2 AND2X2_6544 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_21_), .Y(alu__abc_42281_new_n2026_));
AND2X2 AND2X2_6545 ( .A(alu__abc_42281_new_n124_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n2027_));
AND2X2 AND2X2_6546 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n118_), .Y(alu__abc_42281_new_n2028_));
AND2X2 AND2X2_6547 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n123_), .Y(alu__abc_42281_new_n2029_));
AND2X2 AND2X2_6548 ( .A(alu__abc_42281_new_n1962_), .B(alu__abc_42281_new_n126_), .Y(alu__abc_42281_new_n2038_));
AND2X2 AND2X2_6549 ( .A(alu__abc_42281_new_n2039_), .B(alu__abc_42281_new_n134_), .Y(alu__abc_42281_new_n2041_));
AND2X2 AND2X2_655 ( .A(_abc_44694_new_n1522__bF_buf1), .B(epc_q_13_), .Y(_abc_44694_new_n1838_));
AND2X2 AND2X2_6550 ( .A(alu__abc_42281_new_n2042_), .B(alu__abc_42281_new_n942__bF_buf2), .Y(alu__abc_42281_new_n2043_));
AND2X2 AND2X2_6551 ( .A(alu__abc_42281_new_n2043_), .B(alu__abc_42281_new_n2040_), .Y(alu__abc_42281_new_n2044_));
AND2X2 AND2X2_6552 ( .A(alu__abc_42281_new_n811_), .B(alu__abc_42281_new_n665_), .Y(alu__abc_42281_new_n2046_));
AND2X2 AND2X2_6553 ( .A(alu__abc_42281_new_n2047_), .B(alu__abc_42281_new_n952__bF_buf2), .Y(alu__abc_42281_new_n2048_));
AND2X2 AND2X2_6554 ( .A(alu__abc_42281_new_n2048_), .B(alu__abc_42281_new_n2045_), .Y(alu__abc_42281_new_n2049_));
AND2X2 AND2X2_6555 ( .A(alu__abc_42281_new_n664_), .B(alu__abc_42281_new_n926__bF_buf2), .Y(alu__abc_42281_new_n2050_));
AND2X2 AND2X2_6556 ( .A(alu__abc_42281_new_n910_), .B(alu__abc_42281_new_n913_), .Y(alu__abc_42281_new_n2051_));
AND2X2 AND2X2_6557 ( .A(alu__abc_42281_new_n2052_), .B(alu__abc_42281_new_n2053_), .Y(alu__abc_42281_new_n2054_));
AND2X2 AND2X2_6558 ( .A(alu__abc_42281_new_n2055_), .B(alu__abc_42281_new_n2056_), .Y(alu__abc_42281_new_n2057_));
AND2X2 AND2X2_6559 ( .A(alu__abc_42281_new_n2057_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n2058_));
AND2X2 AND2X2_656 ( .A(_abc_44694_new_n1348__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_13_), .Y(_abc_44694_new_n1839_));
AND2X2 AND2X2_6560 ( .A(alu__abc_42281_new_n1732_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n2059_));
AND2X2 AND2X2_6561 ( .A(alu__abc_42281_new_n2062_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n2063_));
AND2X2 AND2X2_6562 ( .A(alu__abc_42281_new_n2061_), .B(alu__abc_42281_new_n2063_), .Y(alu__abc_42281_new_n2064_));
AND2X2 AND2X2_6563 ( .A(alu__abc_42281_new_n2065_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2066_));
AND2X2 AND2X2_6564 ( .A(alu__abc_42281_new_n950__bF_buf2), .B(alu_a_i_22_), .Y(alu__abc_42281_new_n2067_));
AND2X2 AND2X2_6565 ( .A(alu__abc_42281_new_n133_), .B(alu__abc_42281_new_n941__bF_buf2), .Y(alu__abc_42281_new_n2068_));
AND2X2 AND2X2_6566 ( .A(alu__abc_42281_new_n928__bF_buf2), .B(alu__abc_42281_new_n132_), .Y(alu__abc_42281_new_n2069_));
AND2X2 AND2X2_6567 ( .A(alu__abc_42281_new_n939__bF_buf2), .B(alu__abc_42281_new_n127_), .Y(alu__abc_42281_new_n2071_));
AND2X2 AND2X2_6568 ( .A(alu__abc_42281_new_n1998_), .B(alu__abc_42281_new_n665_), .Y(alu__abc_42281_new_n2080_));
AND2X2 AND2X2_6569 ( .A(alu__abc_42281_new_n2080_), .B(alu__abc_42281_new_n820_), .Y(alu__abc_42281_new_n2081_));
AND2X2 AND2X2_657 ( .A(_abc_44694_new_n1207__bF_buf0), .B(_abc_44694_new_n1841_), .Y(_abc_44694_new_n1842_));
AND2X2 AND2X2_6570 ( .A(alu__abc_42281_new_n2082_), .B(alu__abc_42281_new_n2079_), .Y(alu__abc_42281_new_n2083_));
AND2X2 AND2X2_6571 ( .A(alu__abc_42281_new_n2083_), .B(alu__abc_42281_new_n952__bF_buf1), .Y(alu__abc_42281_new_n2084_));
AND2X2 AND2X2_6572 ( .A(alu__abc_42281_new_n2088_), .B(alu__abc_42281_new_n942__bF_buf1), .Y(alu__abc_42281_new_n2089_));
AND2X2 AND2X2_6573 ( .A(alu__abc_42281_new_n2089_), .B(alu__abc_42281_new_n2087_), .Y(alu__abc_42281_new_n2090_));
AND2X2 AND2X2_6574 ( .A(alu__abc_42281_new_n820_), .B(alu__abc_42281_new_n926__bF_buf1), .Y(alu__abc_42281_new_n2091_));
AND2X2 AND2X2_6575 ( .A(alu__abc_42281_new_n995_), .B(alu__abc_42281_new_n998_), .Y(alu__abc_42281_new_n2092_));
AND2X2 AND2X2_6576 ( .A(alu__abc_42281_new_n2093_), .B(alu__abc_42281_new_n2094_), .Y(alu__abc_42281_new_n2095_));
AND2X2 AND2X2_6577 ( .A(alu__abc_42281_new_n2096_), .B(alu__abc_42281_new_n2097_), .Y(alu__abc_42281_new_n2098_));
AND2X2 AND2X2_6578 ( .A(alu__abc_42281_new_n2098_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n2099_));
AND2X2 AND2X2_6579 ( .A(alu__abc_42281_new_n1777_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n2100_));
AND2X2 AND2X2_658 ( .A(_abc_44694_new_n1837_), .B(_abc_44694_new_n1842_), .Y(_abc_44694_new_n1843_));
AND2X2 AND2X2_6580 ( .A(alu__abc_42281_new_n2103_), .B(alu__abc_42281_new_n935_), .Y(alu__abc_42281_new_n2104_));
AND2X2 AND2X2_6581 ( .A(alu__abc_42281_new_n2104_), .B(alu__abc_42281_new_n2102_), .Y(alu__abc_42281_new_n2105_));
AND2X2 AND2X2_6582 ( .A(alu__abc_42281_new_n2106_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2107_));
AND2X2 AND2X2_6583 ( .A(alu__abc_42281_new_n950__bF_buf1), .B(alu_a_i_23_), .Y(alu__abc_42281_new_n2108_));
AND2X2 AND2X2_6584 ( .A(alu__abc_42281_new_n141_), .B(alu__abc_42281_new_n941__bF_buf1), .Y(alu__abc_42281_new_n2109_));
AND2X2 AND2X2_6585 ( .A(alu__abc_42281_new_n928__bF_buf1), .B(alu__abc_42281_new_n140_), .Y(alu__abc_42281_new_n2110_));
AND2X2 AND2X2_6586 ( .A(alu__abc_42281_new_n939__bF_buf1), .B(alu__abc_42281_new_n135_), .Y(alu__abc_42281_new_n2112_));
AND2X2 AND2X2_6587 ( .A(alu__abc_42281_new_n2046_), .B(alu__abc_42281_new_n820_), .Y(alu__abc_42281_new_n2120_));
AND2X2 AND2X2_6588 ( .A(alu__abc_42281_new_n2120_), .B(alu__abc_42281_new_n650_), .Y(alu__abc_42281_new_n2122_));
AND2X2 AND2X2_6589 ( .A(alu__abc_42281_new_n2123_), .B(alu__abc_42281_new_n952__bF_buf0), .Y(alu__abc_42281_new_n2124_));
AND2X2 AND2X2_659 ( .A(_abc_44694_new_n1845_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n1846_));
AND2X2 AND2X2_6590 ( .A(alu__abc_42281_new_n2124_), .B(alu__abc_42281_new_n2121_), .Y(alu__abc_42281_new_n2125_));
AND2X2 AND2X2_6591 ( .A(alu__abc_42281_new_n2128_), .B(alu__abc_42281_new_n942__bF_buf0), .Y(alu__abc_42281_new_n2129_));
AND2X2 AND2X2_6592 ( .A(alu__abc_42281_new_n2129_), .B(alu__abc_42281_new_n2126_), .Y(alu__abc_42281_new_n2130_));
AND2X2 AND2X2_6593 ( .A(alu__abc_42281_new_n650_), .B(alu__abc_42281_new_n926__bF_buf0), .Y(alu__abc_42281_new_n2131_));
AND2X2 AND2X2_6594 ( .A(alu__abc_42281_new_n2132_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2133_));
AND2X2 AND2X2_6595 ( .A(alu__abc_42281_new_n1469_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2134_));
AND2X2 AND2X2_6596 ( .A(alu__abc_42281_new_n914_), .B(alu__abc_42281_new_n877_), .Y(alu__abc_42281_new_n2136_));
AND2X2 AND2X2_6597 ( .A(alu__abc_42281_new_n2137_), .B(alu__abc_42281_new_n2138_), .Y(alu__abc_42281_new_n2139_));
AND2X2 AND2X2_6598 ( .A(alu__abc_42281_new_n2140_), .B(alu__abc_42281_new_n2141_), .Y(alu__abc_42281_new_n2142_));
AND2X2 AND2X2_6599 ( .A(alu__abc_42281_new_n2143_), .B(alu__abc_42281_new_n936__bF_buf2), .Y(alu__abc_42281_new_n2144_));
AND2X2 AND2X2_66 ( .A(_abc_44694_new_n671_), .B(alu_p_o_3_), .Y(_abc_44694_new_n731_));
AND2X2 AND2X2_660 ( .A(_abc_44694_new_n1844_), .B(_abc_44694_new_n1846_), .Y(_0epc_q_31_0__13_));
AND2X2 AND2X2_6600 ( .A(alu__abc_42281_new_n2144_), .B(alu__abc_42281_new_n2135_), .Y(alu__abc_42281_new_n2145_));
AND2X2 AND2X2_6601 ( .A(alu__abc_42281_new_n950__bF_buf0), .B(alu_a_i_24_), .Y(alu__abc_42281_new_n2146_));
AND2X2 AND2X2_6602 ( .A(alu__abc_42281_new_n195_), .B(alu__abc_42281_new_n941__bF_buf0), .Y(alu__abc_42281_new_n2147_));
AND2X2 AND2X2_6603 ( .A(alu__abc_42281_new_n928__bF_buf0), .B(alu__abc_42281_new_n194_), .Y(alu__abc_42281_new_n2148_));
AND2X2 AND2X2_6604 ( .A(alu__abc_42281_new_n939__bF_buf0), .B(alu__abc_42281_new_n189_), .Y(alu__abc_42281_new_n2149_));
AND2X2 AND2X2_6605 ( .A(alu__abc_42281_new_n2122_), .B(alu__abc_42281_new_n671_), .Y(alu__abc_42281_new_n2159_));
AND2X2 AND2X2_6606 ( .A(alu__abc_42281_new_n2161_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n2162_));
AND2X2 AND2X2_6607 ( .A(alu__abc_42281_new_n2162_), .B(alu__abc_42281_new_n2160_), .Y(alu__abc_42281_new_n2163_));
AND2X2 AND2X2_6608 ( .A(alu__abc_42281_new_n2128_), .B(alu__abc_42281_new_n489_), .Y(alu__abc_42281_new_n2164_));
AND2X2 AND2X2_6609 ( .A(alu__abc_42281_new_n2167_), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n2168_));
AND2X2 AND2X2_661 ( .A(_abc_44694_new_n1810_), .B(pc_q_14_), .Y(_abc_44694_new_n1849_));
AND2X2 AND2X2_6610 ( .A(alu__abc_42281_new_n2168_), .B(alu__abc_42281_new_n2166_), .Y(alu__abc_42281_new_n2169_));
AND2X2 AND2X2_6611 ( .A(alu__abc_42281_new_n671_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n2170_));
AND2X2 AND2X2_6612 ( .A(alu__abc_42281_new_n2171_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2172_));
AND2X2 AND2X2_6613 ( .A(alu__abc_42281_new_n1512_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2173_));
AND2X2 AND2X2_6614 ( .A(alu__abc_42281_new_n999_), .B(alu__abc_42281_new_n972_), .Y(alu__abc_42281_new_n2174_));
AND2X2 AND2X2_6615 ( .A(alu__abc_42281_new_n2175_), .B(alu__abc_42281_new_n2176_), .Y(alu__abc_42281_new_n2177_));
AND2X2 AND2X2_6616 ( .A(alu__abc_42281_new_n2177_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n2178_));
AND2X2 AND2X2_6617 ( .A(alu__abc_42281_new_n2015_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n2179_));
AND2X2 AND2X2_6618 ( .A(alu__abc_42281_new_n2182_), .B(alu__abc_42281_new_n2181_), .Y(alu__abc_42281_new_n2183_));
AND2X2 AND2X2_6619 ( .A(alu__abc_42281_new_n2183_), .B(alu__abc_42281_new_n936__bF_buf1), .Y(alu__abc_42281_new_n2184_));
AND2X2 AND2X2_662 ( .A(_abc_44694_new_n1850_), .B(_abc_44694_new_n1848_), .Y(_abc_44694_new_n1851_));
AND2X2 AND2X2_6620 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_25_), .Y(alu__abc_42281_new_n2185_));
AND2X2 AND2X2_6621 ( .A(alu__abc_42281_new_n187_), .B(alu__abc_42281_new_n941__bF_buf4), .Y(alu__abc_42281_new_n2186_));
AND2X2 AND2X2_6622 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n186_), .Y(alu__abc_42281_new_n2187_));
AND2X2 AND2X2_6623 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n181_), .Y(alu__abc_42281_new_n2188_));
AND2X2 AND2X2_6624 ( .A(alu__abc_42281_new_n2081_), .B(alu__abc_42281_new_n650_), .Y(alu__abc_42281_new_n2199_));
AND2X2 AND2X2_6625 ( .A(alu__abc_42281_new_n2199_), .B(alu__abc_42281_new_n671_), .Y(alu__abc_42281_new_n2200_));
AND2X2 AND2X2_6626 ( .A(alu__abc_42281_new_n2200_), .B(alu__abc_42281_new_n815_), .Y(alu__abc_42281_new_n2201_));
AND2X2 AND2X2_6627 ( .A(alu__abc_42281_new_n2202_), .B(alu__abc_42281_new_n2198_), .Y(alu__abc_42281_new_n2203_));
AND2X2 AND2X2_6628 ( .A(alu__abc_42281_new_n2203_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n2204_));
AND2X2 AND2X2_6629 ( .A(alu__abc_42281_new_n2128_), .B(alu__abc_42281_new_n490_), .Y(alu__abc_42281_new_n2205_));
AND2X2 AND2X2_663 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1852_), .Y(_abc_44694_new_n1853_));
AND2X2 AND2X2_6630 ( .A(alu__abc_42281_new_n2209_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n2210_));
AND2X2 AND2X2_6631 ( .A(alu__abc_42281_new_n2210_), .B(alu__abc_42281_new_n2207_), .Y(alu__abc_42281_new_n2211_));
AND2X2 AND2X2_6632 ( .A(alu__abc_42281_new_n815_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n2212_));
AND2X2 AND2X2_6633 ( .A(alu__abc_42281_new_n2213_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2214_));
AND2X2 AND2X2_6634 ( .A(alu__abc_42281_new_n878_), .B(alu__abc_42281_new_n881_), .Y(alu__abc_42281_new_n2215_));
AND2X2 AND2X2_6635 ( .A(alu__abc_42281_new_n2216_), .B(alu__abc_42281_new_n2217_), .Y(alu__abc_42281_new_n2218_));
AND2X2 AND2X2_6636 ( .A(alu__abc_42281_new_n2218_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n2219_));
AND2X2 AND2X2_6637 ( .A(alu__abc_42281_new_n2054_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n2220_));
AND2X2 AND2X2_6638 ( .A(alu__abc_42281_new_n2223_), .B(alu__abc_42281_new_n2222_), .Y(alu__abc_42281_new_n2224_));
AND2X2 AND2X2_6639 ( .A(alu__abc_42281_new_n2224_), .B(alu__abc_42281_new_n936__bF_buf0), .Y(alu__abc_42281_new_n2225_));
AND2X2 AND2X2_664 ( .A(_abc_44694_new_n1019__bF_buf2), .B(epc_q_14_), .Y(_abc_44694_new_n1855_));
AND2X2 AND2X2_6640 ( .A(alu__abc_42281_new_n1558_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2226_));
AND2X2 AND2X2_6641 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_26_), .Y(alu__abc_42281_new_n2227_));
AND2X2 AND2X2_6642 ( .A(alu__abc_42281_new_n204_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n2228_));
AND2X2 AND2X2_6643 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n198_), .Y(alu__abc_42281_new_n2229_));
AND2X2 AND2X2_6644 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n203_), .Y(alu__abc_42281_new_n2230_));
AND2X2 AND2X2_6645 ( .A(alu__abc_42281_new_n2159_), .B(alu__abc_42281_new_n815_), .Y(alu__abc_42281_new_n2240_));
AND2X2 AND2X2_6646 ( .A(alu__abc_42281_new_n2201_), .B(alu__abc_42281_new_n646_), .Y(alu__abc_42281_new_n2242_));
AND2X2 AND2X2_6647 ( .A(alu__abc_42281_new_n2243_), .B(alu__abc_42281_new_n2241_), .Y(alu__abc_42281_new_n2244_));
AND2X2 AND2X2_6648 ( .A(alu__abc_42281_new_n2244_), .B(alu__abc_42281_new_n952__bF_buf2), .Y(alu__abc_42281_new_n2245_));
AND2X2 AND2X2_6649 ( .A(alu__abc_42281_new_n646_), .B(alu__abc_42281_new_n926__bF_buf2), .Y(alu__abc_42281_new_n2246_));
AND2X2 AND2X2_665 ( .A(_abc_44694_new_n1827_), .B(_abc_44694_new_n1819_), .Y(_abc_44694_new_n1856_));
AND2X2 AND2X2_6650 ( .A(alu__abc_42281_new_n2207_), .B(alu__abc_42281_new_n2247_), .Y(alu__abc_42281_new_n2248_));
AND2X2 AND2X2_6651 ( .A(alu__abc_42281_new_n2251_), .B(alu__abc_42281_new_n942__bF_buf2), .Y(alu__abc_42281_new_n2252_));
AND2X2 AND2X2_6652 ( .A(alu__abc_42281_new_n2252_), .B(alu__abc_42281_new_n2250_), .Y(alu__abc_42281_new_n2253_));
AND2X2 AND2X2_6653 ( .A(alu__abc_42281_new_n2254_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2255_));
AND2X2 AND2X2_6654 ( .A(alu__abc_42281_new_n1601_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2256_));
AND2X2 AND2X2_6655 ( .A(alu__abc_42281_new_n950__bF_buf2), .B(alu_a_i_27_), .Y(alu__abc_42281_new_n2257_));
AND2X2 AND2X2_6656 ( .A(alu__abc_42281_new_n928__bF_buf2), .B(alu__abc_42281_new_n211_), .Y(alu__abc_42281_new_n2258_));
AND2X2 AND2X2_6657 ( .A(alu__abc_42281_new_n212_), .B(alu__abc_42281_new_n941__bF_buf2), .Y(alu__abc_42281_new_n2259_));
AND2X2 AND2X2_6658 ( .A(alu__abc_42281_new_n939__bF_buf2), .B(alu__abc_42281_new_n206_), .Y(alu__abc_42281_new_n2261_));
AND2X2 AND2X2_6659 ( .A(alu__abc_42281_new_n973_), .B(alu__abc_42281_new_n976_), .Y(alu__abc_42281_new_n2265_));
AND2X2 AND2X2_666 ( .A(_abc_44694_new_n1825_), .B(_abc_44694_new_n1856_), .Y(_abc_44694_new_n1857_));
AND2X2 AND2X2_6660 ( .A(alu__abc_42281_new_n2266_), .B(alu__abc_42281_new_n2267_), .Y(alu__abc_42281_new_n2268_));
AND2X2 AND2X2_6661 ( .A(alu__abc_42281_new_n2268_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n2269_));
AND2X2 AND2X2_6662 ( .A(alu__abc_42281_new_n2095_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n2270_));
AND2X2 AND2X2_6663 ( .A(alu__abc_42281_new_n2272_), .B(alu__abc_42281_new_n936__bF_buf4), .Y(alu__abc_42281_new_n2273_));
AND2X2 AND2X2_6664 ( .A(alu__abc_42281_new_n2273_), .B(alu__abc_42281_new_n2264_), .Y(alu__abc_42281_new_n2274_));
AND2X2 AND2X2_6665 ( .A(alu__abc_42281_new_n2242_), .B(alu__abc_42281_new_n639_), .Y(alu__abc_42281_new_n2282_));
AND2X2 AND2X2_6666 ( .A(alu__abc_42281_new_n2283_), .B(alu__abc_42281_new_n2281_), .Y(alu__abc_42281_new_n2284_));
AND2X2 AND2X2_6667 ( .A(alu__abc_42281_new_n2284_), .B(alu__abc_42281_new_n952__bF_buf1), .Y(alu__abc_42281_new_n2285_));
AND2X2 AND2X2_6668 ( .A(alu__abc_42281_new_n495_), .B(alu__abc_42281_new_n223_), .Y(alu__abc_42281_new_n2287_));
AND2X2 AND2X2_6669 ( .A(alu__abc_42281_new_n2288_), .B(alu__abc_42281_new_n942__bF_buf1), .Y(alu__abc_42281_new_n2289_));
AND2X2 AND2X2_667 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_44694_new_n1860_));
AND2X2 AND2X2_6670 ( .A(alu__abc_42281_new_n2289_), .B(alu__abc_42281_new_n2286_), .Y(alu__abc_42281_new_n2290_));
AND2X2 AND2X2_6671 ( .A(alu__abc_42281_new_n639_), .B(alu__abc_42281_new_n926__bF_buf1), .Y(alu__abc_42281_new_n2291_));
AND2X2 AND2X2_6672 ( .A(alu__abc_42281_new_n2292_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2293_));
AND2X2 AND2X2_6673 ( .A(alu__abc_42281_new_n882_), .B(alu__abc_42281_new_n887_), .Y(alu__abc_42281_new_n2295_));
AND2X2 AND2X2_6674 ( .A(alu__abc_42281_new_n2295_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n2296_));
AND2X2 AND2X2_6675 ( .A(alu__abc_42281_new_n2215_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n2297_));
AND2X2 AND2X2_6676 ( .A(alu__abc_42281_new_n2300_), .B(alu__abc_42281_new_n2299_), .Y(alu__abc_42281_new_n2301_));
AND2X2 AND2X2_6677 ( .A(alu__abc_42281_new_n2302_), .B(alu__abc_42281_new_n936__bF_buf3), .Y(alu__abc_42281_new_n2303_));
AND2X2 AND2X2_6678 ( .A(alu__abc_42281_new_n2303_), .B(alu__abc_42281_new_n2294_), .Y(alu__abc_42281_new_n2304_));
AND2X2 AND2X2_6679 ( .A(alu__abc_42281_new_n1646_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2305_));
AND2X2 AND2X2_668 ( .A(_abc_44694_new_n1861_), .B(_abc_44694_new_n1859_), .Y(_abc_44694_new_n1862_));
AND2X2 AND2X2_6680 ( .A(alu__abc_42281_new_n950__bF_buf1), .B(alu_a_i_28_), .Y(alu__abc_42281_new_n2306_));
AND2X2 AND2X2_6681 ( .A(alu__abc_42281_new_n222_), .B(alu__abc_42281_new_n941__bF_buf1), .Y(alu__abc_42281_new_n2307_));
AND2X2 AND2X2_6682 ( .A(alu__abc_42281_new_n928__bF_buf1), .B(alu__abc_42281_new_n221_), .Y(alu__abc_42281_new_n2308_));
AND2X2 AND2X2_6683 ( .A(alu__abc_42281_new_n939__bF_buf1), .B(alu__abc_42281_new_n216_), .Y(alu__abc_42281_new_n2309_));
AND2X2 AND2X2_6684 ( .A(alu__abc_42281_new_n2240_), .B(alu__abc_42281_new_n647_), .Y(alu__abc_42281_new_n2319_));
AND2X2 AND2X2_6685 ( .A(alu__abc_42281_new_n2319_), .B(alu__abc_42281_new_n637_), .Y(alu__abc_42281_new_n2321_));
AND2X2 AND2X2_6686 ( .A(alu__abc_42281_new_n2322_), .B(alu__abc_42281_new_n952__bF_buf0), .Y(alu__abc_42281_new_n2323_));
AND2X2 AND2X2_6687 ( .A(alu__abc_42281_new_n2323_), .B(alu__abc_42281_new_n2320_), .Y(alu__abc_42281_new_n2324_));
AND2X2 AND2X2_6688 ( .A(alu__abc_42281_new_n2288_), .B(alu__abc_42281_new_n501_), .Y(alu__abc_42281_new_n2325_));
AND2X2 AND2X2_6689 ( .A(alu__abc_42281_new_n2328_), .B(alu__abc_42281_new_n942__bF_buf0), .Y(alu__abc_42281_new_n2329_));
AND2X2 AND2X2_669 ( .A(_abc_44694_new_n1858_), .B(_abc_44694_new_n1862_), .Y(_abc_44694_new_n1863_));
AND2X2 AND2X2_6690 ( .A(alu__abc_42281_new_n2329_), .B(alu__abc_42281_new_n2326_), .Y(alu__abc_42281_new_n2330_));
AND2X2 AND2X2_6691 ( .A(alu__abc_42281_new_n637_), .B(alu__abc_42281_new_n926__bF_buf0), .Y(alu__abc_42281_new_n2331_));
AND2X2 AND2X2_6692 ( .A(alu__abc_42281_new_n2332_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2333_));
AND2X2 AND2X2_6693 ( .A(alu__abc_42281_new_n1690_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2334_));
AND2X2 AND2X2_6694 ( .A(alu__abc_42281_new_n977_), .B(alu__abc_42281_new_n2335_), .Y(alu__abc_42281_new_n2336_));
AND2X2 AND2X2_6695 ( .A(alu__abc_42281_new_n2337_), .B(alu__abc_42281_new_n2338_), .Y(alu__abc_42281_new_n2339_));
AND2X2 AND2X2_6696 ( .A(alu__abc_42281_new_n2340_), .B(alu__abc_42281_new_n2341_), .Y(alu__abc_42281_new_n2342_));
AND2X2 AND2X2_6697 ( .A(alu__abc_42281_new_n2343_), .B(alu__abc_42281_new_n2344_), .Y(alu__abc_42281_new_n2345_));
AND2X2 AND2X2_6698 ( .A(alu__abc_42281_new_n2345_), .B(alu__abc_42281_new_n936__bF_buf2), .Y(alu__abc_42281_new_n2346_));
AND2X2 AND2X2_6699 ( .A(alu__abc_42281_new_n950__bF_buf0), .B(alu_a_i_29_), .Y(alu__abc_42281_new_n2347_));
AND2X2 AND2X2_67 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[3] ), .Y(_abc_44694_new_n732_));
AND2X2 AND2X2_670 ( .A(_abc_44694_new_n1865_), .B(_abc_44694_new_n1194__bF_buf0), .Y(_abc_44694_new_n1866_));
AND2X2 AND2X2_6700 ( .A(alu__abc_42281_new_n230_), .B(alu__abc_42281_new_n941__bF_buf0), .Y(alu__abc_42281_new_n2348_));
AND2X2 AND2X2_6701 ( .A(alu__abc_42281_new_n928__bF_buf0), .B(alu__abc_42281_new_n229_), .Y(alu__abc_42281_new_n2349_));
AND2X2 AND2X2_6702 ( .A(alu__abc_42281_new_n939__bF_buf0), .B(alu__abc_42281_new_n224_), .Y(alu__abc_42281_new_n2350_));
AND2X2 AND2X2_6703 ( .A(alu__abc_42281_new_n2321_), .B(alu__abc_42281_new_n630_), .Y(alu__abc_42281_new_n2360_));
AND2X2 AND2X2_6704 ( .A(alu__abc_42281_new_n2362_), .B(alu__abc_42281_new_n952__bF_buf4), .Y(alu__abc_42281_new_n2363_));
AND2X2 AND2X2_6705 ( .A(alu__abc_42281_new_n2363_), .B(alu__abc_42281_new_n2361_), .Y(alu__abc_42281_new_n2364_));
AND2X2 AND2X2_6706 ( .A(alu__abc_42281_new_n2366_), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n2367_));
AND2X2 AND2X2_6707 ( .A(alu__abc_42281_new_n2367_), .B(alu__abc_42281_new_n2365_), .Y(alu__abc_42281_new_n2368_));
AND2X2 AND2X2_6708 ( .A(alu__abc_42281_new_n630_), .B(alu__abc_42281_new_n926__bF_buf4), .Y(alu__abc_42281_new_n2369_));
AND2X2 AND2X2_6709 ( .A(alu__abc_42281_new_n2370_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2371_));
AND2X2 AND2X2_671 ( .A(_abc_44694_new_n1866_), .B(_abc_44694_new_n1864_), .Y(_abc_44694_new_n1867_));
AND2X2 AND2X2_6710 ( .A(alu__abc_42281_new_n888_), .B(alu__abc_42281_new_n891_), .Y(alu__abc_42281_new_n2372_));
AND2X2 AND2X2_6711 ( .A(alu__abc_42281_new_n2372_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n2373_));
AND2X2 AND2X2_6712 ( .A(alu__abc_42281_new_n2295_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n2374_));
AND2X2 AND2X2_6713 ( .A(alu__abc_42281_new_n2377_), .B(alu__abc_42281_new_n2376_), .Y(alu__abc_42281_new_n2378_));
AND2X2 AND2X2_6714 ( .A(alu__abc_42281_new_n2380_), .B(alu__abc_42281_new_n2379_), .Y(alu__abc_42281_new_n2381_));
AND2X2 AND2X2_6715 ( .A(alu__abc_42281_new_n2381_), .B(alu__abc_42281_new_n936__bF_buf1), .Y(alu__abc_42281_new_n2382_));
AND2X2 AND2X2_6716 ( .A(alu__abc_42281_new_n1735_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2383_));
AND2X2 AND2X2_6717 ( .A(alu__abc_42281_new_n950__bF_buf4), .B(alu_a_i_30_), .Y(alu__abc_42281_new_n2384_));
AND2X2 AND2X2_6718 ( .A(alu__abc_42281_new_n239_), .B(alu__abc_42281_new_n941__bF_buf4), .Y(alu__abc_42281_new_n2385_));
AND2X2 AND2X2_6719 ( .A(alu__abc_42281_new_n939__bF_buf4), .B(alu__abc_42281_new_n233_), .Y(alu__abc_42281_new_n2386_));
AND2X2 AND2X2_672 ( .A(_abc_44694_new_n1868_), .B(_abc_44694_new_n1340__bF_buf0), .Y(_abc_44694_new_n1869_));
AND2X2 AND2X2_6720 ( .A(alu__abc_42281_new_n928__bF_buf4), .B(alu__abc_42281_new_n238_), .Y(alu__abc_42281_new_n2387_));
AND2X2 AND2X2_6721 ( .A(alu__abc_42281_new_n2398_), .B(alu__abc_42281_new_n952__bF_buf3), .Y(alu__abc_42281_new_n2399_));
AND2X2 AND2X2_6722 ( .A(alu__abc_42281_new_n2397_), .B(alu__abc_42281_new_n2399_), .Y(alu__abc_42281_new_n2400_));
AND2X2 AND2X2_6723 ( .A(alu__abc_42281_new_n628_), .B(alu__abc_42281_new_n926__bF_buf3), .Y(alu__abc_42281_new_n2401_));
AND2X2 AND2X2_6724 ( .A(alu__abc_42281_new_n2402_), .B(alu__abc_42281_new_n2403_), .Y(alu__abc_42281_new_n2404_));
AND2X2 AND2X2_6725 ( .A(alu__abc_42281_new_n2404_), .B(alu__abc_42281_new_n942__bF_buf3), .Y(alu__abc_42281_new_n2405_));
AND2X2 AND2X2_6726 ( .A(alu__abc_42281_new_n2406_), .B(alu__abc_42281_new_n1803_), .Y(alu__abc_42281_new_n2407_));
AND2X2 AND2X2_6727 ( .A(alu__abc_42281_new_n2409_), .B(alu__abc_42281_new_n2410_), .Y(alu__abc_42281_new_n2411_));
AND2X2 AND2X2_6728 ( .A(alu__abc_42281_new_n2412_), .B(alu__abc_42281_new_n2413_), .Y(alu__abc_42281_new_n2414_));
AND2X2 AND2X2_6729 ( .A(alu__abc_42281_new_n2415_), .B(alu__abc_42281_new_n2416_), .Y(alu__abc_42281_new_n2417_));
AND2X2 AND2X2_673 ( .A(_abc_44694_new_n1337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n1870_));
AND2X2 AND2X2_6730 ( .A(alu__abc_42281_new_n2417_), .B(alu__abc_42281_new_n936__bF_buf0), .Y(alu__abc_42281_new_n2418_));
AND2X2 AND2X2_6731 ( .A(alu__abc_42281_new_n1779_), .B(alu__abc_42281_new_n1818_), .Y(alu__abc_42281_new_n2419_));
AND2X2 AND2X2_6732 ( .A(alu__abc_42281_new_n950__bF_buf3), .B(alu_a_i_31_), .Y(alu__abc_42281_new_n2420_));
AND2X2 AND2X2_6733 ( .A(alu__abc_42281_new_n512_), .B(alu__abc_42281_new_n941__bF_buf3), .Y(alu__abc_42281_new_n2421_));
AND2X2 AND2X2_6734 ( .A(alu__abc_42281_new_n939__bF_buf3), .B(alu__abc_42281_new_n241_), .Y(alu__abc_42281_new_n2422_));
AND2X2 AND2X2_6735 ( .A(alu__abc_42281_new_n928__bF_buf3), .B(alu__abc_42281_new_n530_), .Y(alu__abc_42281_new_n2423_));
AND2X2 AND2X2_6736 ( .A(alu__abc_42281_new_n2434_), .B(alu__abc_42281_new_n2433_), .Y(alu_greater_than_signed_o));
AND2X2 AND2X2_6737 ( .A(alu__abc_42281_new_n1136_), .B(alu__abc_42281_new_n2436_), .Y(alu__abc_42281_new_n2437_));
AND2X2 AND2X2_6738 ( .A(alu__abc_42281_new_n2438_), .B(alu__abc_42281_new_n302_), .Y(alu__abc_42281_new_n2439_));
AND2X2 AND2X2_6739 ( .A(alu__abc_42281_new_n293_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n2440_));
AND2X2 AND2X2_674 ( .A(_abc_44694_new_n1872_), .B(_abc_44694_new_n1854_), .Y(_abc_44694_new_n1873_));
AND2X2 AND2X2_6740 ( .A(alu__abc_42281_new_n301_), .B(alu__abc_42281_new_n2440_), .Y(alu__abc_42281_new_n2441_));
AND2X2 AND2X2_6741 ( .A(alu__abc_42281_new_n2443_), .B(alu__abc_42281_new_n278_), .Y(alu__abc_42281_new_n2444_));
AND2X2 AND2X2_6742 ( .A(alu__abc_42281_new_n253_), .B(alu_b_i_6_), .Y(alu__abc_42281_new_n2445_));
AND2X2 AND2X2_6743 ( .A(alu__abc_42281_new_n262_), .B(alu__abc_42281_new_n2445_), .Y(alu__abc_42281_new_n2446_));
AND2X2 AND2X2_6744 ( .A(alu__abc_42281_new_n272_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n2448_));
AND2X2 AND2X2_6745 ( .A(alu__abc_42281_new_n268_), .B(alu__abc_42281_new_n2448_), .Y(alu__abc_42281_new_n2449_));
AND2X2 AND2X2_6746 ( .A(alu__abc_42281_new_n2450_), .B(alu__abc_42281_new_n263_), .Y(alu__abc_42281_new_n2451_));
AND2X2 AND2X2_6747 ( .A(alu__abc_42281_new_n2453_), .B(alu__abc_42281_new_n375_), .Y(alu__abc_42281_new_n2454_));
AND2X2 AND2X2_6748 ( .A(alu__abc_42281_new_n351_), .B(alu_b_i_11_), .Y(alu__abc_42281_new_n2455_));
AND2X2 AND2X2_6749 ( .A(alu__abc_42281_new_n343_), .B(alu_b_i_10_), .Y(alu__abc_42281_new_n2456_));
AND2X2 AND2X2_675 ( .A(_abc_44694_new_n1522__bF_buf0), .B(epc_q_14_), .Y(_abc_44694_new_n1875_));
AND2X2 AND2X2_6750 ( .A(alu__abc_42281_new_n355_), .B(alu__abc_42281_new_n2456_), .Y(alu__abc_42281_new_n2457_));
AND2X2 AND2X2_6751 ( .A(alu__abc_42281_new_n360_), .B(alu_b_i_8_), .Y(alu__abc_42281_new_n2459_));
AND2X2 AND2X2_6752 ( .A(alu__abc_42281_new_n2460_), .B(alu__abc_42281_new_n416_), .Y(alu__abc_42281_new_n2461_));
AND2X2 AND2X2_6753 ( .A(alu__abc_42281_new_n356_), .B(alu__abc_42281_new_n2461_), .Y(alu__abc_42281_new_n2462_));
AND2X2 AND2X2_6754 ( .A(alu__abc_42281_new_n2463_), .B(alu__abc_42281_new_n339_), .Y(alu__abc_42281_new_n2464_));
AND2X2 AND2X2_6755 ( .A(alu__abc_42281_new_n333_), .B(alu_b_i_15_), .Y(alu__abc_42281_new_n2465_));
AND2X2 AND2X2_6756 ( .A(alu__abc_42281_new_n325_), .B(alu_b_i_14_), .Y(alu__abc_42281_new_n2466_));
AND2X2 AND2X2_6757 ( .A(alu__abc_42281_new_n337_), .B(alu__abc_42281_new_n2466_), .Y(alu__abc_42281_new_n2467_));
AND2X2 AND2X2_6758 ( .A(alu__abc_42281_new_n308_), .B(alu_b_i_12_), .Y(alu__abc_42281_new_n2469_));
AND2X2 AND2X2_6759 ( .A(alu__abc_42281_new_n2470_), .B(alu__abc_42281_new_n431_), .Y(alu__abc_42281_new_n2471_));
AND2X2 AND2X2_676 ( .A(_abc_44694_new_n1348__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_14_), .Y(_abc_44694_new_n1876_));
AND2X2 AND2X2_6760 ( .A(alu__abc_42281_new_n338_), .B(alu__abc_42281_new_n2471_), .Y(alu__abc_42281_new_n2472_));
AND2X2 AND2X2_6761 ( .A(alu__abc_42281_new_n2475_), .B(alu__abc_42281_new_n249_), .Y(alu__abc_42281_new_n2476_));
AND2X2 AND2X2_6762 ( .A(alu__abc_42281_new_n209_), .B(alu_b_i_27_), .Y(alu__abc_42281_new_n2477_));
AND2X2 AND2X2_6763 ( .A(alu__abc_42281_new_n201_), .B(alu_b_i_26_), .Y(alu__abc_42281_new_n2478_));
AND2X2 AND2X2_6764 ( .A(alu__abc_42281_new_n213_), .B(alu__abc_42281_new_n2478_), .Y(alu__abc_42281_new_n2479_));
AND2X2 AND2X2_6765 ( .A(alu__abc_42281_new_n192_), .B(alu_b_i_24_), .Y(alu__abc_42281_new_n2481_));
AND2X2 AND2X2_6766 ( .A(alu__abc_42281_new_n2482_), .B(alu__abc_42281_new_n487_), .Y(alu__abc_42281_new_n2483_));
AND2X2 AND2X2_6767 ( .A(alu__abc_42281_new_n214_), .B(alu__abc_42281_new_n2483_), .Y(alu__abc_42281_new_n2484_));
AND2X2 AND2X2_6768 ( .A(alu__abc_42281_new_n2485_), .B(alu__abc_42281_new_n247_), .Y(alu__abc_42281_new_n2486_));
AND2X2 AND2X2_6769 ( .A(alu__abc_42281_new_n243_), .B(alu_b_i_31_), .Y(alu__abc_42281_new_n2487_));
AND2X2 AND2X2_677 ( .A(_abc_44694_new_n1207__bF_buf5), .B(_abc_44694_new_n1878_), .Y(_abc_44694_new_n1879_));
AND2X2 AND2X2_6770 ( .A(alu__abc_42281_new_n236_), .B(alu_b_i_30_), .Y(alu__abc_42281_new_n2488_));
AND2X2 AND2X2_6771 ( .A(alu__abc_42281_new_n245_), .B(alu__abc_42281_new_n2488_), .Y(alu__abc_42281_new_n2489_));
AND2X2 AND2X2_6772 ( .A(alu__abc_42281_new_n219_), .B(alu_b_i_28_), .Y(alu__abc_42281_new_n2491_));
AND2X2 AND2X2_6773 ( .A(alu__abc_42281_new_n2492_), .B(alu__abc_42281_new_n499_), .Y(alu__abc_42281_new_n2493_));
AND2X2 AND2X2_6774 ( .A(alu__abc_42281_new_n246_), .B(alu__abc_42281_new_n2493_), .Y(alu__abc_42281_new_n2494_));
AND2X2 AND2X2_6775 ( .A(alu__abc_42281_new_n156_), .B(alu_b_i_19_), .Y(alu__abc_42281_new_n2497_));
AND2X2 AND2X2_6776 ( .A(alu__abc_42281_new_n148_), .B(alu_b_i_18_), .Y(alu__abc_42281_new_n2498_));
AND2X2 AND2X2_6777 ( .A(alu__abc_42281_new_n160_), .B(alu__abc_42281_new_n2498_), .Y(alu__abc_42281_new_n2499_));
AND2X2 AND2X2_6778 ( .A(alu__abc_42281_new_n165_), .B(alu_b_i_16_), .Y(alu__abc_42281_new_n2501_));
AND2X2 AND2X2_6779 ( .A(alu__abc_42281_new_n2502_), .B(alu__abc_42281_new_n448_), .Y(alu__abc_42281_new_n2503_));
AND2X2 AND2X2_678 ( .A(_abc_44694_new_n1874_), .B(_abc_44694_new_n1879_), .Y(_abc_44694_new_n1880_));
AND2X2 AND2X2_6780 ( .A(alu__abc_42281_new_n161_), .B(alu__abc_42281_new_n2503_), .Y(alu__abc_42281_new_n2504_));
AND2X2 AND2X2_6781 ( .A(alu__abc_42281_new_n2505_), .B(alu__abc_42281_new_n144_), .Y(alu__abc_42281_new_n2506_));
AND2X2 AND2X2_6782 ( .A(alu__abc_42281_new_n138_), .B(alu_b_i_23_), .Y(alu__abc_42281_new_n2507_));
AND2X2 AND2X2_6783 ( .A(alu__abc_42281_new_n130_), .B(alu_b_i_22_), .Y(alu__abc_42281_new_n2508_));
AND2X2 AND2X2_6784 ( .A(alu__abc_42281_new_n142_), .B(alu__abc_42281_new_n2508_), .Y(alu__abc_42281_new_n2509_));
AND2X2 AND2X2_6785 ( .A(alu__abc_42281_new_n113_), .B(alu_b_i_20_), .Y(alu__abc_42281_new_n2511_));
AND2X2 AND2X2_6786 ( .A(alu__abc_42281_new_n2512_), .B(alu__abc_42281_new_n463_), .Y(alu__abc_42281_new_n2513_));
AND2X2 AND2X2_6787 ( .A(alu__abc_42281_new_n143_), .B(alu__abc_42281_new_n2513_), .Y(alu__abc_42281_new_n2514_));
AND2X2 AND2X2_6788 ( .A(alu__abc_42281_new_n2516_), .B(alu__abc_42281_new_n248_), .Y(alu__abc_42281_new_n2517_));
AND2X2 AND2X2_6789 ( .A(alu__abc_42281_new_n2519_), .B(alu__abc_42281_new_n2433_), .Y(alu_less_than_o));
AND2X2 AND2X2_679 ( .A(_abc_44694_new_n1882_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n1883_));
AND2X2 AND2X2_68 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[19] ), .Y(_abc_44694_new_n733_));
AND2X2 AND2X2_680 ( .A(_abc_44694_new_n1881_), .B(_abc_44694_new_n1883_), .Y(_0epc_q_31_0__14_));
AND2X2 AND2X2_681 ( .A(_abc_44694_new_n1849_), .B(pc_q_15_), .Y(_abc_44694_new_n1886_));
AND2X2 AND2X2_682 ( .A(_abc_44694_new_n1887_), .B(_abc_44694_new_n1885_), .Y(_abc_44694_new_n1888_));
AND2X2 AND2X2_683 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1889_), .Y(_abc_44694_new_n1890_));
AND2X2 AND2X2_684 ( .A(_abc_44694_new_n1019__bF_buf1), .B(epc_q_15_), .Y(_abc_44694_new_n1892_));
AND2X2 AND2X2_685 ( .A(_abc_44694_new_n1864_), .B(_abc_44694_new_n1861_), .Y(_abc_44694_new_n1893_));
AND2X2 AND2X2_686 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_44694_new_n1896_));
AND2X2 AND2X2_687 ( .A(_abc_44694_new_n1897_), .B(_abc_44694_new_n1895_), .Y(_abc_44694_new_n1898_));
AND2X2 AND2X2_688 ( .A(_abc_44694_new_n1901_), .B(_abc_44694_new_n1194__bF_buf4), .Y(_abc_44694_new_n1902_));
AND2X2 AND2X2_689 ( .A(_abc_44694_new_n1902_), .B(_abc_44694_new_n1899_), .Y(_abc_44694_new_n1903_));
AND2X2 AND2X2_69 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[19] ), .Y(_abc_44694_new_n736_));
AND2X2 AND2X2_690 ( .A(_abc_44694_new_n1904_), .B(_abc_44694_new_n1340__bF_buf4), .Y(_abc_44694_new_n1905_));
AND2X2 AND2X2_691 ( .A(_abc_44694_new_n1337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n1906_));
AND2X2 AND2X2_692 ( .A(_abc_44694_new_n1908_), .B(_abc_44694_new_n1891_), .Y(_abc_44694_new_n1909_));
AND2X2 AND2X2_693 ( .A(_abc_44694_new_n1522__bF_buf4), .B(epc_q_15_), .Y(_abc_44694_new_n1911_));
AND2X2 AND2X2_694 ( .A(_abc_44694_new_n1348__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n1912_));
AND2X2 AND2X2_695 ( .A(_abc_44694_new_n1207__bF_buf4), .B(_abc_44694_new_n1914_), .Y(_abc_44694_new_n1915_));
AND2X2 AND2X2_696 ( .A(_abc_44694_new_n1910_), .B(_abc_44694_new_n1915_), .Y(_abc_44694_new_n1916_));
AND2X2 AND2X2_697 ( .A(_abc_44694_new_n1918_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n1919_));
AND2X2 AND2X2_698 ( .A(_abc_44694_new_n1917_), .B(_abc_44694_new_n1919_), .Y(_0epc_q_31_0__15_));
AND2X2 AND2X2_699 ( .A(_abc_44694_new_n1886_), .B(pc_q_16_), .Y(_abc_44694_new_n1922_));
AND2X2 AND2X2_7 ( .A(_abc_44694_new_n628_), .B(_abc_44694_new_n622_), .Y(inst_trap_w));
AND2X2 AND2X2_70 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[11] ), .Y(_abc_44694_new_n737_));
AND2X2 AND2X2_700 ( .A(_abc_44694_new_n1923_), .B(_abc_44694_new_n1921_), .Y(_abc_44694_new_n1924_));
AND2X2 AND2X2_701 ( .A(_abc_44694_new_n1535_), .B(_abc_44694_new_n1925_), .Y(_abc_44694_new_n1926_));
AND2X2 AND2X2_702 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_16_), .Y(_abc_44694_new_n1928_));
AND2X2 AND2X2_703 ( .A(_abc_44694_new_n1862_), .B(_abc_44694_new_n1898_), .Y(_abc_44694_new_n1929_));
AND2X2 AND2X2_704 ( .A(_abc_44694_new_n1823_), .B(_abc_44694_new_n1929_), .Y(_abc_44694_new_n1930_));
AND2X2 AND2X2_705 ( .A(_abc_44694_new_n1779_), .B(_abc_44694_new_n1930_), .Y(_abc_44694_new_n1931_));
AND2X2 AND2X2_706 ( .A(_abc_44694_new_n1895_), .B(_abc_44694_new_n1860_), .Y(_abc_44694_new_n1932_));
AND2X2 AND2X2_707 ( .A(_abc_44694_new_n1934_), .B(_abc_44694_new_n1929_), .Y(_abc_44694_new_n1935_));
AND2X2 AND2X2_708 ( .A(_abc_44694_new_n1780_), .B(_abc_44694_new_n1930_), .Y(_abc_44694_new_n1938_));
AND2X2 AND2X2_709 ( .A(_abc_44694_new_n1624_), .B(_abc_44694_new_n1938_), .Y(_abc_44694_new_n1939_));
AND2X2 AND2X2_71 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[27] ), .Y(_abc_44694_new_n739_));
AND2X2 AND2X2_710 ( .A(pc_q_16_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_44694_new_n1942_));
AND2X2 AND2X2_711 ( .A(_abc_44694_new_n1943_), .B(_abc_44694_new_n1941_), .Y(_abc_44694_new_n1944_));
AND2X2 AND2X2_712 ( .A(_abc_44694_new_n1940_), .B(_abc_44694_new_n1944_), .Y(_abc_44694_new_n1946_));
AND2X2 AND2X2_713 ( .A(_abc_44694_new_n1947_), .B(_abc_44694_new_n1194__bF_buf3), .Y(_abc_44694_new_n1948_));
AND2X2 AND2X2_714 ( .A(_abc_44694_new_n1948_), .B(_abc_44694_new_n1945_), .Y(_abc_44694_new_n1949_));
AND2X2 AND2X2_715 ( .A(_abc_44694_new_n1950_), .B(_abc_44694_new_n1340__bF_buf3), .Y(_abc_44694_new_n1951_));
AND2X2 AND2X2_716 ( .A(_abc_44694_new_n1337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_44694_new_n1952_));
AND2X2 AND2X2_717 ( .A(_abc_44694_new_n1954_), .B(_abc_44694_new_n1927_), .Y(_abc_44694_new_n1955_));
AND2X2 AND2X2_718 ( .A(_abc_44694_new_n1522__bF_buf3), .B(epc_q_16_), .Y(_abc_44694_new_n1957_));
AND2X2 AND2X2_719 ( .A(_abc_44694_new_n1348__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_44694_new_n1958_));
AND2X2 AND2X2_72 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[3] ), .Y(_abc_44694_new_n740_));
AND2X2 AND2X2_720 ( .A(_abc_44694_new_n1207__bF_buf3), .B(_abc_44694_new_n1960_), .Y(_abc_44694_new_n1961_));
AND2X2 AND2X2_721 ( .A(_abc_44694_new_n1956_), .B(_abc_44694_new_n1961_), .Y(_abc_44694_new_n1962_));
AND2X2 AND2X2_722 ( .A(_abc_44694_new_n1964_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n1965_));
AND2X2 AND2X2_723 ( .A(_abc_44694_new_n1963_), .B(_abc_44694_new_n1965_), .Y(_0epc_q_31_0__16_));
AND2X2 AND2X2_724 ( .A(_abc_44694_new_n1922_), .B(pc_q_17_), .Y(_abc_44694_new_n1968_));
AND2X2 AND2X2_725 ( .A(_abc_44694_new_n1969_), .B(_abc_44694_new_n1967_), .Y(_abc_44694_new_n1970_));
AND2X2 AND2X2_726 ( .A(_abc_44694_new_n1971_), .B(_abc_44694_new_n1535_), .Y(_abc_44694_new_n1972_));
AND2X2 AND2X2_727 ( .A(_abc_44694_new_n1019__bF_buf4), .B(epc_q_17_), .Y(_abc_44694_new_n1974_));
AND2X2 AND2X2_728 ( .A(pc_q_17_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf4_), .Y(_abc_44694_new_n1976_));
AND2X2 AND2X2_729 ( .A(_abc_44694_new_n1977_), .B(_abc_44694_new_n1975_), .Y(_abc_44694_new_n1978_));
AND2X2 AND2X2_73 ( .A(_abc_44694_new_n743_), .B(state_q_1_bF_buf3_), .Y(_abc_44694_new_n744_));
AND2X2 AND2X2_730 ( .A(_abc_44694_new_n1947_), .B(_abc_44694_new_n1943_), .Y(_abc_44694_new_n1979_));
AND2X2 AND2X2_731 ( .A(_abc_44694_new_n1980_), .B(_abc_44694_new_n1978_), .Y(_abc_44694_new_n1981_));
AND2X2 AND2X2_732 ( .A(_abc_44694_new_n1983_), .B(_abc_44694_new_n1194__bF_buf2), .Y(_abc_44694_new_n1984_));
AND2X2 AND2X2_733 ( .A(_abc_44694_new_n1984_), .B(_abc_44694_new_n1982_), .Y(_abc_44694_new_n1985_));
AND2X2 AND2X2_734 ( .A(_abc_44694_new_n1986_), .B(_abc_44694_new_n1340__bF_buf2), .Y(_abc_44694_new_n1987_));
AND2X2 AND2X2_735 ( .A(_abc_44694_new_n1337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_44694_new_n1988_));
AND2X2 AND2X2_736 ( .A(_abc_44694_new_n1990_), .B(_abc_44694_new_n1973_), .Y(_abc_44694_new_n1991_));
AND2X2 AND2X2_737 ( .A(_abc_44694_new_n1522__bF_buf2), .B(epc_q_17_), .Y(_abc_44694_new_n1993_));
AND2X2 AND2X2_738 ( .A(_abc_44694_new_n1348__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_44694_new_n1994_));
AND2X2 AND2X2_739 ( .A(_abc_44694_new_n1207__bF_buf2), .B(_abc_44694_new_n1996_), .Y(_abc_44694_new_n1997_));
AND2X2 AND2X2_74 ( .A(_abc_44694_new_n735_), .B(_abc_44694_new_n744_), .Y(_abc_44694_new_n745_));
AND2X2 AND2X2_740 ( .A(_abc_44694_new_n1992_), .B(_abc_44694_new_n1997_), .Y(_abc_44694_new_n1998_));
AND2X2 AND2X2_741 ( .A(_abc_44694_new_n2000_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n2001_));
AND2X2 AND2X2_742 ( .A(_abc_44694_new_n1999_), .B(_abc_44694_new_n2001_), .Y(_0epc_q_31_0__17_));
AND2X2 AND2X2_743 ( .A(_abc_44694_new_n1968_), .B(pc_q_18_), .Y(_abc_44694_new_n2004_));
AND2X2 AND2X2_744 ( .A(_abc_44694_new_n2005_), .B(_abc_44694_new_n2003_), .Y(_abc_44694_new_n2006_));
AND2X2 AND2X2_745 ( .A(_abc_44694_new_n2006_), .B(_abc_44694_new_n1382__bF_buf3), .Y(_abc_44694_new_n2007_));
AND2X2 AND2X2_746 ( .A(_abc_44694_new_n1019__bF_buf3), .B(epc_q_18_), .Y(_abc_44694_new_n2010_));
AND2X2 AND2X2_747 ( .A(_abc_44694_new_n1982_), .B(_abc_44694_new_n1977_), .Y(_abc_44694_new_n2011_));
AND2X2 AND2X2_748 ( .A(pc_q_18_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_44694_new_n2014_));
AND2X2 AND2X2_749 ( .A(_abc_44694_new_n2015_), .B(_abc_44694_new_n2013_), .Y(_abc_44694_new_n2016_));
AND2X2 AND2X2_75 ( .A(_abc_44694_new_n671_), .B(alu_p_o_4_), .Y(_abc_44694_new_n747_));
AND2X2 AND2X2_750 ( .A(_abc_44694_new_n2012_), .B(_abc_44694_new_n2016_), .Y(_abc_44694_new_n2017_));
AND2X2 AND2X2_751 ( .A(_abc_44694_new_n2019_), .B(_abc_44694_new_n1194__bF_buf1), .Y(_abc_44694_new_n2020_));
AND2X2 AND2X2_752 ( .A(_abc_44694_new_n2020_), .B(_abc_44694_new_n2018_), .Y(_abc_44694_new_n2021_));
AND2X2 AND2X2_753 ( .A(_abc_44694_new_n2022_), .B(_abc_44694_new_n1340__bF_buf1), .Y(_abc_44694_new_n2023_));
AND2X2 AND2X2_754 ( .A(_abc_44694_new_n1337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_44694_new_n2024_));
AND2X2 AND2X2_755 ( .A(_abc_44694_new_n2026_), .B(_abc_44694_new_n2009_), .Y(_abc_44694_new_n2027_));
AND2X2 AND2X2_756 ( .A(_abc_44694_new_n1522__bF_buf1), .B(epc_q_18_), .Y(_abc_44694_new_n2029_));
AND2X2 AND2X2_757 ( .A(_abc_44694_new_n1348__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_44694_new_n2030_));
AND2X2 AND2X2_758 ( .A(_abc_44694_new_n1207__bF_buf1), .B(_abc_44694_new_n2032_), .Y(_abc_44694_new_n2033_));
AND2X2 AND2X2_759 ( .A(_abc_44694_new_n2028_), .B(_abc_44694_new_n2033_), .Y(_abc_44694_new_n2034_));
AND2X2 AND2X2_76 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[4] ), .Y(_abc_44694_new_n748_));
AND2X2 AND2X2_760 ( .A(_abc_44694_new_n2036_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n2037_));
AND2X2 AND2X2_761 ( .A(_abc_44694_new_n2035_), .B(_abc_44694_new_n2037_), .Y(_0epc_q_31_0__18_));
AND2X2 AND2X2_762 ( .A(_abc_44694_new_n2004_), .B(pc_q_19_), .Y(_abc_44694_new_n2040_));
AND2X2 AND2X2_763 ( .A(_abc_44694_new_n2041_), .B(_abc_44694_new_n2039_), .Y(_abc_44694_new_n2042_));
AND2X2 AND2X2_764 ( .A(_abc_44694_new_n2042_), .B(_abc_44694_new_n1382__bF_buf2), .Y(_abc_44694_new_n2043_));
AND2X2 AND2X2_765 ( .A(_abc_44694_new_n1019__bF_buf2), .B(epc_q_19_), .Y(_abc_44694_new_n2046_));
AND2X2 AND2X2_766 ( .A(_abc_44694_new_n2018_), .B(_abc_44694_new_n2015_), .Y(_abc_44694_new_n2047_));
AND2X2 AND2X2_767 ( .A(pc_q_19_), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_44694_new_n2049_));
AND2X2 AND2X2_768 ( .A(_abc_44694_new_n2050_), .B(_abc_44694_new_n2048_), .Y(_abc_44694_new_n2051_));
AND2X2 AND2X2_769 ( .A(_abc_44694_new_n2055_), .B(_abc_44694_new_n1194__bF_buf0), .Y(_abc_44694_new_n2056_));
AND2X2 AND2X2_77 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[20] ), .Y(_abc_44694_new_n749_));
AND2X2 AND2X2_770 ( .A(_abc_44694_new_n2056_), .B(_abc_44694_new_n2053_), .Y(_abc_44694_new_n2057_));
AND2X2 AND2X2_771 ( .A(_abc_44694_new_n2058_), .B(_abc_44694_new_n1340__bF_buf0), .Y(_abc_44694_new_n2059_));
AND2X2 AND2X2_772 ( .A(_abc_44694_new_n1337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_44694_new_n2060_));
AND2X2 AND2X2_773 ( .A(_abc_44694_new_n2062_), .B(_abc_44694_new_n2045_), .Y(_abc_44694_new_n2063_));
AND2X2 AND2X2_774 ( .A(_abc_44694_new_n1522__bF_buf0), .B(epc_q_19_), .Y(_abc_44694_new_n2065_));
AND2X2 AND2X2_775 ( .A(_abc_44694_new_n1348__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_44694_new_n2066_));
AND2X2 AND2X2_776 ( .A(_abc_44694_new_n1207__bF_buf0), .B(_abc_44694_new_n2068_), .Y(_abc_44694_new_n2069_));
AND2X2 AND2X2_777 ( .A(_abc_44694_new_n2064_), .B(_abc_44694_new_n2069_), .Y(_abc_44694_new_n2070_));
AND2X2 AND2X2_778 ( .A(_abc_44694_new_n2072_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n2073_));
AND2X2 AND2X2_779 ( .A(_abc_44694_new_n2071_), .B(_abc_44694_new_n2073_), .Y(_0epc_q_31_0__19_));
AND2X2 AND2X2_78 ( .A(_abc_44694_new_n750_), .B(_abc_44694_new_n673__bF_buf0), .Y(_abc_44694_new_n751_));
AND2X2 AND2X2_780 ( .A(_abc_44694_new_n2040_), .B(pc_q_20_), .Y(_abc_44694_new_n2076_));
AND2X2 AND2X2_781 ( .A(_abc_44694_new_n2077_), .B(_abc_44694_new_n2075_), .Y(_abc_44694_new_n2078_));
AND2X2 AND2X2_782 ( .A(_abc_44694_new_n2078_), .B(_abc_44694_new_n1382__bF_buf1), .Y(_abc_44694_new_n2079_));
AND2X2 AND2X2_783 ( .A(_abc_44694_new_n1019__bF_buf1), .B(epc_q_20_), .Y(_abc_44694_new_n2082_));
AND2X2 AND2X2_784 ( .A(_abc_44694_new_n1975_), .B(_abc_44694_new_n1942_), .Y(_abc_44694_new_n2083_));
AND2X2 AND2X2_785 ( .A(_abc_44694_new_n2016_), .B(_abc_44694_new_n2051_), .Y(_abc_44694_new_n2085_));
AND2X2 AND2X2_786 ( .A(_abc_44694_new_n2085_), .B(_abc_44694_new_n2084_), .Y(_abc_44694_new_n2086_));
AND2X2 AND2X2_787 ( .A(_abc_44694_new_n2048_), .B(_abc_44694_new_n2014_), .Y(_abc_44694_new_n2087_));
AND2X2 AND2X2_788 ( .A(_abc_44694_new_n1944_), .B(_abc_44694_new_n1978_), .Y(_abc_44694_new_n2092_));
AND2X2 AND2X2_789 ( .A(_abc_44694_new_n2092_), .B(_abc_44694_new_n2085_), .Y(_abc_44694_new_n2093_));
AND2X2 AND2X2_79 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[28] ), .Y(_abc_44694_new_n752_));
AND2X2 AND2X2_790 ( .A(_abc_44694_new_n2095_), .B(_abc_44694_new_n2090_), .Y(_abc_44694_new_n2096_));
AND2X2 AND2X2_791 ( .A(pc_q_20_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_44694_new_n2099_));
AND2X2 AND2X2_792 ( .A(_abc_44694_new_n2100_), .B(_abc_44694_new_n2098_), .Y(_abc_44694_new_n2101_));
AND2X2 AND2X2_793 ( .A(_abc_44694_new_n2097_), .B(_abc_44694_new_n2101_), .Y(_abc_44694_new_n2102_));
AND2X2 AND2X2_794 ( .A(_abc_44694_new_n2104_), .B(_abc_44694_new_n1194__bF_buf4), .Y(_abc_44694_new_n2105_));
AND2X2 AND2X2_795 ( .A(_abc_44694_new_n2105_), .B(_abc_44694_new_n2103_), .Y(_abc_44694_new_n2106_));
AND2X2 AND2X2_796 ( .A(_abc_44694_new_n2107_), .B(_abc_44694_new_n1340__bF_buf4), .Y(_abc_44694_new_n2108_));
AND2X2 AND2X2_797 ( .A(_abc_44694_new_n1337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_44694_new_n2109_));
AND2X2 AND2X2_798 ( .A(_abc_44694_new_n2111_), .B(_abc_44694_new_n2081_), .Y(_abc_44694_new_n2112_));
AND2X2 AND2X2_799 ( .A(_abc_44694_new_n1522__bF_buf4), .B(epc_q_20_), .Y(_abc_44694_new_n2114_));
AND2X2 AND2X2_8 ( .A(_abc_44694_new_n631_), .B(inst_r_2_), .Y(_abc_44694_new_n632_));
AND2X2 AND2X2_80 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[12] ), .Y(_abc_44694_new_n753_));
AND2X2 AND2X2_800 ( .A(_abc_44694_new_n1348__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_44694_new_n2115_));
AND2X2 AND2X2_801 ( .A(_abc_44694_new_n1207__bF_buf5), .B(_abc_44694_new_n2117_), .Y(_abc_44694_new_n2118_));
AND2X2 AND2X2_802 ( .A(_abc_44694_new_n2113_), .B(_abc_44694_new_n2118_), .Y(_abc_44694_new_n2119_));
AND2X2 AND2X2_803 ( .A(_abc_44694_new_n2121_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n2122_));
AND2X2 AND2X2_804 ( .A(_abc_44694_new_n2120_), .B(_abc_44694_new_n2122_), .Y(_0epc_q_31_0__20_));
AND2X2 AND2X2_805 ( .A(_abc_44694_new_n2076_), .B(pc_q_21_), .Y(_abc_44694_new_n2125_));
AND2X2 AND2X2_806 ( .A(_abc_44694_new_n2126_), .B(_abc_44694_new_n2124_), .Y(_abc_44694_new_n2127_));
AND2X2 AND2X2_807 ( .A(_abc_44694_new_n2127_), .B(_abc_44694_new_n1382__bF_buf0), .Y(_abc_44694_new_n2128_));
AND2X2 AND2X2_808 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_21_), .Y(_abc_44694_new_n2131_));
AND2X2 AND2X2_809 ( .A(pc_q_21_), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_44694_new_n2133_));
AND2X2 AND2X2_81 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[20] ), .Y(_abc_44694_new_n755_));
AND2X2 AND2X2_810 ( .A(_abc_44694_new_n2134_), .B(_abc_44694_new_n2132_), .Y(_abc_44694_new_n2135_));
AND2X2 AND2X2_811 ( .A(_abc_44694_new_n2101_), .B(_abc_44694_new_n2135_), .Y(_abc_44694_new_n2138_));
AND2X2 AND2X2_812 ( .A(_abc_44694_new_n2097_), .B(_abc_44694_new_n2138_), .Y(_abc_44694_new_n2139_));
AND2X2 AND2X2_813 ( .A(_abc_44694_new_n2135_), .B(_abc_44694_new_n2099_), .Y(_abc_44694_new_n2141_));
AND2X2 AND2X2_814 ( .A(_abc_44694_new_n1194__bF_buf3), .B(_abc_44694_new_n2142_), .Y(_abc_44694_new_n2143_));
AND2X2 AND2X2_815 ( .A(_abc_44694_new_n2140_), .B(_abc_44694_new_n2143_), .Y(_abc_44694_new_n2144_));
AND2X2 AND2X2_816 ( .A(_abc_44694_new_n2144_), .B(_abc_44694_new_n2137_), .Y(_abc_44694_new_n2145_));
AND2X2 AND2X2_817 ( .A(_abc_44694_new_n2146_), .B(_abc_44694_new_n1340__bF_buf3), .Y(_abc_44694_new_n2147_));
AND2X2 AND2X2_818 ( .A(_abc_44694_new_n1337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_44694_new_n2148_));
AND2X2 AND2X2_819 ( .A(_abc_44694_new_n2150_), .B(_abc_44694_new_n2130_), .Y(_abc_44694_new_n2151_));
AND2X2 AND2X2_82 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[4] ), .Y(_abc_44694_new_n756_));
AND2X2 AND2X2_820 ( .A(_abc_44694_new_n1522__bF_buf3), .B(epc_q_21_), .Y(_abc_44694_new_n2153_));
AND2X2 AND2X2_821 ( .A(_abc_44694_new_n1348__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_44694_new_n2154_));
AND2X2 AND2X2_822 ( .A(_abc_44694_new_n1207__bF_buf4), .B(_abc_44694_new_n2156_), .Y(_abc_44694_new_n2157_));
AND2X2 AND2X2_823 ( .A(_abc_44694_new_n2152_), .B(_abc_44694_new_n2157_), .Y(_abc_44694_new_n2158_));
AND2X2 AND2X2_824 ( .A(_abc_44694_new_n2160_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n2161_));
AND2X2 AND2X2_825 ( .A(_abc_44694_new_n2159_), .B(_abc_44694_new_n2161_), .Y(_0epc_q_31_0__21_));
AND2X2 AND2X2_826 ( .A(_abc_44694_new_n2125_), .B(pc_q_22_), .Y(_abc_44694_new_n2164_));
AND2X2 AND2X2_827 ( .A(_abc_44694_new_n2165_), .B(_abc_44694_new_n2163_), .Y(_abc_44694_new_n2166_));
AND2X2 AND2X2_828 ( .A(_abc_44694_new_n2166_), .B(_abc_44694_new_n1382__bF_buf3), .Y(_abc_44694_new_n2167_));
AND2X2 AND2X2_829 ( .A(_abc_44694_new_n1019__bF_buf4), .B(epc_q_22_), .Y(_abc_44694_new_n2170_));
AND2X2 AND2X2_83 ( .A(_abc_44694_new_n758_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n759_));
AND2X2 AND2X2_830 ( .A(_abc_44694_new_n2142_), .B(_abc_44694_new_n2134_), .Y(_abc_44694_new_n2171_));
AND2X2 AND2X2_831 ( .A(_abc_44694_new_n2140_), .B(_abc_44694_new_n2171_), .Y(_abc_44694_new_n2172_));
AND2X2 AND2X2_832 ( .A(pc_q_22_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf2_), .Y(_abc_44694_new_n2175_));
AND2X2 AND2X2_833 ( .A(_abc_44694_new_n2176_), .B(_abc_44694_new_n2174_), .Y(_abc_44694_new_n2177_));
AND2X2 AND2X2_834 ( .A(_abc_44694_new_n2173_), .B(_abc_44694_new_n2177_), .Y(_abc_44694_new_n2178_));
AND2X2 AND2X2_835 ( .A(_abc_44694_new_n2180_), .B(_abc_44694_new_n1194__bF_buf2), .Y(_abc_44694_new_n2181_));
AND2X2 AND2X2_836 ( .A(_abc_44694_new_n2181_), .B(_abc_44694_new_n2179_), .Y(_abc_44694_new_n2182_));
AND2X2 AND2X2_837 ( .A(_abc_44694_new_n2183_), .B(_abc_44694_new_n1340__bF_buf2), .Y(_abc_44694_new_n2184_));
AND2X2 AND2X2_838 ( .A(_abc_44694_new_n1337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_44694_new_n2185_));
AND2X2 AND2X2_839 ( .A(_abc_44694_new_n2187_), .B(_abc_44694_new_n2169_), .Y(_abc_44694_new_n2188_));
AND2X2 AND2X2_84 ( .A(_abc_44694_new_n760_), .B(state_q_1_bF_buf2_), .Y(_abc_44694_new_n761_));
AND2X2 AND2X2_840 ( .A(_abc_44694_new_n1522__bF_buf2), .B(epc_q_22_), .Y(_abc_44694_new_n2190_));
AND2X2 AND2X2_841 ( .A(_abc_44694_new_n1348__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_44694_new_n2191_));
AND2X2 AND2X2_842 ( .A(_abc_44694_new_n1207__bF_buf3), .B(_abc_44694_new_n2193_), .Y(_abc_44694_new_n2194_));
AND2X2 AND2X2_843 ( .A(_abc_44694_new_n2189_), .B(_abc_44694_new_n2194_), .Y(_abc_44694_new_n2195_));
AND2X2 AND2X2_844 ( .A(_abc_44694_new_n2197_), .B(enable_i_bF_buf1), .Y(_abc_44694_new_n2198_));
AND2X2 AND2X2_845 ( .A(_abc_44694_new_n2196_), .B(_abc_44694_new_n2198_), .Y(_0epc_q_31_0__22_));
AND2X2 AND2X2_846 ( .A(_abc_44694_new_n2164_), .B(pc_q_23_), .Y(_abc_44694_new_n2201_));
AND2X2 AND2X2_847 ( .A(_abc_44694_new_n2202_), .B(_abc_44694_new_n2200_), .Y(_abc_44694_new_n2203_));
AND2X2 AND2X2_848 ( .A(_abc_44694_new_n2203_), .B(_abc_44694_new_n1382__bF_buf2), .Y(_abc_44694_new_n2204_));
AND2X2 AND2X2_849 ( .A(_abc_44694_new_n1019__bF_buf3), .B(epc_q_23_), .Y(_abc_44694_new_n2207_));
AND2X2 AND2X2_85 ( .A(_abc_44694_new_n671_), .B(alu_p_o_5_), .Y(_abc_44694_new_n763_));
AND2X2 AND2X2_850 ( .A(_abc_44694_new_n2179_), .B(_abc_44694_new_n2176_), .Y(_abc_44694_new_n2208_));
AND2X2 AND2X2_851 ( .A(opcode_q_21_), .B(pc_q_23_), .Y(_abc_44694_new_n2211_));
AND2X2 AND2X2_852 ( .A(_abc_44694_new_n2212_), .B(_abc_44694_new_n2210_), .Y(_abc_44694_new_n2213_));
AND2X2 AND2X2_853 ( .A(_abc_44694_new_n2216_), .B(_abc_44694_new_n1194__bF_buf1), .Y(_abc_44694_new_n2217_));
AND2X2 AND2X2_854 ( .A(_abc_44694_new_n2217_), .B(_abc_44694_new_n2214_), .Y(_abc_44694_new_n2218_));
AND2X2 AND2X2_855 ( .A(_abc_44694_new_n2219_), .B(_abc_44694_new_n1340__bF_buf1), .Y(_abc_44694_new_n2220_));
AND2X2 AND2X2_856 ( .A(_abc_44694_new_n1337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_44694_new_n2221_));
AND2X2 AND2X2_857 ( .A(_abc_44694_new_n2223_), .B(_abc_44694_new_n2206_), .Y(_abc_44694_new_n2224_));
AND2X2 AND2X2_858 ( .A(_abc_44694_new_n1522__bF_buf1), .B(epc_q_23_), .Y(_abc_44694_new_n2226_));
AND2X2 AND2X2_859 ( .A(_abc_44694_new_n1348__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_44694_new_n2227_));
AND2X2 AND2X2_86 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[5] ), .Y(_abc_44694_new_n764_));
AND2X2 AND2X2_860 ( .A(_abc_44694_new_n1207__bF_buf2), .B(_abc_44694_new_n2229_), .Y(_abc_44694_new_n2230_));
AND2X2 AND2X2_861 ( .A(_abc_44694_new_n2225_), .B(_abc_44694_new_n2230_), .Y(_abc_44694_new_n2231_));
AND2X2 AND2X2_862 ( .A(_abc_44694_new_n2233_), .B(enable_i_bF_buf0), .Y(_abc_44694_new_n2234_));
AND2X2 AND2X2_863 ( .A(_abc_44694_new_n2232_), .B(_abc_44694_new_n2234_), .Y(_0epc_q_31_0__23_));
AND2X2 AND2X2_864 ( .A(_abc_44694_new_n2201_), .B(pc_q_24_), .Y(_abc_44694_new_n2237_));
AND2X2 AND2X2_865 ( .A(_abc_44694_new_n2238_), .B(_abc_44694_new_n2236_), .Y(_abc_44694_new_n2239_));
AND2X2 AND2X2_866 ( .A(_abc_44694_new_n2239_), .B(_abc_44694_new_n1382__bF_buf1), .Y(_abc_44694_new_n2240_));
AND2X2 AND2X2_867 ( .A(_abc_44694_new_n2177_), .B(_abc_44694_new_n2213_), .Y(_abc_44694_new_n2242_));
AND2X2 AND2X2_868 ( .A(_abc_44694_new_n2138_), .B(_abc_44694_new_n2242_), .Y(_abc_44694_new_n2243_));
AND2X2 AND2X2_869 ( .A(_abc_44694_new_n2093_), .B(_abc_44694_new_n2243_), .Y(_abc_44694_new_n2244_));
AND2X2 AND2X2_87 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[21] ), .Y(_abc_44694_new_n765_));
AND2X2 AND2X2_870 ( .A(_abc_44694_new_n1940_), .B(_abc_44694_new_n2244_), .Y(_abc_44694_new_n2245_));
AND2X2 AND2X2_871 ( .A(_abc_44694_new_n2246_), .B(_abc_44694_new_n2242_), .Y(_abc_44694_new_n2247_));
AND2X2 AND2X2_872 ( .A(_abc_44694_new_n2089_), .B(_abc_44694_new_n2243_), .Y(_abc_44694_new_n2248_));
AND2X2 AND2X2_873 ( .A(_abc_44694_new_n2210_), .B(_abc_44694_new_n2175_), .Y(_abc_44694_new_n2249_));
AND2X2 AND2X2_874 ( .A(opcode_q_22_), .B(pc_q_24_), .Y(_abc_44694_new_n2255_));
AND2X2 AND2X2_875 ( .A(_abc_44694_new_n2256_), .B(_abc_44694_new_n2254_), .Y(_abc_44694_new_n2257_));
AND2X2 AND2X2_876 ( .A(_abc_44694_new_n2253_), .B(_abc_44694_new_n2257_), .Y(_abc_44694_new_n2259_));
AND2X2 AND2X2_877 ( .A(_abc_44694_new_n2260_), .B(_abc_44694_new_n1194__bF_buf0), .Y(_abc_44694_new_n2261_));
AND2X2 AND2X2_878 ( .A(_abc_44694_new_n2261_), .B(_abc_44694_new_n2258_), .Y(_abc_44694_new_n2262_));
AND2X2 AND2X2_879 ( .A(_abc_44694_new_n1019__bF_buf2), .B(epc_q_24_), .Y(_abc_44694_new_n2263_));
AND2X2 AND2X2_88 ( .A(_abc_44694_new_n766_), .B(_abc_44694_new_n673__bF_buf4), .Y(_abc_44694_new_n767_));
AND2X2 AND2X2_880 ( .A(_abc_44694_new_n2264_), .B(_abc_44694_new_n1340__bF_buf0), .Y(_abc_44694_new_n2265_));
AND2X2 AND2X2_881 ( .A(_abc_44694_new_n1337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_44694_new_n2266_));
AND2X2 AND2X2_882 ( .A(_abc_44694_new_n2269_), .B(_abc_44694_new_n2268_), .Y(_abc_44694_new_n2270_));
AND2X2 AND2X2_883 ( .A(_abc_44694_new_n1522__bF_buf0), .B(epc_q_24_), .Y(_abc_44694_new_n2272_));
AND2X2 AND2X2_884 ( .A(_abc_44694_new_n1348__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_44694_new_n2273_));
AND2X2 AND2X2_885 ( .A(_abc_44694_new_n1207__bF_buf1), .B(_abc_44694_new_n2275_), .Y(_abc_44694_new_n2276_));
AND2X2 AND2X2_886 ( .A(_abc_44694_new_n2271_), .B(_abc_44694_new_n2276_), .Y(_abc_44694_new_n2277_));
AND2X2 AND2X2_887 ( .A(_abc_44694_new_n2279_), .B(enable_i_bF_buf7), .Y(_abc_44694_new_n2280_));
AND2X2 AND2X2_888 ( .A(_abc_44694_new_n2278_), .B(_abc_44694_new_n2280_), .Y(_0epc_q_31_0__24_));
AND2X2 AND2X2_889 ( .A(_abc_44694_new_n2237_), .B(pc_q_25_), .Y(_abc_44694_new_n2283_));
AND2X2 AND2X2_89 ( .A(_abc_44694_new_n681_), .B(\mem_dat_i[29] ), .Y(_abc_44694_new_n768_));
AND2X2 AND2X2_890 ( .A(_abc_44694_new_n2284_), .B(_abc_44694_new_n2282_), .Y(_abc_44694_new_n2285_));
AND2X2 AND2X2_891 ( .A(_abc_44694_new_n2285_), .B(_abc_44694_new_n1382__bF_buf0), .Y(_abc_44694_new_n2286_));
AND2X2 AND2X2_892 ( .A(opcode_q_23_), .B(pc_q_25_), .Y(_abc_44694_new_n2289_));
AND2X2 AND2X2_893 ( .A(_abc_44694_new_n2290_), .B(_abc_44694_new_n2288_), .Y(_abc_44694_new_n2291_));
AND2X2 AND2X2_894 ( .A(_abc_44694_new_n2257_), .B(_abc_44694_new_n2291_), .Y(_abc_44694_new_n2294_));
AND2X2 AND2X2_895 ( .A(_abc_44694_new_n2253_), .B(_abc_44694_new_n2294_), .Y(_abc_44694_new_n2295_));
AND2X2 AND2X2_896 ( .A(_abc_44694_new_n2291_), .B(_abc_44694_new_n2255_), .Y(_abc_44694_new_n2297_));
AND2X2 AND2X2_897 ( .A(_abc_44694_new_n1194__bF_buf4), .B(_abc_44694_new_n2298_), .Y(_abc_44694_new_n2299_));
AND2X2 AND2X2_898 ( .A(_abc_44694_new_n2296_), .B(_abc_44694_new_n2299_), .Y(_abc_44694_new_n2300_));
AND2X2 AND2X2_899 ( .A(_abc_44694_new_n2300_), .B(_abc_44694_new_n2293_), .Y(_abc_44694_new_n2301_));
AND2X2 AND2X2_9 ( .A(inst_r_4_), .B(inst_r_5_), .Y(_abc_44694_new_n633_));
AND2X2 AND2X2_90 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[13] ), .Y(_abc_44694_new_n769_));
AND2X2 AND2X2_900 ( .A(_abc_44694_new_n1019__bF_buf1), .B(epc_q_25_), .Y(_abc_44694_new_n2302_));
AND2X2 AND2X2_901 ( .A(_abc_44694_new_n2303_), .B(_abc_44694_new_n1340__bF_buf4), .Y(_abc_44694_new_n2304_));
AND2X2 AND2X2_902 ( .A(_abc_44694_new_n1337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_44694_new_n2305_));
AND2X2 AND2X2_903 ( .A(_abc_44694_new_n2308_), .B(_abc_44694_new_n2307_), .Y(_abc_44694_new_n2309_));
AND2X2 AND2X2_904 ( .A(_abc_44694_new_n1522__bF_buf4), .B(epc_q_25_), .Y(_abc_44694_new_n2311_));
AND2X2 AND2X2_905 ( .A(_abc_44694_new_n1348__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_44694_new_n2312_));
AND2X2 AND2X2_906 ( .A(_abc_44694_new_n1207__bF_buf0), .B(_abc_44694_new_n2314_), .Y(_abc_44694_new_n2315_));
AND2X2 AND2X2_907 ( .A(_abc_44694_new_n2310_), .B(_abc_44694_new_n2315_), .Y(_abc_44694_new_n2316_));
AND2X2 AND2X2_908 ( .A(_abc_44694_new_n2318_), .B(enable_i_bF_buf6), .Y(_abc_44694_new_n2319_));
AND2X2 AND2X2_909 ( .A(_abc_44694_new_n2317_), .B(_abc_44694_new_n2319_), .Y(_0epc_q_31_0__25_));
AND2X2 AND2X2_91 ( .A(_abc_44694_new_n689_), .B(\mem_dat_i[21] ), .Y(_abc_44694_new_n771_));
AND2X2 AND2X2_910 ( .A(_abc_44694_new_n2283_), .B(pc_q_26_), .Y(_abc_44694_new_n2322_));
AND2X2 AND2X2_911 ( .A(_abc_44694_new_n2323_), .B(_abc_44694_new_n2321_), .Y(_abc_44694_new_n2324_));
AND2X2 AND2X2_912 ( .A(_abc_44694_new_n2324_), .B(_abc_44694_new_n1382__bF_buf3), .Y(_abc_44694_new_n2325_));
AND2X2 AND2X2_913 ( .A(_abc_44694_new_n2298_), .B(_abc_44694_new_n2290_), .Y(_abc_44694_new_n2327_));
AND2X2 AND2X2_914 ( .A(opcode_q_24_), .B(pc_q_26_), .Y(_abc_44694_new_n2331_));
AND2X2 AND2X2_915 ( .A(_abc_44694_new_n2332_), .B(_abc_44694_new_n2330_), .Y(_abc_44694_new_n2333_));
AND2X2 AND2X2_916 ( .A(_abc_44694_new_n2329_), .B(_abc_44694_new_n2333_), .Y(_abc_44694_new_n2335_));
AND2X2 AND2X2_917 ( .A(_abc_44694_new_n2336_), .B(_abc_44694_new_n1194__bF_buf3), .Y(_abc_44694_new_n2337_));
AND2X2 AND2X2_918 ( .A(_abc_44694_new_n2337_), .B(_abc_44694_new_n2334_), .Y(_abc_44694_new_n2338_));
AND2X2 AND2X2_919 ( .A(_abc_44694_new_n1019__bF_buf0), .B(epc_q_26_), .Y(_abc_44694_new_n2339_));
AND2X2 AND2X2_92 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[5] ), .Y(_abc_44694_new_n772_));
AND2X2 AND2X2_920 ( .A(_abc_44694_new_n2340_), .B(_abc_44694_new_n1340__bF_buf3), .Y(_abc_44694_new_n2341_));
AND2X2 AND2X2_921 ( .A(_abc_44694_new_n1337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_44694_new_n2342_));
AND2X2 AND2X2_922 ( .A(_abc_44694_new_n2345_), .B(_abc_44694_new_n2344_), .Y(_abc_44694_new_n2346_));
AND2X2 AND2X2_923 ( .A(_abc_44694_new_n1522__bF_buf3), .B(epc_q_26_), .Y(_abc_44694_new_n2348_));
AND2X2 AND2X2_924 ( .A(_abc_44694_new_n1348__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_44694_new_n2349_));
AND2X2 AND2X2_925 ( .A(_abc_44694_new_n1207__bF_buf5), .B(_abc_44694_new_n2351_), .Y(_abc_44694_new_n2352_));
AND2X2 AND2X2_926 ( .A(_abc_44694_new_n2347_), .B(_abc_44694_new_n2352_), .Y(_abc_44694_new_n2353_));
AND2X2 AND2X2_927 ( .A(_abc_44694_new_n2355_), .B(enable_i_bF_buf5), .Y(_abc_44694_new_n2356_));
AND2X2 AND2X2_928 ( .A(_abc_44694_new_n2354_), .B(_abc_44694_new_n2356_), .Y(_0epc_q_31_0__26_));
AND2X2 AND2X2_929 ( .A(_abc_44694_new_n2322_), .B(pc_q_27_), .Y(_abc_44694_new_n2359_));
AND2X2 AND2X2_93 ( .A(_abc_44694_new_n774_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n775_));
AND2X2 AND2X2_930 ( .A(_abc_44694_new_n2360_), .B(_abc_44694_new_n2358_), .Y(_abc_44694_new_n2361_));
AND2X2 AND2X2_931 ( .A(_abc_44694_new_n2361_), .B(_abc_44694_new_n1382__bF_buf2), .Y(_abc_44694_new_n2362_));
AND2X2 AND2X2_932 ( .A(opcode_q_25_), .B(pc_q_27_), .Y(_abc_44694_new_n2365_));
AND2X2 AND2X2_933 ( .A(_abc_44694_new_n2366_), .B(_abc_44694_new_n2364_), .Y(_abc_44694_new_n2367_));
AND2X2 AND2X2_934 ( .A(_abc_44694_new_n2333_), .B(_abc_44694_new_n2367_), .Y(_abc_44694_new_n2370_));
AND2X2 AND2X2_935 ( .A(_abc_44694_new_n2329_), .B(_abc_44694_new_n2370_), .Y(_abc_44694_new_n2371_));
AND2X2 AND2X2_936 ( .A(_abc_44694_new_n2367_), .B(_abc_44694_new_n2331_), .Y(_abc_44694_new_n2373_));
AND2X2 AND2X2_937 ( .A(_abc_44694_new_n1194__bF_buf2), .B(_abc_44694_new_n2374_), .Y(_abc_44694_new_n2375_));
AND2X2 AND2X2_938 ( .A(_abc_44694_new_n2372_), .B(_abc_44694_new_n2375_), .Y(_abc_44694_new_n2376_));
AND2X2 AND2X2_939 ( .A(_abc_44694_new_n2376_), .B(_abc_44694_new_n2369_), .Y(_abc_44694_new_n2377_));
AND2X2 AND2X2_94 ( .A(_abc_44694_new_n776_), .B(state_q_1_bF_buf1_), .Y(_abc_44694_new_n777_));
AND2X2 AND2X2_940 ( .A(_abc_44694_new_n1019__bF_buf4), .B(epc_q_27_), .Y(_abc_44694_new_n2378_));
AND2X2 AND2X2_941 ( .A(_abc_44694_new_n2379_), .B(_abc_44694_new_n1340__bF_buf2), .Y(_abc_44694_new_n2380_));
AND2X2 AND2X2_942 ( .A(_abc_44694_new_n1337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_44694_new_n2381_));
AND2X2 AND2X2_943 ( .A(_abc_44694_new_n2384_), .B(_abc_44694_new_n2383_), .Y(_abc_44694_new_n2385_));
AND2X2 AND2X2_944 ( .A(_abc_44694_new_n1522__bF_buf2), .B(epc_q_27_), .Y(_abc_44694_new_n2387_));
AND2X2 AND2X2_945 ( .A(_abc_44694_new_n1348__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_44694_new_n2388_));
AND2X2 AND2X2_946 ( .A(_abc_44694_new_n1207__bF_buf4), .B(_abc_44694_new_n2390_), .Y(_abc_44694_new_n2391_));
AND2X2 AND2X2_947 ( .A(_abc_44694_new_n2386_), .B(_abc_44694_new_n2391_), .Y(_abc_44694_new_n2392_));
AND2X2 AND2X2_948 ( .A(_abc_44694_new_n2394_), .B(enable_i_bF_buf4), .Y(_abc_44694_new_n2395_));
AND2X2 AND2X2_949 ( .A(_abc_44694_new_n2393_), .B(_abc_44694_new_n2395_), .Y(_0epc_q_31_0__27_));
AND2X2 AND2X2_95 ( .A(_abc_44694_new_n671_), .B(alu_p_o_6_), .Y(_abc_44694_new_n779_));
AND2X2 AND2X2_950 ( .A(_abc_44694_new_n2359_), .B(pc_q_28_), .Y(_abc_44694_new_n2398_));
AND2X2 AND2X2_951 ( .A(_abc_44694_new_n2399_), .B(_abc_44694_new_n2397_), .Y(_abc_44694_new_n2400_));
AND2X2 AND2X2_952 ( .A(_abc_44694_new_n2400_), .B(_abc_44694_new_n1382__bF_buf1), .Y(_abc_44694_new_n2401_));
AND2X2 AND2X2_953 ( .A(_abc_44694_new_n2374_), .B(_abc_44694_new_n2366_), .Y(_abc_44694_new_n2403_));
AND2X2 AND2X2_954 ( .A(opcode_q_25_), .B(pc_q_28_), .Y(_abc_44694_new_n2407_));
AND2X2 AND2X2_955 ( .A(_abc_44694_new_n2408_), .B(_abc_44694_new_n2406_), .Y(_abc_44694_new_n2409_));
AND2X2 AND2X2_956 ( .A(_abc_44694_new_n2405_), .B(_abc_44694_new_n2409_), .Y(_abc_44694_new_n2411_));
AND2X2 AND2X2_957 ( .A(_abc_44694_new_n2412_), .B(_abc_44694_new_n1194__bF_buf1), .Y(_abc_44694_new_n2413_));
AND2X2 AND2X2_958 ( .A(_abc_44694_new_n2413_), .B(_abc_44694_new_n2410_), .Y(_abc_44694_new_n2414_));
AND2X2 AND2X2_959 ( .A(_abc_44694_new_n1019__bF_buf3), .B(epc_q_28_), .Y(_abc_44694_new_n2415_));
AND2X2 AND2X2_96 ( .A(_abc_44694_new_n678_), .B(\mem_dat_i[6] ), .Y(_abc_44694_new_n780_));
AND2X2 AND2X2_960 ( .A(_abc_44694_new_n2416_), .B(_abc_44694_new_n1340__bF_buf1), .Y(_abc_44694_new_n2417_));
AND2X2 AND2X2_961 ( .A(_abc_44694_new_n1337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_44694_new_n2418_));
AND2X2 AND2X2_962 ( .A(_abc_44694_new_n2421_), .B(_abc_44694_new_n2420_), .Y(_abc_44694_new_n2422_));
AND2X2 AND2X2_963 ( .A(_abc_44694_new_n1522__bF_buf1), .B(epc_q_28_), .Y(_abc_44694_new_n2424_));
AND2X2 AND2X2_964 ( .A(_abc_44694_new_n1348__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_44694_new_n2425_));
AND2X2 AND2X2_965 ( .A(_abc_44694_new_n1207__bF_buf3), .B(_abc_44694_new_n2427_), .Y(_abc_44694_new_n2428_));
AND2X2 AND2X2_966 ( .A(_abc_44694_new_n2423_), .B(_abc_44694_new_n2428_), .Y(_abc_44694_new_n2429_));
AND2X2 AND2X2_967 ( .A(_abc_44694_new_n2431_), .B(enable_i_bF_buf3), .Y(_abc_44694_new_n2432_));
AND2X2 AND2X2_968 ( .A(_abc_44694_new_n2430_), .B(_abc_44694_new_n2432_), .Y(_0epc_q_31_0__28_));
AND2X2 AND2X2_969 ( .A(_abc_44694_new_n2398_), .B(pc_q_29_), .Y(_abc_44694_new_n2435_));
AND2X2 AND2X2_97 ( .A(_abc_44694_new_n682_), .B(\mem_dat_i[22] ), .Y(_abc_44694_new_n781_));
AND2X2 AND2X2_970 ( .A(_abc_44694_new_n2436_), .B(_abc_44694_new_n2434_), .Y(_abc_44694_new_n2437_));
AND2X2 AND2X2_971 ( .A(_abc_44694_new_n2437_), .B(_abc_44694_new_n1382__bF_buf0), .Y(_abc_44694_new_n2438_));
AND2X2 AND2X2_972 ( .A(_abc_44694_new_n2412_), .B(_abc_44694_new_n2408_), .Y(_abc_44694_new_n2440_));
AND2X2 AND2X2_973 ( .A(opcode_q_25_), .B(pc_q_29_), .Y(_abc_44694_new_n2443_));
AND2X2 AND2X2_974 ( .A(_abc_44694_new_n2444_), .B(_abc_44694_new_n2442_), .Y(_abc_44694_new_n2445_));
AND2X2 AND2X2_975 ( .A(_abc_44694_new_n2448_), .B(_abc_44694_new_n1194__bF_buf0), .Y(_abc_44694_new_n2449_));
AND2X2 AND2X2_976 ( .A(_abc_44694_new_n2449_), .B(_abc_44694_new_n2446_), .Y(_abc_44694_new_n2450_));
AND2X2 AND2X2_977 ( .A(_abc_44694_new_n1019__bF_buf2), .B(epc_q_29_), .Y(_abc_44694_new_n2451_));
AND2X2 AND2X2_978 ( .A(_abc_44694_new_n2453_), .B(_abc_44694_new_n2454_), .Y(_abc_44694_new_n2455_));
AND2X2 AND2X2_979 ( .A(_abc_44694_new_n2457_), .B(_abc_44694_new_n2456_), .Y(_abc_44694_new_n2458_));
AND2X2 AND2X2_98 ( .A(_abc_44694_new_n691_), .B(\mem_dat_i[6] ), .Y(_abc_44694_new_n784_));
AND2X2 AND2X2_980 ( .A(_abc_44694_new_n1522__bF_buf0), .B(epc_q_29_), .Y(_abc_44694_new_n2460_));
AND2X2 AND2X2_981 ( .A(_abc_44694_new_n1348__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_44694_new_n2461_));
AND2X2 AND2X2_982 ( .A(_abc_44694_new_n1207__bF_buf2), .B(_abc_44694_new_n2463_), .Y(_abc_44694_new_n2464_));
AND2X2 AND2X2_983 ( .A(_abc_44694_new_n2459_), .B(_abc_44694_new_n2464_), .Y(_abc_44694_new_n2465_));
AND2X2 AND2X2_984 ( .A(_abc_44694_new_n2467_), .B(enable_i_bF_buf2), .Y(_abc_44694_new_n2468_));
AND2X2 AND2X2_985 ( .A(_abc_44694_new_n2466_), .B(_abc_44694_new_n2468_), .Y(_0epc_q_31_0__29_));
AND2X2 AND2X2_986 ( .A(_abc_44694_new_n2435_), .B(pc_q_30_), .Y(_abc_44694_new_n2471_));
AND2X2 AND2X2_987 ( .A(_abc_44694_new_n2472_), .B(_abc_44694_new_n2470_), .Y(_abc_44694_new_n2473_));
AND2X2 AND2X2_988 ( .A(_abc_44694_new_n2473_), .B(_abc_44694_new_n1382__bF_buf3), .Y(_abc_44694_new_n2474_));
AND2X2 AND2X2_989 ( .A(_abc_44694_new_n2411_), .B(_abc_44694_new_n2445_), .Y(_abc_44694_new_n2476_));
AND2X2 AND2X2_99 ( .A(_abc_44694_new_n675_), .B(\mem_dat_i[14] ), .Y(_abc_44694_new_n785_));
AND2X2 AND2X2_990 ( .A(_abc_44694_new_n2408_), .B(_abc_44694_new_n2444_), .Y(_abc_44694_new_n2477_));
AND2X2 AND2X2_991 ( .A(_abc_44694_new_n2481_), .B(opcode_q_25_), .Y(_abc_44694_new_n2482_));
AND2X2 AND2X2_992 ( .A(_abc_44694_new_n623_), .B(pc_q_30_), .Y(_abc_44694_new_n2484_));
AND2X2 AND2X2_993 ( .A(_abc_44694_new_n2483_), .B(_abc_44694_new_n2485_), .Y(_abc_44694_new_n2486_));
AND2X2 AND2X2_994 ( .A(_abc_44694_new_n2489_), .B(_abc_44694_new_n1194__bF_buf4), .Y(_abc_44694_new_n2490_));
AND2X2 AND2X2_995 ( .A(_abc_44694_new_n2490_), .B(_abc_44694_new_n2487_), .Y(_abc_44694_new_n2491_));
AND2X2 AND2X2_996 ( .A(_abc_44694_new_n1019__bF_buf1), .B(epc_q_30_), .Y(_abc_44694_new_n2492_));
AND2X2 AND2X2_997 ( .A(_abc_44694_new_n2493_), .B(_abc_44694_new_n1340__bF_buf4), .Y(_abc_44694_new_n2494_));
AND2X2 AND2X2_998 ( .A(_abc_44694_new_n1337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_44694_new_n2495_));
AND2X2 AND2X2_999 ( .A(_abc_44694_new_n2498_), .B(_abc_44694_new_n2497_), .Y(_abc_44694_new_n2499_));
BUFX2 BUFX2_1 ( .A(_abc_44694_new_n1186_), .Y(_abc_44694_new_n1186__bF_buf3));
BUFX2 BUFX2_10 ( .A(_abc_44694_new_n3546_), .Y(_abc_44694_new_n3546__bF_buf2));
BUFX2 BUFX2_100 ( .A(1'h1), .Y(\mem_cti_o[0] ));
BUFX2 BUFX2_101 ( .A(1'h1), .Y(\mem_cti_o[1] ));
BUFX2 BUFX2_102 ( .A(1'h1), .Y(\mem_cti_o[2] ));
BUFX2 BUFX2_103 ( .A(_auto_iopadmap_cc_368_execute_48748), .Y(mem_cyc_o));
BUFX2 BUFX2_104 ( .A(_auto_iopadmap_cc_368_execute_48750_0_), .Y(\mem_dat_o[0] ));
BUFX2 BUFX2_105 ( .A(_auto_iopadmap_cc_368_execute_48750_1_), .Y(\mem_dat_o[1] ));
BUFX2 BUFX2_106 ( .A(_auto_iopadmap_cc_368_execute_48750_2_), .Y(\mem_dat_o[2] ));
BUFX2 BUFX2_107 ( .A(_auto_iopadmap_cc_368_execute_48750_3_), .Y(\mem_dat_o[3] ));
BUFX2 BUFX2_108 ( .A(_auto_iopadmap_cc_368_execute_48750_4_), .Y(\mem_dat_o[4] ));
BUFX2 BUFX2_109 ( .A(_auto_iopadmap_cc_368_execute_48750_5_), .Y(\mem_dat_o[5] ));
BUFX2 BUFX2_11 ( .A(_abc_44694_new_n3546_), .Y(_abc_44694_new_n3546__bF_buf1));
BUFX2 BUFX2_110 ( .A(_auto_iopadmap_cc_368_execute_48750_6_), .Y(\mem_dat_o[6] ));
BUFX2 BUFX2_111 ( .A(_auto_iopadmap_cc_368_execute_48750_7_), .Y(\mem_dat_o[7] ));
BUFX2 BUFX2_112 ( .A(_auto_iopadmap_cc_368_execute_48750_8_), .Y(\mem_dat_o[8] ));
BUFX2 BUFX2_113 ( .A(_auto_iopadmap_cc_368_execute_48750_9_), .Y(\mem_dat_o[9] ));
BUFX2 BUFX2_114 ( .A(_auto_iopadmap_cc_368_execute_48750_10_), .Y(\mem_dat_o[10] ));
BUFX2 BUFX2_115 ( .A(_auto_iopadmap_cc_368_execute_48750_11_), .Y(\mem_dat_o[11] ));
BUFX2 BUFX2_116 ( .A(_auto_iopadmap_cc_368_execute_48750_12_), .Y(\mem_dat_o[12] ));
BUFX2 BUFX2_117 ( .A(_auto_iopadmap_cc_368_execute_48750_13_), .Y(\mem_dat_o[13] ));
BUFX2 BUFX2_118 ( .A(_auto_iopadmap_cc_368_execute_48750_14_), .Y(\mem_dat_o[14] ));
BUFX2 BUFX2_119 ( .A(_auto_iopadmap_cc_368_execute_48750_15_), .Y(\mem_dat_o[15] ));
BUFX2 BUFX2_12 ( .A(_abc_44694_new_n3546_), .Y(_abc_44694_new_n3546__bF_buf0));
BUFX2 BUFX2_120 ( .A(_auto_iopadmap_cc_368_execute_48750_16_), .Y(\mem_dat_o[16] ));
BUFX2 BUFX2_121 ( .A(_auto_iopadmap_cc_368_execute_48750_17_), .Y(\mem_dat_o[17] ));
BUFX2 BUFX2_122 ( .A(_auto_iopadmap_cc_368_execute_48750_18_), .Y(\mem_dat_o[18] ));
BUFX2 BUFX2_123 ( .A(_auto_iopadmap_cc_368_execute_48750_19_), .Y(\mem_dat_o[19] ));
BUFX2 BUFX2_124 ( .A(_auto_iopadmap_cc_368_execute_48750_20_), .Y(\mem_dat_o[20] ));
BUFX2 BUFX2_125 ( .A(_auto_iopadmap_cc_368_execute_48750_21_), .Y(\mem_dat_o[21] ));
BUFX2 BUFX2_126 ( .A(_auto_iopadmap_cc_368_execute_48750_22_), .Y(\mem_dat_o[22] ));
BUFX2 BUFX2_127 ( .A(_auto_iopadmap_cc_368_execute_48750_23_), .Y(\mem_dat_o[23] ));
BUFX2 BUFX2_128 ( .A(_auto_iopadmap_cc_368_execute_48750_24_), .Y(\mem_dat_o[24] ));
BUFX2 BUFX2_129 ( .A(_auto_iopadmap_cc_368_execute_48750_25_), .Y(\mem_dat_o[25] ));
BUFX2 BUFX2_13 ( .A(alu__abc_42281_new_n876_), .Y(alu__abc_42281_new_n876__bF_buf3));
BUFX2 BUFX2_130 ( .A(_auto_iopadmap_cc_368_execute_48750_26_), .Y(\mem_dat_o[26] ));
BUFX2 BUFX2_131 ( .A(_auto_iopadmap_cc_368_execute_48750_27_), .Y(\mem_dat_o[27] ));
BUFX2 BUFX2_132 ( .A(_auto_iopadmap_cc_368_execute_48750_28_), .Y(\mem_dat_o[28] ));
BUFX2 BUFX2_133 ( .A(_auto_iopadmap_cc_368_execute_48750_29_), .Y(\mem_dat_o[29] ));
BUFX2 BUFX2_134 ( .A(_auto_iopadmap_cc_368_execute_48750_30_), .Y(\mem_dat_o[30] ));
BUFX2 BUFX2_135 ( .A(_auto_iopadmap_cc_368_execute_48750_31_), .Y(\mem_dat_o[31] ));
BUFX2 BUFX2_136 ( .A(_auto_iopadmap_cc_368_execute_48783_0_), .Y(\mem_sel_o[0] ));
BUFX2 BUFX2_137 ( .A(_auto_iopadmap_cc_368_execute_48783_1_), .Y(\mem_sel_o[1] ));
BUFX2 BUFX2_138 ( .A(_auto_iopadmap_cc_368_execute_48783_2_), .Y(\mem_sel_o[2] ));
BUFX2 BUFX2_139 ( .A(_auto_iopadmap_cc_368_execute_48783_3_), .Y(\mem_sel_o[3] ));
BUFX2 BUFX2_14 ( .A(alu__abc_42281_new_n876_), .Y(alu__abc_42281_new_n876__bF_buf2));
BUFX2 BUFX2_140 ( .A(_auto_iopadmap_cc_368_execute_48788), .Y(mem_stb_o));
BUFX2 BUFX2_141 ( .A(_auto_iopadmap_cc_368_execute_48790), .Y(mem_we_o));
BUFX2 BUFX2_15 ( .A(alu__abc_42281_new_n876_), .Y(alu__abc_42281_new_n876__bF_buf1));
BUFX2 BUFX2_16 ( .A(alu__abc_42281_new_n876_), .Y(alu__abc_42281_new_n876__bF_buf0));
BUFX2 BUFX2_17 ( .A(_abc_44694_new_n1382_), .Y(_abc_44694_new_n1382__bF_buf3));
BUFX2 BUFX2_18 ( .A(_abc_44694_new_n1382_), .Y(_abc_44694_new_n1382__bF_buf2));
BUFX2 BUFX2_19 ( .A(_abc_44694_new_n1382_), .Y(_abc_44694_new_n1382__bF_buf1));
BUFX2 BUFX2_2 ( .A(_abc_44694_new_n1186_), .Y(_abc_44694_new_n1186__bF_buf2));
BUFX2 BUFX2_20 ( .A(_abc_44694_new_n1382_), .Y(_abc_44694_new_n1382__bF_buf0));
BUFX2 BUFX2_21 ( .A(_abc_44694_new_n2546_), .Y(_abc_44694_new_n2546__bF_buf1));
BUFX2 BUFX2_22 ( .A(_abc_44694_new_n2546_), .Y(_abc_44694_new_n2546__bF_buf0));
BUFX2 BUFX2_23 ( .A(_abc_44694_new_n1185_), .Y(_abc_44694_new_n1185__bF_buf2));
BUFX2 BUFX2_24 ( .A(_abc_44694_new_n1185_), .Y(_abc_44694_new_n1185__bF_buf1));
BUFX2 BUFX2_25 ( .A(_abc_44694_new_n1185_), .Y(_abc_44694_new_n1185__bF_buf0));
BUFX2 BUFX2_26 ( .A(_abc_44694_new_n677_), .Y(_abc_44694_new_n677__bF_buf2));
BUFX2 BUFX2_27 ( .A(_abc_44694_new_n677_), .Y(_abc_44694_new_n677__bF_buf1));
BUFX2 BUFX2_28 ( .A(_abc_44694_new_n677_), .Y(_abc_44694_new_n677__bF_buf0));
BUFX2 BUFX2_29 ( .A(_abc_44694_new_n668_), .Y(_abc_44694_new_n668__bF_buf1));
BUFX2 BUFX2_3 ( .A(_abc_44694_new_n1186_), .Y(_abc_44694_new_n1186__bF_buf1));
BUFX2 BUFX2_30 ( .A(_abc_44694_new_n668_), .Y(_abc_44694_new_n668__bF_buf0));
BUFX2 BUFX2_31 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0_));
BUFX2 BUFX2_32 ( .A(_abc_44694_new_n1087_), .Y(_abc_44694_new_n1087__bF_buf1));
BUFX2 BUFX2_33 ( .A(_abc_44694_new_n1087_), .Y(_abc_44694_new_n1087__bF_buf0));
BUFX2 BUFX2_34 ( .A(_abc_44694_new_n3518_), .Y(_abc_44694_new_n3518__bF_buf0));
BUFX2 BUFX2_35 ( .A(_abc_44694_new_n1181_), .Y(_abc_44694_new_n1181__bF_buf1));
BUFX2 BUFX2_36 ( .A(_abc_44694_new_n1181_), .Y(_abc_44694_new_n1181__bF_buf0));
BUFX2 BUFX2_37 ( .A(_abc_44694_new_n1084_), .Y(_abc_44694_new_n1084__bF_buf1));
BUFX2 BUFX2_38 ( .A(_abc_44694_new_n1084_), .Y(_abc_44694_new_n1084__bF_buf0));
BUFX2 BUFX2_39 ( .A(_abc_44694_new_n3515_), .Y(_abc_44694_new_n3515__bF_buf3));
BUFX2 BUFX2_4 ( .A(_abc_44694_new_n1186_), .Y(_abc_44694_new_n1186__bF_buf0));
BUFX2 BUFX2_40 ( .A(_abc_44694_new_n3515_), .Y(_abc_44694_new_n3515__bF_buf2));
BUFX2 BUFX2_41 ( .A(_abc_44694_new_n3515_), .Y(_abc_44694_new_n3515__bF_buf1));
BUFX2 BUFX2_42 ( .A(_abc_44694_new_n3515_), .Y(_abc_44694_new_n3515__bF_buf0));
BUFX2 BUFX2_43 ( .A(_abc_44694_new_n1522_), .Y(_abc_44694_new_n1522__bF_buf2));
BUFX2 BUFX2_44 ( .A(_abc_44694_new_n1522_), .Y(_abc_44694_new_n1522__bF_buf1));
BUFX2 BUFX2_45 ( .A(_abc_44694_new_n1522_), .Y(_abc_44694_new_n1522__bF_buf0));
BUFX2 BUFX2_46 ( .A(state_q_5_), .Y(state_q_5_bF_buf3_));
BUFX2 BUFX2_47 ( .A(state_q_5_), .Y(state_q_5_bF_buf2_));
BUFX2 BUFX2_48 ( .A(state_q_5_), .Y(state_q_5_bF_buf1_));
BUFX2 BUFX2_49 ( .A(alu__abc_42281_new_n936_), .Y(alu__abc_42281_new_n936__bF_buf4));
BUFX2 BUFX2_5 ( .A(_abc_44694_new_n2826_), .Y(_abc_44694_new_n2826__bF_buf3));
BUFX2 BUFX2_50 ( .A(alu__abc_42281_new_n936_), .Y(alu__abc_42281_new_n936__bF_buf3));
BUFX2 BUFX2_51 ( .A(alu__abc_42281_new_n936_), .Y(alu__abc_42281_new_n936__bF_buf2));
BUFX2 BUFX2_52 ( .A(alu__abc_42281_new_n936_), .Y(alu__abc_42281_new_n936__bF_buf1));
BUFX2 BUFX2_53 ( .A(alu__abc_42281_new_n936_), .Y(alu__abc_42281_new_n936__bF_buf0));
BUFX2 BUFX2_54 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_));
BUFX2 BUFX2_55 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank_ra_i_4_bF_buf2_));
BUFX2 BUFX2_56 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank_ra_i_4_bF_buf1_));
BUFX2 BUFX2_57 ( .A(_abc_44694_new_n2779_), .Y(_abc_44694_new_n2779__bF_buf3));
BUFX2 BUFX2_58 ( .A(_abc_44694_new_n2779_), .Y(_abc_44694_new_n2779__bF_buf2));
BUFX2 BUFX2_59 ( .A(_abc_44694_new_n2779_), .Y(_abc_44694_new_n2779__bF_buf1));
BUFX2 BUFX2_6 ( .A(_abc_44694_new_n2826_), .Y(_abc_44694_new_n2826__bF_buf2));
BUFX2 BUFX2_60 ( .A(_abc_44694_new_n2779_), .Y(_abc_44694_new_n2779__bF_buf0));
BUFX2 BUFX2_61 ( .A(_abc_44694_new_n4064_), .Y(_abc_44694_new_n4064__bF_buf4));
BUFX2 BUFX2_62 ( .A(_abc_44694_new_n4064_), .Y(_abc_44694_new_n4064__bF_buf3));
BUFX2 BUFX2_63 ( .A(_abc_44694_new_n4064_), .Y(_abc_44694_new_n4064__bF_buf2));
BUFX2 BUFX2_64 ( .A(_abc_44694_new_n4064_), .Y(_abc_44694_new_n4064__bF_buf1));
BUFX2 BUFX2_65 ( .A(_abc_44694_new_n4064_), .Y(_abc_44694_new_n4064__bF_buf0));
BUFX2 BUFX2_66 ( .A(_auto_iopadmap_cc_368_execute_48707), .Y(break_o));
BUFX2 BUFX2_67 ( .A(_auto_iopadmap_cc_368_execute_48709), .Y(fault_o));
BUFX2 BUFX2_68 ( .A(_auto_iopadmap_cc_368_execute_48711_0_), .Y(\mem_addr_o[0] ));
BUFX2 BUFX2_69 ( .A(_auto_iopadmap_cc_368_execute_48711_1_), .Y(\mem_addr_o[1] ));
BUFX2 BUFX2_7 ( .A(_abc_44694_new_n2826_), .Y(_abc_44694_new_n2826__bF_buf1));
BUFX2 BUFX2_70 ( .A(_auto_iopadmap_cc_368_execute_48711_2_), .Y(\mem_addr_o[2] ));
BUFX2 BUFX2_71 ( .A(_auto_iopadmap_cc_368_execute_48711_3_), .Y(\mem_addr_o[3] ));
BUFX2 BUFX2_72 ( .A(_auto_iopadmap_cc_368_execute_48711_4_), .Y(\mem_addr_o[4] ));
BUFX2 BUFX2_73 ( .A(_auto_iopadmap_cc_368_execute_48711_5_), .Y(\mem_addr_o[5] ));
BUFX2 BUFX2_74 ( .A(_auto_iopadmap_cc_368_execute_48711_6_), .Y(\mem_addr_o[6] ));
BUFX2 BUFX2_75 ( .A(_auto_iopadmap_cc_368_execute_48711_7_), .Y(\mem_addr_o[7] ));
BUFX2 BUFX2_76 ( .A(_auto_iopadmap_cc_368_execute_48711_8_), .Y(\mem_addr_o[8] ));
BUFX2 BUFX2_77 ( .A(_auto_iopadmap_cc_368_execute_48711_9_), .Y(\mem_addr_o[9] ));
BUFX2 BUFX2_78 ( .A(_auto_iopadmap_cc_368_execute_48711_10_), .Y(\mem_addr_o[10] ));
BUFX2 BUFX2_79 ( .A(_auto_iopadmap_cc_368_execute_48711_11_), .Y(\mem_addr_o[11] ));
BUFX2 BUFX2_8 ( .A(_abc_44694_new_n2826_), .Y(_abc_44694_new_n2826__bF_buf0));
BUFX2 BUFX2_80 ( .A(_auto_iopadmap_cc_368_execute_48711_12_), .Y(\mem_addr_o[12] ));
BUFX2 BUFX2_81 ( .A(_auto_iopadmap_cc_368_execute_48711_13_), .Y(\mem_addr_o[13] ));
BUFX2 BUFX2_82 ( .A(_auto_iopadmap_cc_368_execute_48711_14_), .Y(\mem_addr_o[14] ));
BUFX2 BUFX2_83 ( .A(_auto_iopadmap_cc_368_execute_48711_15_), .Y(\mem_addr_o[15] ));
BUFX2 BUFX2_84 ( .A(_auto_iopadmap_cc_368_execute_48711_16_), .Y(\mem_addr_o[16] ));
BUFX2 BUFX2_85 ( .A(_auto_iopadmap_cc_368_execute_48711_17_), .Y(\mem_addr_o[17] ));
BUFX2 BUFX2_86 ( .A(_auto_iopadmap_cc_368_execute_48711_18_), .Y(\mem_addr_o[18] ));
BUFX2 BUFX2_87 ( .A(_auto_iopadmap_cc_368_execute_48711_19_), .Y(\mem_addr_o[19] ));
BUFX2 BUFX2_88 ( .A(_auto_iopadmap_cc_368_execute_48711_20_), .Y(\mem_addr_o[20] ));
BUFX2 BUFX2_89 ( .A(_auto_iopadmap_cc_368_execute_48711_21_), .Y(\mem_addr_o[21] ));
BUFX2 BUFX2_9 ( .A(_abc_44694_new_n3546_), .Y(_abc_44694_new_n3546__bF_buf3));
BUFX2 BUFX2_90 ( .A(_auto_iopadmap_cc_368_execute_48711_22_), .Y(\mem_addr_o[22] ));
BUFX2 BUFX2_91 ( .A(_auto_iopadmap_cc_368_execute_48711_23_), .Y(\mem_addr_o[23] ));
BUFX2 BUFX2_92 ( .A(_auto_iopadmap_cc_368_execute_48711_24_), .Y(\mem_addr_o[24] ));
BUFX2 BUFX2_93 ( .A(_auto_iopadmap_cc_368_execute_48711_25_), .Y(\mem_addr_o[25] ));
BUFX2 BUFX2_94 ( .A(_auto_iopadmap_cc_368_execute_48711_26_), .Y(\mem_addr_o[26] ));
BUFX2 BUFX2_95 ( .A(_auto_iopadmap_cc_368_execute_48711_27_), .Y(\mem_addr_o[27] ));
BUFX2 BUFX2_96 ( .A(_auto_iopadmap_cc_368_execute_48711_28_), .Y(\mem_addr_o[28] ));
BUFX2 BUFX2_97 ( .A(_auto_iopadmap_cc_368_execute_48711_29_), .Y(\mem_addr_o[29] ));
BUFX2 BUFX2_98 ( .A(_auto_iopadmap_cc_368_execute_48711_30_), .Y(\mem_addr_o[30] ));
BUFX2 BUFX2_99 ( .A(_auto_iopadmap_cc_368_execute_48711_31_), .Y(\mem_addr_o[31] ));
BUFX4 BUFX4_1 ( .A(clk_i), .Y(clk_i_hier0_bF_buf9));
BUFX4 BUFX4_10 ( .A(clk_i), .Y(clk_i_hier0_bF_buf0));
BUFX4 BUFX4_100 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_));
BUFX4 BUFX4_1000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf1));
BUFX4 BUFX4_1001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf0));
BUFX4 BUFX4_1002 ( .A(_abc_44694_new_n673_), .Y(_abc_44694_new_n673__bF_buf4));
BUFX4 BUFX4_1003 ( .A(_abc_44694_new_n673_), .Y(_abc_44694_new_n673__bF_buf3));
BUFX4 BUFX4_1004 ( .A(_abc_44694_new_n673_), .Y(_abc_44694_new_n673__bF_buf2));
BUFX4 BUFX4_1005 ( .A(_abc_44694_new_n673_), .Y(_abc_44694_new_n673__bF_buf1));
BUFX4 BUFX4_1006 ( .A(_abc_44694_new_n673_), .Y(_abc_44694_new_n673__bF_buf0));
BUFX4 BUFX4_1007 ( .A(_abc_44694_new_n1084_), .Y(_abc_44694_new_n1084__bF_buf3));
BUFX4 BUFX4_1008 ( .A(_abc_44694_new_n1084_), .Y(_abc_44694_new_n1084__bF_buf2));
BUFX4 BUFX4_1009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf4));
BUFX4 BUFX4_101 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_));
BUFX4 BUFX4_1010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf3));
BUFX4 BUFX4_1011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf2));
BUFX4 BUFX4_1012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf1));
BUFX4 BUFX4_1013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5585__bF_buf0));
BUFX4 BUFX4_1014 ( .A(_abc_44694_new_n1178_), .Y(_abc_44694_new_n1178__bF_buf4));
BUFX4 BUFX4_1015 ( .A(_abc_44694_new_n1178_), .Y(_abc_44694_new_n1178__bF_buf3));
BUFX4 BUFX4_1016 ( .A(_abc_44694_new_n1178_), .Y(_abc_44694_new_n1178__bF_buf2));
BUFX4 BUFX4_1017 ( .A(_abc_44694_new_n1178_), .Y(_abc_44694_new_n1178__bF_buf1));
BUFX4 BUFX4_1018 ( .A(_abc_44694_new_n1178_), .Y(_abc_44694_new_n1178__bF_buf0));
BUFX4 BUFX4_1019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4));
BUFX4 BUFX4_102 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_));
BUFX4 BUFX4_1020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3));
BUFX4 BUFX4_1021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2));
BUFX4 BUFX4_1022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1));
BUFX4 BUFX4_1023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0));
BUFX4 BUFX4_1024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4));
BUFX4 BUFX4_1025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3));
BUFX4 BUFX4_1026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2));
BUFX4 BUFX4_1027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1));
BUFX4 BUFX4_1028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0));
BUFX4 BUFX4_1029 ( .A(_abc_44694_new_n1522_), .Y(_abc_44694_new_n1522__bF_buf4));
BUFX4 BUFX4_103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7));
BUFX4 BUFX4_1030 ( .A(_abc_44694_new_n1522_), .Y(_abc_44694_new_n1522__bF_buf3));
BUFX4 BUFX4_1031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4));
BUFX4 BUFX4_1032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3));
BUFX4 BUFX4_1033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2));
BUFX4 BUFX4_1034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1));
BUFX4 BUFX4_1035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0));
BUFX4 BUFX4_1036 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_));
BUFX4 BUFX4_1037 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_));
BUFX4 BUFX4_1038 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_));
BUFX4 BUFX4_1039 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_));
BUFX4 BUFX4_104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf6));
BUFX4 BUFX4_1040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf4));
BUFX4 BUFX4_1041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf3));
BUFX4 BUFX4_1042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf2));
BUFX4 BUFX4_1043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf1));
BUFX4 BUFX4_1044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5603_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5603__bF_buf0));
BUFX4 BUFX4_1045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf4));
BUFX4 BUFX4_1046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf3));
BUFX4 BUFX4_1047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf2));
BUFX4 BUFX4_1048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf1));
BUFX4 BUFX4_1049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7575__bF_buf0));
BUFX4 BUFX4_105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5));
BUFX4 BUFX4_1050 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf6));
BUFX4 BUFX4_1051 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf5));
BUFX4 BUFX4_1052 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf4));
BUFX4 BUFX4_1053 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf3));
BUFX4 BUFX4_1054 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf2));
BUFX4 BUFX4_1055 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf1));
BUFX4 BUFX4_1056 ( .A(alu__abc_42281_new_n281_), .Y(alu__abc_42281_new_n281__bF_buf0));
BUFX4 BUFX4_1057 ( .A(_abc_44694_new_n3512_), .Y(_abc_44694_new_n3512__bF_buf4));
BUFX4 BUFX4_1058 ( .A(_abc_44694_new_n3512_), .Y(_abc_44694_new_n3512__bF_buf3));
BUFX4 BUFX4_1059 ( .A(_abc_44694_new_n3512_), .Y(_abc_44694_new_n3512__bF_buf2));
BUFX4 BUFX4_106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf4));
BUFX4 BUFX4_1060 ( .A(_abc_44694_new_n3512_), .Y(_abc_44694_new_n3512__bF_buf1));
BUFX4 BUFX4_1061 ( .A(_abc_44694_new_n3512_), .Y(_abc_44694_new_n3512__bF_buf0));
BUFX4 BUFX4_1062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf4));
BUFX4 BUFX4_1063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf3));
BUFX4 BUFX4_1064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf2));
BUFX4 BUFX4_1065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf1));
BUFX4 BUFX4_1066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5582__bF_buf0));
BUFX4 BUFX4_1067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf4));
BUFX4 BUFX4_1068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf3));
BUFX4 BUFX4_1069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf2));
BUFX4 BUFX4_107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3));
BUFX4 BUFX4_1070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf1));
BUFX4 BUFX4_1071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5638__bF_buf0));
BUFX4 BUFX4_1072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7));
BUFX4 BUFX4_1073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf6));
BUFX4 BUFX4_1074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5));
BUFX4 BUFX4_1075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf4));
BUFX4 BUFX4_1076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3));
BUFX4 BUFX4_1077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf2));
BUFX4 BUFX4_1078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1));
BUFX4 BUFX4_1079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf0));
BUFX4 BUFX4_108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf2));
BUFX4 BUFX4_1080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4));
BUFX4 BUFX4_1081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3));
BUFX4 BUFX4_1082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2));
BUFX4 BUFX4_1083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1));
BUFX4 BUFX4_1084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0));
BUFX4 BUFX4_1085 ( .A(state_q_5_), .Y(state_q_5_bF_buf0_));
BUFX4 BUFX4_1086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf4));
BUFX4 BUFX4_1087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf3));
BUFX4 BUFX4_1088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf2));
BUFX4 BUFX4_1089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf1));
BUFX4 BUFX4_109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1));
BUFX4 BUFX4_1090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7631_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7631__bF_buf0));
BUFX4 BUFX4_1091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4));
BUFX4 BUFX4_1092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3));
BUFX4 BUFX4_1093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2));
BUFX4 BUFX4_1094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1));
BUFX4 BUFX4_1095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0));
BUFX4 BUFX4_1096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf4));
BUFX4 BUFX4_1097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf3));
BUFX4 BUFX4_1098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf2));
BUFX4 BUFX4_1099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf1));
BUFX4 BUFX4_11 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3));
BUFX4 BUFX4_110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf0));
BUFX4 BUFX4_1100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5600__bF_buf0));
BUFX4 BUFX4_1101 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7));
BUFX4 BUFX4_1102 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf6));
BUFX4 BUFX4_1103 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5));
BUFX4 BUFX4_1104 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf4));
BUFX4 BUFX4_1105 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3));
BUFX4 BUFX4_1106 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf2));
BUFX4 BUFX4_1107 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1));
BUFX4 BUFX4_1108 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424), .Y(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf0));
BUFX4 BUFX4_1109 ( .A(_abc_44694_new_n817_), .Y(_abc_44694_new_n817__bF_buf3));
BUFX4 BUFX4_111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf4));
BUFX4 BUFX4_1110 ( .A(_abc_44694_new_n817_), .Y(_abc_44694_new_n817__bF_buf2));
BUFX4 BUFX4_1111 ( .A(_abc_44694_new_n817_), .Y(_abc_44694_new_n817__bF_buf1));
BUFX4 BUFX4_1112 ( .A(_abc_44694_new_n817_), .Y(_abc_44694_new_n817__bF_buf0));
BUFX4 BUFX4_1113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf4));
BUFX4 BUFX4_1114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf3));
BUFX4 BUFX4_1115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf2));
BUFX4 BUFX4_1116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf1));
BUFX4 BUFX4_1117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5635_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5635__bF_buf0));
BUFX4 BUFX4_1118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4));
BUFX4 BUFX4_1119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3));
BUFX4 BUFX4_112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf3));
BUFX4 BUFX4_1120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2));
BUFX4 BUFX4_1121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1));
BUFX4 BUFX4_1122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0));
BUFX4 BUFX4_1123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4));
BUFX4 BUFX4_1124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3));
BUFX4 BUFX4_1125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2));
BUFX4 BUFX4_1126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1));
BUFX4 BUFX4_1127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0));
BUFX4 BUFX4_1128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf4));
BUFX4 BUFX4_1129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf3));
BUFX4 BUFX4_113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf2));
BUFX4 BUFX4_1130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf2));
BUFX4 BUFX4_1131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf1));
BUFX4 BUFX4_1132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7625_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7625__bF_buf0));
BUFX4 BUFX4_1133 ( .A(alu__abc_42281_new_n942_), .Y(alu__abc_42281_new_n942__bF_buf4));
BUFX4 BUFX4_1134 ( .A(alu__abc_42281_new_n942_), .Y(alu__abc_42281_new_n942__bF_buf3));
BUFX4 BUFX4_1135 ( .A(alu__abc_42281_new_n942_), .Y(alu__abc_42281_new_n942__bF_buf2));
BUFX4 BUFX4_1136 ( .A(alu__abc_42281_new_n942_), .Y(alu__abc_42281_new_n942__bF_buf1));
BUFX4 BUFX4_1137 ( .A(alu__abc_42281_new_n942_), .Y(alu__abc_42281_new_n942__bF_buf0));
BUFX4 BUFX4_1138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4));
BUFX4 BUFX4_1139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3));
BUFX4 BUFX4_114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf1));
BUFX4 BUFX4_1140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2));
BUFX4 BUFX4_1141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1));
BUFX4 BUFX4_1142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0));
BUFX4 BUFX4_1143 ( .A(alu__abc_42281_new_n939_), .Y(alu__abc_42281_new_n939__bF_buf4));
BUFX4 BUFX4_1144 ( .A(alu__abc_42281_new_n939_), .Y(alu__abc_42281_new_n939__bF_buf3));
BUFX4 BUFX4_1145 ( .A(alu__abc_42281_new_n939_), .Y(alu__abc_42281_new_n939__bF_buf2));
BUFX4 BUFX4_1146 ( .A(alu__abc_42281_new_n939_), .Y(alu__abc_42281_new_n939__bF_buf1));
BUFX4 BUFX4_1147 ( .A(alu__abc_42281_new_n939_), .Y(alu__abc_42281_new_n939__bF_buf0));
BUFX4 BUFX4_1148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4));
BUFX4 BUFX4_1149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3));
BUFX4 BUFX4_115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7633__bF_buf0));
BUFX4 BUFX4_1150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2));
BUFX4 BUFX4_1151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1));
BUFX4 BUFX4_1152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0));
BUFX4 BUFX4_1153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4));
BUFX4 BUFX4_1154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3));
BUFX4 BUFX4_1155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2));
BUFX4 BUFX4_1156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1));
BUFX4 BUFX4_1157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0));
BUFX4 BUFX4_1158 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf7));
BUFX4 BUFX4_1159 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf6));
BUFX4 BUFX4_116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7));
BUFX4 BUFX4_1160 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf5));
BUFX4 BUFX4_1161 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf4));
BUFX4 BUFX4_1162 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf3));
BUFX4 BUFX4_1163 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf2));
BUFX4 BUFX4_1164 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf1));
BUFX4 BUFX4_1165 ( .A(REGFILE_SIM_reg_bank_wr_i), .Y(REGFILE_SIM_reg_bank_wr_i_bF_buf0));
BUFX4 BUFX4_1166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf4));
BUFX4 BUFX4_1167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf3));
BUFX4 BUFX4_1168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf2));
BUFX4 BUFX4_1169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf1));
BUFX4 BUFX4_117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf6));
BUFX4 BUFX4_1170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7619_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7619__bF_buf0));
BUFX4 BUFX4_1171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf4));
BUFX4 BUFX4_1172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf3));
BUFX4 BUFX4_1173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf2));
BUFX4 BUFX4_1174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf1));
BUFX4 BUFX4_1175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5626_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5626__bF_buf0));
BUFX4 BUFX4_1176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf4));
BUFX4 BUFX4_1177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf3));
BUFX4 BUFX4_1178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf2));
BUFX4 BUFX4_1179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf1));
BUFX4 BUFX4_118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5));
BUFX4 BUFX4_1180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7598__bF_buf0));
BUFX4 BUFX4_1181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf4));
BUFX4 BUFX4_1182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf3));
BUFX4 BUFX4_1183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf2));
BUFX4 BUFX4_1184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf1));
BUFX4 BUFX4_1185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7654_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7654__bF_buf0));
BUFX4 BUFX4_1186 ( .A(REGFILE_SIM_reg_bank_ra_i_4_), .Y(REGFILE_SIM_reg_bank_ra_i_4_bF_buf0_));
BUFX4 BUFX4_1187 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf6_));
BUFX4 BUFX4_1188 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf5_));
BUFX4 BUFX4_1189 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf4_));
BUFX4 BUFX4_119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf4));
BUFX4 BUFX4_1190 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf3_));
BUFX4 BUFX4_1191 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf2_));
BUFX4 BUFX4_1192 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf1_));
BUFX4 BUFX4_1193 ( .A(alu_b_i_3_), .Y(alu_b_i_3_bF_buf0_));
BUFX4 BUFX4_1194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf4));
BUFX4 BUFX4_1195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf3));
BUFX4 BUFX4_1196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf2));
BUFX4 BUFX4_1197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf1));
BUFX4 BUFX4_1198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5623__bF_buf0));
BUFX4 BUFX4_1199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf4));
BUFX4 BUFX4_12 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf2));
BUFX4 BUFX4_120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3));
BUFX4 BUFX4_1200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf3));
BUFX4 BUFX4_1201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf2));
BUFX4 BUFX4_1202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf1));
BUFX4 BUFX4_1203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7595_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7595__bF_buf0));
BUFX4 BUFX4_1204 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_));
BUFX4 BUFX4_1205 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_));
BUFX4 BUFX4_1206 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_));
BUFX4 BUFX4_1207 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_));
BUFX4 BUFX4_1208 ( .A(_abc_44694_new_n1348_), .Y(_abc_44694_new_n1348__bF_buf5));
BUFX4 BUFX4_1209 ( .A(_abc_44694_new_n1348_), .Y(_abc_44694_new_n1348__bF_buf4));
BUFX4 BUFX4_121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf2));
BUFX4 BUFX4_1210 ( .A(_abc_44694_new_n1348_), .Y(_abc_44694_new_n1348__bF_buf3));
BUFX4 BUFX4_1211 ( .A(_abc_44694_new_n1348_), .Y(_abc_44694_new_n1348__bF_buf2));
BUFX4 BUFX4_1212 ( .A(_abc_44694_new_n1348_), .Y(_abc_44694_new_n1348__bF_buf1));
BUFX4 BUFX4_1213 ( .A(_abc_44694_new_n1348_), .Y(_abc_44694_new_n1348__bF_buf0));
BUFX4 BUFX4_1214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4));
BUFX4 BUFX4_1215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3));
BUFX4 BUFX4_1216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2));
BUFX4 BUFX4_1217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1));
BUFX4 BUFX4_1218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0));
BUFX4 BUFX4_1219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf4));
BUFX4 BUFX4_122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1));
BUFX4 BUFX4_1220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf3));
BUFX4 BUFX4_1221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf2));
BUFX4 BUFX4_1222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf1));
BUFX4 BUFX4_1223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7613__bF_buf0));
BUFX4 BUFX4_1224 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf4_));
BUFX4 BUFX4_1225 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf3_));
BUFX4 BUFX4_1226 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf2_));
BUFX4 BUFX4_1227 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf1_));
BUFX4 BUFX4_1228 ( .A(alu_b_i_0_), .Y(alu_b_i_0_bF_buf0_));
BUFX4 BUFX4_1229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf4));
BUFX4 BUFX4_123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf0));
BUFX4 BUFX4_1230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf3));
BUFX4 BUFX4_1231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf2));
BUFX4 BUFX4_1232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf1));
BUFX4 BUFX4_1233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7592__bF_buf0));
BUFX4 BUFX4_1234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf4));
BUFX4 BUFX4_1235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf3));
BUFX4 BUFX4_1236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf2));
BUFX4 BUFX4_1237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf1));
BUFX4 BUFX4_1238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7648__bF_buf0));
BUFX4 BUFX4_1239 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_));
BUFX4 BUFX4_124 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_));
BUFX4 BUFX4_1240 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_));
BUFX4 BUFX4_1241 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_));
BUFX4 BUFX4_1242 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_));
BUFX4 BUFX4_1243 ( .A(_abc_44694_new_n2779_), .Y(_abc_44694_new_n2779__bF_buf4));
BUFX4 BUFX4_1244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf4));
BUFX4 BUFX4_1245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf3));
BUFX4 BUFX4_1246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf2));
BUFX4 BUFX4_1247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf1));
BUFX4 BUFX4_1248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5617_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5617__bF_buf0));
BUFX4 BUFX4_1249 ( .A(_abc_44694_new_n1019_), .Y(_abc_44694_new_n1019__bF_buf4));
BUFX4 BUFX4_125 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_));
BUFX4 BUFX4_1250 ( .A(_abc_44694_new_n1019_), .Y(_abc_44694_new_n1019__bF_buf3));
BUFX4 BUFX4_1251 ( .A(_abc_44694_new_n1019_), .Y(_abc_44694_new_n1019__bF_buf2));
BUFX4 BUFX4_1252 ( .A(_abc_44694_new_n1019_), .Y(_abc_44694_new_n1019__bF_buf1));
BUFX4 BUFX4_1253 ( .A(_abc_44694_new_n1019_), .Y(_abc_44694_new_n1019__bF_buf0));
BUFX4 BUFX4_1254 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_));
BUFX4 BUFX4_1255 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_));
BUFX4 BUFX4_1256 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_));
BUFX4 BUFX4_1257 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_));
BUFX4 BUFX4_1258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf4));
BUFX4 BUFX4_1259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf3));
BUFX4 BUFX4_126 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_));
BUFX4 BUFX4_1260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf2));
BUFX4 BUFX4_1261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf1));
BUFX4 BUFX4_1262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7610__bF_buf0));
BUFX4 BUFX4_1263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4));
BUFX4 BUFX4_1264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3));
BUFX4 BUFX4_1265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2));
BUFX4 BUFX4_1266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1));
BUFX4 BUFX4_1267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0));
BUFX4 BUFX4_1268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf4));
BUFX4 BUFX4_1269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf3));
BUFX4 BUFX4_127 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_));
BUFX4 BUFX4_1270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf2));
BUFX4 BUFX4_1271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf1));
BUFX4 BUFX4_1272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5558__bF_buf0));
BUFX4 BUFX4_1273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf4));
BUFX4 BUFX4_1274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf3));
BUFX4 BUFX4_1275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf2));
BUFX4 BUFX4_1276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf1));
BUFX4 BUFX4_1277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5596_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5596__bF_buf0));
BUFX4 BUFX4_1278 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf7));
BUFX4 BUFX4_1279 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf6));
BUFX4 BUFX4_128 ( .A(alu__abc_42281_new_n950_), .Y(alu__abc_42281_new_n950__bF_buf4));
BUFX4 BUFX4_1280 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf5));
BUFX4 BUFX4_1281 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf4));
BUFX4 BUFX4_1282 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf3));
BUFX4 BUFX4_1283 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf2));
BUFX4 BUFX4_1284 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf1));
BUFX4 BUFX4_1285 ( .A(_abc_44694_new_n1210_), .Y(_abc_44694_new_n1210__bF_buf0));
BUFX4 BUFX4_129 ( .A(alu__abc_42281_new_n950_), .Y(alu__abc_42281_new_n950__bF_buf3));
BUFX4 BUFX4_13 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf1));
BUFX4 BUFX4_130 ( .A(alu__abc_42281_new_n950_), .Y(alu__abc_42281_new_n950__bF_buf2));
BUFX4 BUFX4_131 ( .A(alu__abc_42281_new_n950_), .Y(alu__abc_42281_new_n950__bF_buf1));
BUFX4 BUFX4_132 ( .A(alu__abc_42281_new_n950_), .Y(alu__abc_42281_new_n950__bF_buf0));
BUFX4 BUFX4_133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf4));
BUFX4 BUFX4_134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf3));
BUFX4 BUFX4_135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf2));
BUFX4 BUFX4_136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf1));
BUFX4 BUFX4_137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5640__bF_buf0));
BUFX4 BUFX4_138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf4));
BUFX4 BUFX4_139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf3));
BUFX4 BUFX4_14 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf0));
BUFX4 BUFX4_140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf2));
BUFX4 BUFX4_141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf1));
BUFX4 BUFX4_142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5543__bF_buf0));
BUFX4 BUFX4_143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4));
BUFX4 BUFX4_144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3));
BUFX4 BUFX4_145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2));
BUFX4 BUFX4_146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1));
BUFX4 BUFX4_147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0));
BUFX4 BUFX4_148 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf114));
BUFX4 BUFX4_149 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf113));
BUFX4 BUFX4_15 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8));
BUFX4 BUFX4_150 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf112));
BUFX4 BUFX4_151 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf111));
BUFX4 BUFX4_152 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf110));
BUFX4 BUFX4_153 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf109));
BUFX4 BUFX4_154 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf108));
BUFX4 BUFX4_155 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf107));
BUFX4 BUFX4_156 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf106));
BUFX4 BUFX4_157 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf105));
BUFX4 BUFX4_158 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf104));
BUFX4 BUFX4_159 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf103));
BUFX4 BUFX4_16 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7));
BUFX4 BUFX4_160 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf102));
BUFX4 BUFX4_161 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf101));
BUFX4 BUFX4_162 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf100));
BUFX4 BUFX4_163 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf99));
BUFX4 BUFX4_164 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf98));
BUFX4 BUFX4_165 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf97));
BUFX4 BUFX4_166 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf96));
BUFX4 BUFX4_167 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf95));
BUFX4 BUFX4_168 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf94));
BUFX4 BUFX4_169 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf93));
BUFX4 BUFX4_17 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6));
BUFX4 BUFX4_170 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf92));
BUFX4 BUFX4_171 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf91));
BUFX4 BUFX4_172 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf90));
BUFX4 BUFX4_173 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf89));
BUFX4 BUFX4_174 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf88));
BUFX4 BUFX4_175 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf87));
BUFX4 BUFX4_176 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf86));
BUFX4 BUFX4_177 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf85));
BUFX4 BUFX4_178 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf84));
BUFX4 BUFX4_179 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf83));
BUFX4 BUFX4_18 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5));
BUFX4 BUFX4_180 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf82));
BUFX4 BUFX4_181 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf81));
BUFX4 BUFX4_182 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf80));
BUFX4 BUFX4_183 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf79));
BUFX4 BUFX4_184 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf78));
BUFX4 BUFX4_185 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf77));
BUFX4 BUFX4_186 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf76));
BUFX4 BUFX4_187 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf75));
BUFX4 BUFX4_188 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf74));
BUFX4 BUFX4_189 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf73));
BUFX4 BUFX4_19 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4));
BUFX4 BUFX4_190 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf72));
BUFX4 BUFX4_191 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf71));
BUFX4 BUFX4_192 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf70));
BUFX4 BUFX4_193 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf69));
BUFX4 BUFX4_194 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf68));
BUFX4 BUFX4_195 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf67));
BUFX4 BUFX4_196 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf66));
BUFX4 BUFX4_197 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf65));
BUFX4 BUFX4_198 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf64));
BUFX4 BUFX4_199 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf63));
BUFX4 BUFX4_2 ( .A(clk_i), .Y(clk_i_hier0_bF_buf8));
BUFX4 BUFX4_20 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3));
BUFX4 BUFX4_200 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf62));
BUFX4 BUFX4_201 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf61));
BUFX4 BUFX4_202 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf60));
BUFX4 BUFX4_203 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf59));
BUFX4 BUFX4_204 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf58));
BUFX4 BUFX4_205 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf57));
BUFX4 BUFX4_206 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf56));
BUFX4 BUFX4_207 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf55));
BUFX4 BUFX4_208 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf54));
BUFX4 BUFX4_209 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf53));
BUFX4 BUFX4_21 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2));
BUFX4 BUFX4_210 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf52));
BUFX4 BUFX4_211 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf51));
BUFX4 BUFX4_212 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf50));
BUFX4 BUFX4_213 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf49));
BUFX4 BUFX4_214 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf48));
BUFX4 BUFX4_215 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf47));
BUFX4 BUFX4_216 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf46));
BUFX4 BUFX4_217 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf45));
BUFX4 BUFX4_218 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf44));
BUFX4 BUFX4_219 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf43));
BUFX4 BUFX4_22 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1));
BUFX4 BUFX4_220 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf42));
BUFX4 BUFX4_221 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf41));
BUFX4 BUFX4_222 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf40));
BUFX4 BUFX4_223 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf39));
BUFX4 BUFX4_224 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf38));
BUFX4 BUFX4_225 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf37));
BUFX4 BUFX4_226 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf36));
BUFX4 BUFX4_227 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf35));
BUFX4 BUFX4_228 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf34));
BUFX4 BUFX4_229 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf33));
BUFX4 BUFX4_23 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0));
BUFX4 BUFX4_230 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf32));
BUFX4 BUFX4_231 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf31));
BUFX4 BUFX4_232 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf30));
BUFX4 BUFX4_233 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf29));
BUFX4 BUFX4_234 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf28));
BUFX4 BUFX4_235 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf27));
BUFX4 BUFX4_236 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf26));
BUFX4 BUFX4_237 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf25));
BUFX4 BUFX4_238 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf24));
BUFX4 BUFX4_239 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf23));
BUFX4 BUFX4_24 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf4));
BUFX4 BUFX4_240 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf22));
BUFX4 BUFX4_241 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf21));
BUFX4 BUFX4_242 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf20));
BUFX4 BUFX4_243 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf19));
BUFX4 BUFX4_244 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf18));
BUFX4 BUFX4_245 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf17));
BUFX4 BUFX4_246 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf16));
BUFX4 BUFX4_247 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf15));
BUFX4 BUFX4_248 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf14));
BUFX4 BUFX4_249 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf13));
BUFX4 BUFX4_25 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf3));
BUFX4 BUFX4_250 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf12));
BUFX4 BUFX4_251 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf11));
BUFX4 BUFX4_252 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf10));
BUFX4 BUFX4_253 ( .A(clk_i_hier0_bF_buf4), .Y(clk_i_bF_buf9));
BUFX4 BUFX4_254 ( .A(clk_i_hier0_bF_buf3), .Y(clk_i_bF_buf8));
BUFX4 BUFX4_255 ( .A(clk_i_hier0_bF_buf2), .Y(clk_i_bF_buf7));
BUFX4 BUFX4_256 ( .A(clk_i_hier0_bF_buf1), .Y(clk_i_bF_buf6));
BUFX4 BUFX4_257 ( .A(clk_i_hier0_bF_buf0), .Y(clk_i_bF_buf5));
BUFX4 BUFX4_258 ( .A(clk_i_hier0_bF_buf9), .Y(clk_i_bF_buf4));
BUFX4 BUFX4_259 ( .A(clk_i_hier0_bF_buf8), .Y(clk_i_bF_buf3));
BUFX4 BUFX4_26 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf2));
BUFX4 BUFX4_260 ( .A(clk_i_hier0_bF_buf7), .Y(clk_i_bF_buf2));
BUFX4 BUFX4_261 ( .A(clk_i_hier0_bF_buf6), .Y(clk_i_bF_buf1));
BUFX4 BUFX4_262 ( .A(clk_i_hier0_bF_buf5), .Y(clk_i_bF_buf0));
BUFX4 BUFX4_263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4));
BUFX4 BUFX4_264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3));
BUFX4 BUFX4_265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2));
BUFX4 BUFX4_266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1));
BUFX4 BUFX4_267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0));
BUFX4 BUFX4_268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4));
BUFX4 BUFX4_269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3));
BUFX4 BUFX4_27 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf1));
BUFX4 BUFX4_270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2));
BUFX4 BUFX4_271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1));
BUFX4 BUFX4_272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0));
BUFX4 BUFX4_273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf4));
BUFX4 BUFX4_274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf3));
BUFX4 BUFX4_275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf2));
BUFX4 BUFX4_276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf1));
BUFX4 BUFX4_277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7627_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7627__bF_buf0));
BUFX4 BUFX4_278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf4));
BUFX4 BUFX4_279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf3));
BUFX4 BUFX4_28 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7645_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7645__bF_buf0));
BUFX4 BUFX4_280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf2));
BUFX4 BUFX4_281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf1));
BUFX4 BUFX4_282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7568__bF_buf0));
BUFX4 BUFX4_283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4));
BUFX4 BUFX4_284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3));
BUFX4 BUFX4_285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2));
BUFX4 BUFX4_286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1));
BUFX4 BUFX4_287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0));
BUFX4 BUFX4_288 ( .A(state_q_1_), .Y(state_q_1_bF_buf4_));
BUFX4 BUFX4_289 ( .A(state_q_1_), .Y(state_q_1_bF_buf3_));
BUFX4 BUFX4_29 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_));
BUFX4 BUFX4_290 ( .A(state_q_1_), .Y(state_q_1_bF_buf2_));
BUFX4 BUFX4_291 ( .A(state_q_1_), .Y(state_q_1_bF_buf1_));
BUFX4 BUFX4_292 ( .A(state_q_1_), .Y(state_q_1_bF_buf0_));
BUFX4 BUFX4_293 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98));
BUFX4 BUFX4_294 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97));
BUFX4 BUFX4_295 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96));
BUFX4 BUFX4_296 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95));
BUFX4 BUFX4_297 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94));
BUFX4 BUFX4_298 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93));
BUFX4 BUFX4_299 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92));
BUFX4 BUFX4_3 ( .A(clk_i), .Y(clk_i_hier0_bF_buf7));
BUFX4 BUFX4_30 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_));
BUFX4 BUFX4_300 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91));
BUFX4 BUFX4_301 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90));
BUFX4 BUFX4_302 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89));
BUFX4 BUFX4_303 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88));
BUFX4 BUFX4_304 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87));
BUFX4 BUFX4_305 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86));
BUFX4 BUFX4_306 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85));
BUFX4 BUFX4_307 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84));
BUFX4 BUFX4_308 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83));
BUFX4 BUFX4_309 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82));
BUFX4 BUFX4_31 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_));
BUFX4 BUFX4_310 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81));
BUFX4 BUFX4_311 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80));
BUFX4 BUFX4_312 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79));
BUFX4 BUFX4_313 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78));
BUFX4 BUFX4_314 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77));
BUFX4 BUFX4_315 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76));
BUFX4 BUFX4_316 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75));
BUFX4 BUFX4_317 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74));
BUFX4 BUFX4_318 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73));
BUFX4 BUFX4_319 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72));
BUFX4 BUFX4_32 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_));
BUFX4 BUFX4_320 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71));
BUFX4 BUFX4_321 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70));
BUFX4 BUFX4_322 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69));
BUFX4 BUFX4_323 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68));
BUFX4 BUFX4_324 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67));
BUFX4 BUFX4_325 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66));
BUFX4 BUFX4_326 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65));
BUFX4 BUFX4_327 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64));
BUFX4 BUFX4_328 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63));
BUFX4 BUFX4_329 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62));
BUFX4 BUFX4_33 ( .A(_abc_44694_new_n1207_), .Y(_abc_44694_new_n1207__bF_buf5));
BUFX4 BUFX4_330 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61));
BUFX4 BUFX4_331 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60));
BUFX4 BUFX4_332 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59));
BUFX4 BUFX4_333 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58));
BUFX4 BUFX4_334 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57));
BUFX4 BUFX4_335 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56));
BUFX4 BUFX4_336 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55));
BUFX4 BUFX4_337 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54));
BUFX4 BUFX4_338 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53));
BUFX4 BUFX4_339 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52));
BUFX4 BUFX4_34 ( .A(_abc_44694_new_n1207_), .Y(_abc_44694_new_n1207__bF_buf4));
BUFX4 BUFX4_340 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51));
BUFX4 BUFX4_341 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50));
BUFX4 BUFX4_342 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49));
BUFX4 BUFX4_343 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48));
BUFX4 BUFX4_344 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47));
BUFX4 BUFX4_345 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46));
BUFX4 BUFX4_346 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45));
BUFX4 BUFX4_347 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44));
BUFX4 BUFX4_348 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43));
BUFX4 BUFX4_349 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42));
BUFX4 BUFX4_35 ( .A(_abc_44694_new_n1207_), .Y(_abc_44694_new_n1207__bF_buf3));
BUFX4 BUFX4_350 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41));
BUFX4 BUFX4_351 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40));
BUFX4 BUFX4_352 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39));
BUFX4 BUFX4_353 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38));
BUFX4 BUFX4_354 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37));
BUFX4 BUFX4_355 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36));
BUFX4 BUFX4_356 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35));
BUFX4 BUFX4_357 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34));
BUFX4 BUFX4_358 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33));
BUFX4 BUFX4_359 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32));
BUFX4 BUFX4_36 ( .A(_abc_44694_new_n1207_), .Y(_abc_44694_new_n1207__bF_buf2));
BUFX4 BUFX4_360 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31));
BUFX4 BUFX4_361 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30));
BUFX4 BUFX4_362 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29));
BUFX4 BUFX4_363 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28));
BUFX4 BUFX4_364 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27));
BUFX4 BUFX4_365 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26));
BUFX4 BUFX4_366 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25));
BUFX4 BUFX4_367 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24));
BUFX4 BUFX4_368 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23));
BUFX4 BUFX4_369 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22));
BUFX4 BUFX4_37 ( .A(_abc_44694_new_n1207_), .Y(_abc_44694_new_n1207__bF_buf1));
BUFX4 BUFX4_370 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21));
BUFX4 BUFX4_371 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20));
BUFX4 BUFX4_372 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19));
BUFX4 BUFX4_373 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18));
BUFX4 BUFX4_374 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17));
BUFX4 BUFX4_375 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16));
BUFX4 BUFX4_376 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15));
BUFX4 BUFX4_377 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14));
BUFX4 BUFX4_378 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13));
BUFX4 BUFX4_379 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12));
BUFX4 BUFX4_38 ( .A(_abc_44694_new_n1207_), .Y(_abc_44694_new_n1207__bF_buf0));
BUFX4 BUFX4_380 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11));
BUFX4 BUFX4_381 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10));
BUFX4 BUFX4_382 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9));
BUFX4 BUFX4_383 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf8), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8));
BUFX4 BUFX4_384 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf7), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7));
BUFX4 BUFX4_385 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf6), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6));
BUFX4 BUFX4_386 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf5), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5));
BUFX4 BUFX4_387 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf4), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4));
BUFX4 BUFX4_388 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3));
BUFX4 BUFX4_389 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf2), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2));
BUFX4 BUFX4_39 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_));
BUFX4 BUFX4_390 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf1), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1));
BUFX4 BUFX4_391 ( .A(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_hier0_bF_buf0), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0));
BUFX4 BUFX4_392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4));
BUFX4 BUFX4_393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3));
BUFX4 BUFX4_394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2));
BUFX4 BUFX4_395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1));
BUFX4 BUFX4_396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0));
BUFX4 BUFX4_397 ( .A(alu__abc_42281_new_n941_), .Y(alu__abc_42281_new_n941__bF_buf4));
BUFX4 BUFX4_398 ( .A(alu__abc_42281_new_n941_), .Y(alu__abc_42281_new_n941__bF_buf3));
BUFX4 BUFX4_399 ( .A(alu__abc_42281_new_n941_), .Y(alu__abc_42281_new_n941__bF_buf2));
BUFX4 BUFX4_4 ( .A(clk_i), .Y(clk_i_hier0_bF_buf6));
BUFX4 BUFX4_40 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_));
BUFX4 BUFX4_400 ( .A(alu__abc_42281_new_n941_), .Y(alu__abc_42281_new_n941__bF_buf1));
BUFX4 BUFX4_401 ( .A(alu__abc_42281_new_n941_), .Y(alu__abc_42281_new_n941__bF_buf0));
BUFX4 BUFX4_402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf4));
BUFX4 BUFX4_403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf3));
BUFX4 BUFX4_404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf2));
BUFX4 BUFX4_405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf1));
BUFX4 BUFX4_406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7659__bF_buf0));
BUFX4 BUFX4_407 ( .A(alu__abc_42281_new_n271_), .Y(alu__abc_42281_new_n271__bF_buf4));
BUFX4 BUFX4_408 ( .A(alu__abc_42281_new_n271_), .Y(alu__abc_42281_new_n271__bF_buf3));
BUFX4 BUFX4_409 ( .A(alu__abc_42281_new_n271_), .Y(alu__abc_42281_new_n271__bF_buf2));
BUFX4 BUFX4_41 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_));
BUFX4 BUFX4_410 ( .A(alu__abc_42281_new_n271_), .Y(alu__abc_42281_new_n271__bF_buf1));
BUFX4 BUFX4_411 ( .A(alu__abc_42281_new_n271_), .Y(alu__abc_42281_new_n271__bF_buf0));
BUFX4 BUFX4_412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4));
BUFX4 BUFX4_413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3));
BUFX4 BUFX4_414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2));
BUFX4 BUFX4_415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1));
BUFX4 BUFX4_416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0));
BUFX4 BUFX4_417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7));
BUFX4 BUFX4_418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf6));
BUFX4 BUFX4_419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5));
BUFX4 BUFX4_42 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_));
BUFX4 BUFX4_420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf4));
BUFX4 BUFX4_421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3));
BUFX4 BUFX4_422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf2));
BUFX4 BUFX4_423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1));
BUFX4 BUFX4_424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf0));
BUFX4 BUFX4_425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf4));
BUFX4 BUFX4_426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf3));
BUFX4 BUFX4_427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf2));
BUFX4 BUFX4_428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf1));
BUFX4 BUFX4_429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5572_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5572__bF_buf0));
BUFX4 BUFX4_43 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf4));
BUFX4 BUFX4_430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf4));
BUFX4 BUFX4_431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf3));
BUFX4 BUFX4_432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf2));
BUFX4 BUFX4_433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf1));
BUFX4 BUFX4_434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5628__bF_buf0));
BUFX4 BUFX4_435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf4));
BUFX4 BUFX4_436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf3));
BUFX4 BUFX4_437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf2));
BUFX4 BUFX4_438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf1));
BUFX4 BUFX4_439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7621__bF_buf0));
BUFX4 BUFX4_44 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf3));
BUFX4 BUFX4_440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf4));
BUFX4 BUFX4_441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf3));
BUFX4 BUFX4_442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf2));
BUFX4 BUFX4_443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf1));
BUFX4 BUFX4_444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7656_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7656__bF_buf0));
BUFX4 BUFX4_445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4));
BUFX4 BUFX4_446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3));
BUFX4 BUFX4_447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2));
BUFX4 BUFX4_448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1));
BUFX4 BUFX4_449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0));
BUFX4 BUFX4_45 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf2));
BUFX4 BUFX4_450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7));
BUFX4 BUFX4_451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf6));
BUFX4 BUFX4_452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5));
BUFX4 BUFX4_453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf4));
BUFX4 BUFX4_454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3));
BUFX4 BUFX4_455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf2));
BUFX4 BUFX4_456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1));
BUFX4 BUFX4_457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf0));
BUFX4 BUFX4_458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4));
BUFX4 BUFX4_459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3));
BUFX4 BUFX4_46 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf1));
BUFX4 BUFX4_460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2));
BUFX4 BUFX4_461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1));
BUFX4 BUFX4_462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0));
BUFX4 BUFX4_463 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_));
BUFX4 BUFX4_464 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_));
BUFX4 BUFX4_465 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_));
BUFX4 BUFX4_466 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_));
BUFX4 BUFX4_467 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf6_));
BUFX4 BUFX4_468 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf5_));
BUFX4 BUFX4_469 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf4_));
BUFX4 BUFX4_47 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5649_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5649__bF_buf0));
BUFX4 BUFX4_470 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf3_));
BUFX4 BUFX4_471 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf2_));
BUFX4 BUFX4_472 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf1_));
BUFX4 BUFX4_473 ( .A(alu_b_i_2_), .Y(alu_b_i_2_bF_buf0_));
BUFX4 BUFX4_474 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_));
BUFX4 BUFX4_475 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_));
BUFX4 BUFX4_476 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_));
BUFX4 BUFX4_477 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_));
BUFX4 BUFX4_478 ( .A(_abc_44694_new_n1347_), .Y(_abc_44694_new_n1347__bF_buf4));
BUFX4 BUFX4_479 ( .A(_abc_44694_new_n1347_), .Y(_abc_44694_new_n1347__bF_buf3));
BUFX4 BUFX4_48 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4));
BUFX4 BUFX4_480 ( .A(_abc_44694_new_n1347_), .Y(_abc_44694_new_n1347__bF_buf2));
BUFX4 BUFX4_481 ( .A(_abc_44694_new_n1347_), .Y(_abc_44694_new_n1347__bF_buf1));
BUFX4 BUFX4_482 ( .A(_abc_44694_new_n1347_), .Y(_abc_44694_new_n1347__bF_buf0));
BUFX4 BUFX4_483 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15));
BUFX4 BUFX4_484 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14));
BUFX4 BUFX4_485 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13));
BUFX4 BUFX4_486 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12));
BUFX4 BUFX4_487 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11));
BUFX4 BUFX4_488 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10));
BUFX4 BUFX4_489 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9));
BUFX4 BUFX4_49 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3));
BUFX4 BUFX4_490 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8));
BUFX4 BUFX4_491 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7));
BUFX4 BUFX4_492 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6));
BUFX4 BUFX4_493 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5));
BUFX4 BUFX4_494 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4));
BUFX4 BUFX4_495 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3));
BUFX4 BUFX4_496 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2));
BUFX4 BUFX4_497 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1));
BUFX4 BUFX4_498 ( .A(_abc_44694_auto_rtlil_cc_1942_NotGate_34306), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0));
BUFX4 BUFX4_499 ( .A(_abc_44694_new_n1194_), .Y(_abc_44694_new_n1194__bF_buf4));
BUFX4 BUFX4_5 ( .A(clk_i), .Y(clk_i_hier0_bF_buf5));
BUFX4 BUFX4_50 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2));
BUFX4 BUFX4_500 ( .A(_abc_44694_new_n1194_), .Y(_abc_44694_new_n1194__bF_buf3));
BUFX4 BUFX4_501 ( .A(_abc_44694_new_n1194_), .Y(_abc_44694_new_n1194__bF_buf2));
BUFX4 BUFX4_502 ( .A(_abc_44694_new_n1194_), .Y(_abc_44694_new_n1194__bF_buf1));
BUFX4 BUFX4_503 ( .A(_abc_44694_new_n1194_), .Y(_abc_44694_new_n1194__bF_buf0));
BUFX4 BUFX4_504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf4));
BUFX4 BUFX4_505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf3));
BUFX4 BUFX4_506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf2));
BUFX4 BUFX4_507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf1));
BUFX4 BUFX4_508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7650_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7650__bF_buf0));
BUFX4 BUFX4_509 ( .A(_abc_44694_new_n2972_), .Y(_abc_44694_new_n2972__bF_buf4));
BUFX4 BUFX4_51 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1));
BUFX4 BUFX4_510 ( .A(_abc_44694_new_n2972_), .Y(_abc_44694_new_n2972__bF_buf3));
BUFX4 BUFX4_511 ( .A(_abc_44694_new_n2972_), .Y(_abc_44694_new_n2972__bF_buf2));
BUFX4 BUFX4_512 ( .A(_abc_44694_new_n2972_), .Y(_abc_44694_new_n2972__bF_buf1));
BUFX4 BUFX4_513 ( .A(_abc_44694_new_n2972_), .Y(_abc_44694_new_n2972__bF_buf0));
BUFX4 BUFX4_514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf4));
BUFX4 BUFX4_515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf3));
BUFX4 BUFX4_516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf2));
BUFX4 BUFX4_517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf1));
BUFX4 BUFX4_518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7553__bF_buf0));
BUFX4 BUFX4_519 ( .A(alu__abc_42281_new_n926_), .Y(alu__abc_42281_new_n926__bF_buf4));
BUFX4 BUFX4_52 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0));
BUFX4 BUFX4_520 ( .A(alu__abc_42281_new_n926_), .Y(alu__abc_42281_new_n926__bF_buf3));
BUFX4 BUFX4_521 ( .A(alu__abc_42281_new_n926_), .Y(alu__abc_42281_new_n926__bF_buf2));
BUFX4 BUFX4_522 ( .A(alu__abc_42281_new_n926_), .Y(alu__abc_42281_new_n926__bF_buf1));
BUFX4 BUFX4_523 ( .A(alu__abc_42281_new_n926_), .Y(alu__abc_42281_new_n926__bF_buf0));
BUFX4 BUFX4_524 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_));
BUFX4 BUFX4_525 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_));
BUFX4 BUFX4_526 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_));
BUFX4 BUFX4_527 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_));
BUFX4 BUFX4_528 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_));
BUFX4 BUFX4_529 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_));
BUFX4 BUFX4_53 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf4));
BUFX4 BUFX4_530 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_));
BUFX4 BUFX4_531 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_));
BUFX4 BUFX4_532 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf6));
BUFX4 BUFX4_533 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf5));
BUFX4 BUFX4_534 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf4));
BUFX4 BUFX4_535 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf3));
BUFX4 BUFX4_536 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf2));
BUFX4 BUFX4_537 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf1));
BUFX4 BUFX4_538 ( .A(alu__abc_42281_new_n294_), .Y(alu__abc_42281_new_n294__bF_buf0));
BUFX4 BUFX4_539 ( .A(_abc_44694_new_n3334_), .Y(_abc_44694_new_n3334__bF_buf5));
BUFX4 BUFX4_54 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf3));
BUFX4 BUFX4_540 ( .A(_abc_44694_new_n3334_), .Y(_abc_44694_new_n3334__bF_buf4));
BUFX4 BUFX4_541 ( .A(_abc_44694_new_n3334_), .Y(_abc_44694_new_n3334__bF_buf3));
BUFX4 BUFX4_542 ( .A(_abc_44694_new_n3334_), .Y(_abc_44694_new_n3334__bF_buf2));
BUFX4 BUFX4_543 ( .A(_abc_44694_new_n3334_), .Y(_abc_44694_new_n3334__bF_buf1));
BUFX4 BUFX4_544 ( .A(_abc_44694_new_n3334_), .Y(_abc_44694_new_n3334__bF_buf0));
BUFX4 BUFX4_545 ( .A(_abc_44694_new_n1400_), .Y(_abc_44694_new_n1400__bF_buf4));
BUFX4 BUFX4_546 ( .A(_abc_44694_new_n1400_), .Y(_abc_44694_new_n1400__bF_buf3));
BUFX4 BUFX4_547 ( .A(_abc_44694_new_n1400_), .Y(_abc_44694_new_n1400__bF_buf2));
BUFX4 BUFX4_548 ( .A(_abc_44694_new_n1400_), .Y(_abc_44694_new_n1400__bF_buf1));
BUFX4 BUFX4_549 ( .A(_abc_44694_new_n1400_), .Y(_abc_44694_new_n1400__bF_buf0));
BUFX4 BUFX4_55 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf2));
BUFX4 BUFX4_550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4));
BUFX4 BUFX4_551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3));
BUFX4 BUFX4_552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2));
BUFX4 BUFX4_553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1));
BUFX4 BUFX4_554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0));
BUFX4 BUFX4_555 ( .A(_abc_44694_new_n3563_), .Y(_abc_44694_new_n3563__bF_buf4));
BUFX4 BUFX4_556 ( .A(_abc_44694_new_n3563_), .Y(_abc_44694_new_n3563__bF_buf3));
BUFX4 BUFX4_557 ( .A(_abc_44694_new_n3563_), .Y(_abc_44694_new_n3563__bF_buf2));
BUFX4 BUFX4_558 ( .A(_abc_44694_new_n3563_), .Y(_abc_44694_new_n3563__bF_buf1));
BUFX4 BUFX4_559 ( .A(_abc_44694_new_n3563_), .Y(_abc_44694_new_n3563__bF_buf0));
BUFX4 BUFX4_56 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf1));
BUFX4 BUFX4_560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf4));
BUFX4 BUFX4_561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf3));
BUFX4 BUFX4_562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf2));
BUFX4 BUFX4_563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf1));
BUFX4 BUFX4_564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7606__bF_buf0));
BUFX4 BUFX4_565 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_));
BUFX4 BUFX4_566 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_));
BUFX4 BUFX4_567 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_));
BUFX4 BUFX4_568 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_));
BUFX4 BUFX4_569 ( .A(_abc_44694_new_n2546_), .Y(_abc_44694_new_n2546__bF_buf4));
BUFX4 BUFX4_57 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7604__bF_buf0));
BUFX4 BUFX4_570 ( .A(_abc_44694_new_n2546_), .Y(_abc_44694_new_n2546__bF_buf3));
BUFX4 BUFX4_571 ( .A(_abc_44694_new_n2546_), .Y(_abc_44694_new_n2546__bF_buf2));
BUFX4 BUFX4_572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf4));
BUFX4 BUFX4_573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf3));
BUFX4 BUFX4_574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf2));
BUFX4 BUFX4_575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf1));
BUFX4 BUFX4_576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5651__bF_buf0));
BUFX4 BUFX4_577 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_));
BUFX4 BUFX4_578 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_));
BUFX4 BUFX4_579 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_));
BUFX4 BUFX4_58 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4));
BUFX4 BUFX4_580 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_));
BUFX4 BUFX4_581 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_));
BUFX4 BUFX4_582 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_));
BUFX4 BUFX4_583 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_));
BUFX4 BUFX4_584 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_));
BUFX4 BUFX4_585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf4));
BUFX4 BUFX4_586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf3));
BUFX4 BUFX4_587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf2));
BUFX4 BUFX4_588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf1));
BUFX4 BUFX4_589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5554__bF_buf0));
BUFX4 BUFX4_59 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3));
BUFX4 BUFX4_590 ( .A(_abc_44694_new_n1185_), .Y(_abc_44694_new_n1185__bF_buf3));
BUFX4 BUFX4_591 ( .A(_abc_44694_new_n677_), .Y(_abc_44694_new_n677__bF_buf3));
BUFX4 BUFX4_592 ( .A(alu__abc_42281_new_n288_), .Y(alu__abc_42281_new_n288__bF_buf4));
BUFX4 BUFX4_593 ( .A(alu__abc_42281_new_n288_), .Y(alu__abc_42281_new_n288__bF_buf3));
BUFX4 BUFX4_594 ( .A(alu__abc_42281_new_n288_), .Y(alu__abc_42281_new_n288__bF_buf2));
BUFX4 BUFX4_595 ( .A(alu__abc_42281_new_n288_), .Y(alu__abc_42281_new_n288__bF_buf1));
BUFX4 BUFX4_596 ( .A(alu__abc_42281_new_n288_), .Y(alu__abc_42281_new_n288__bF_buf0));
BUFX4 BUFX4_597 ( .A(_abc_44694_new_n3519_), .Y(_abc_44694_new_n3519__bF_buf4));
BUFX4 BUFX4_598 ( .A(_abc_44694_new_n3519_), .Y(_abc_44694_new_n3519__bF_buf3));
BUFX4 BUFX4_599 ( .A(_abc_44694_new_n3519_), .Y(_abc_44694_new_n3519__bF_buf2));
BUFX4 BUFX4_6 ( .A(clk_i), .Y(clk_i_hier0_bF_buf4));
BUFX4 BUFX4_60 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2));
BUFX4 BUFX4_600 ( .A(_abc_44694_new_n3519_), .Y(_abc_44694_new_n3519__bF_buf1));
BUFX4 BUFX4_601 ( .A(_abc_44694_new_n3519_), .Y(_abc_44694_new_n3519__bF_buf0));
BUFX4 BUFX4_602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf4));
BUFX4 BUFX4_603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf3));
BUFX4 BUFX4_604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf2));
BUFX4 BUFX4_605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf1));
BUFX4 BUFX4_606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7582__bF_buf0));
BUFX4 BUFX4_607 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_));
BUFX4 BUFX4_608 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_));
BUFX4 BUFX4_609 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_));
BUFX4 BUFX4_61 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1));
BUFX4 BUFX4_610 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_));
BUFX4 BUFX4_611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf4));
BUFX4 BUFX4_612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf3));
BUFX4 BUFX4_613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf2));
BUFX4 BUFX4_614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf1));
BUFX4 BUFX4_615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7638__bF_buf0));
BUFX4 BUFX4_616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7));
BUFX4 BUFX4_617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf6));
BUFX4 BUFX4_618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5));
BUFX4 BUFX4_619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf4));
BUFX4 BUFX4_62 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0));
BUFX4 BUFX4_620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3));
BUFX4 BUFX4_621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf2));
BUFX4 BUFX4_622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1));
BUFX4 BUFX4_623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf0));
BUFX4 BUFX4_624 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_));
BUFX4 BUFX4_625 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_));
BUFX4 BUFX4_626 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_));
BUFX4 BUFX4_627 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_));
BUFX4 BUFX4_628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4));
BUFX4 BUFX4_629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3));
BUFX4 BUFX4_63 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_));
BUFX4 BUFX4_630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2));
BUFX4 BUFX4_631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1));
BUFX4 BUFX4_632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0));
BUFX4 BUFX4_633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf4));
BUFX4 BUFX4_634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf3));
BUFX4 BUFX4_635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf2));
BUFX4 BUFX4_636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf1));
BUFX4 BUFX4_637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5548_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5548__bF_buf0));
BUFX4 BUFX4_638 ( .A(_abc_44694_new_n1179_), .Y(_abc_44694_new_n1179__bF_buf3));
BUFX4 BUFX4_639 ( .A(_abc_44694_new_n1179_), .Y(_abc_44694_new_n1179__bF_buf2));
BUFX4 BUFX4_64 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_));
BUFX4 BUFX4_640 ( .A(_abc_44694_new_n1179_), .Y(_abc_44694_new_n1179__bF_buf1));
BUFX4 BUFX4_641 ( .A(_abc_44694_new_n1179_), .Y(_abc_44694_new_n1179__bF_buf0));
BUFX4 BUFX4_642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4));
BUFX4 BUFX4_643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3));
BUFX4 BUFX4_644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2));
BUFX4 BUFX4_645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1));
BUFX4 BUFX4_646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0));
BUFX4 BUFX4_647 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_));
BUFX4 BUFX4_648 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_));
BUFX4 BUFX4_649 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_));
BUFX4 BUFX4_65 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_));
BUFX4 BUFX4_650 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_));
BUFX4 BUFX4_651 ( .A(alu__abc_42281_new_n952_), .Y(alu__abc_42281_new_n952__bF_buf4));
BUFX4 BUFX4_652 ( .A(alu__abc_42281_new_n952_), .Y(alu__abc_42281_new_n952__bF_buf3));
BUFX4 BUFX4_653 ( .A(alu__abc_42281_new_n952_), .Y(alu__abc_42281_new_n952__bF_buf2));
BUFX4 BUFX4_654 ( .A(alu__abc_42281_new_n952_), .Y(alu__abc_42281_new_n952__bF_buf1));
BUFX4 BUFX4_655 ( .A(alu__abc_42281_new_n952_), .Y(alu__abc_42281_new_n952__bF_buf0));
BUFX4 BUFX4_656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4));
BUFX4 BUFX4_657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3));
BUFX4 BUFX4_658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2));
BUFX4 BUFX4_659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1));
BUFX4 BUFX4_66 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_));
BUFX4 BUFX4_660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0));
BUFX4 BUFX4_661 ( .A(_abc_44694_new_n3513_), .Y(_abc_44694_new_n3513__bF_buf4));
BUFX4 BUFX4_662 ( .A(_abc_44694_new_n3513_), .Y(_abc_44694_new_n3513__bF_buf3));
BUFX4 BUFX4_663 ( .A(_abc_44694_new_n3513_), .Y(_abc_44694_new_n3513__bF_buf2));
BUFX4 BUFX4_664 ( .A(_abc_44694_new_n3513_), .Y(_abc_44694_new_n3513__bF_buf1));
BUFX4 BUFX4_665 ( .A(_abc_44694_new_n3513_), .Y(_abc_44694_new_n3513__bF_buf0));
BUFX4 BUFX4_666 ( .A(_abc_44694_new_n668_), .Y(_abc_44694_new_n668__bF_buf4));
BUFX4 BUFX4_667 ( .A(_abc_44694_new_n668_), .Y(_abc_44694_new_n668__bF_buf3));
BUFX4 BUFX4_668 ( .A(_abc_44694_new_n668_), .Y(_abc_44694_new_n668__bF_buf2));
BUFX4 BUFX4_669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4));
BUFX4 BUFX4_67 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf4));
BUFX4 BUFX4_670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3));
BUFX4 BUFX4_671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2));
BUFX4 BUFX4_672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1));
BUFX4 BUFX4_673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0));
BUFX4 BUFX4_674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4));
BUFX4 BUFX4_675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3));
BUFX4 BUFX4_676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2));
BUFX4 BUFX4_677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1));
BUFX4 BUFX4_678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0));
BUFX4 BUFX4_679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4));
BUFX4 BUFX4_68 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf3));
BUFX4 BUFX4_680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3));
BUFX4 BUFX4_681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2));
BUFX4 BUFX4_682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1));
BUFX4 BUFX4_683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0));
BUFX4 BUFX4_684 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_));
BUFX4 BUFX4_685 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_));
BUFX4 BUFX4_686 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_));
BUFX4 BUFX4_687 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_));
BUFX4 BUFX4_688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4));
BUFX4 BUFX4_689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3));
BUFX4 BUFX4_69 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf2));
BUFX4 BUFX4_690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2));
BUFX4 BUFX4_691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1));
BUFX4 BUFX4_692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0));
BUFX4 BUFX4_693 ( .A(state_q_3_), .Y(state_q_3_bF_buf5_));
BUFX4 BUFX4_694 ( .A(state_q_3_), .Y(state_q_3_bF_buf4_));
BUFX4 BUFX4_695 ( .A(state_q_3_), .Y(state_q_3_bF_buf3_));
BUFX4 BUFX4_696 ( .A(state_q_3_), .Y(state_q_3_bF_buf2_));
BUFX4 BUFX4_697 ( .A(state_q_3_), .Y(state_q_3_bF_buf1_));
BUFX4 BUFX4_698 ( .A(state_q_3_), .Y(state_q_3_bF_buf0_));
BUFX4 BUFX4_699 ( .A(_abc_44694_new_n1399_), .Y(_abc_44694_new_n1399__bF_buf4));
BUFX4 BUFX4_7 ( .A(clk_i), .Y(clk_i_hier0_bF_buf3));
BUFX4 BUFX4_70 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf1));
BUFX4 BUFX4_700 ( .A(_abc_44694_new_n1399_), .Y(_abc_44694_new_n1399__bF_buf3));
BUFX4 BUFX4_701 ( .A(_abc_44694_new_n1399_), .Y(_abc_44694_new_n1399__bF_buf2));
BUFX4 BUFX4_702 ( .A(_abc_44694_new_n1399_), .Y(_abc_44694_new_n1399__bF_buf1));
BUFX4 BUFX4_703 ( .A(_abc_44694_new_n1399_), .Y(_abc_44694_new_n1399__bF_buf0));
BUFX4 BUFX4_704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf4));
BUFX4 BUFX4_705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf3));
BUFX4 BUFX4_706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf2));
BUFX4 BUFX4_707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf1));
BUFX4 BUFX4_708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5633_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5633__bF_buf0));
BUFX4 BUFX4_709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7));
BUFX4 BUFX4_71 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5611_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5611__bF_buf0));
BUFX4 BUFX4_710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf6));
BUFX4 BUFX4_711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5));
BUFX4 BUFX4_712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf4));
BUFX4 BUFX4_713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3));
BUFX4 BUFX4_714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf2));
BUFX4 BUFX4_715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1));
BUFX4 BUFX4_716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf0));
BUFX4 BUFX4_717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4));
BUFX4 BUFX4_718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3));
BUFX4 BUFX4_719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2));
BUFX4 BUFX4_72 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_));
BUFX4 BUFX4_720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1));
BUFX4 BUFX4_721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0));
BUFX4 BUFX4_722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4));
BUFX4 BUFX4_723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3));
BUFX4 BUFX4_724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2));
BUFX4 BUFX4_725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1));
BUFX4 BUFX4_726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0));
BUFX4 BUFX4_727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf4));
BUFX4 BUFX4_728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf3));
BUFX4 BUFX4_729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf2));
BUFX4 BUFX4_73 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_));
BUFX4 BUFX4_730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf1));
BUFX4 BUFX4_731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5574__bF_buf0));
BUFX4 BUFX4_732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7));
BUFX4 BUFX4_733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf6));
BUFX4 BUFX4_734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5));
BUFX4 BUFX4_735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf4));
BUFX4 BUFX4_736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3));
BUFX4 BUFX4_737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf2));
BUFX4 BUFX4_738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1));
BUFX4 BUFX4_739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf0));
BUFX4 BUFX4_74 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_));
BUFX4 BUFX4_740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf4));
BUFX4 BUFX4_741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf3));
BUFX4 BUFX4_742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf2));
BUFX4 BUFX4_743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf1));
BUFX4 BUFX4_744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7661_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7661__bF_buf0));
BUFX4 BUFX4_745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf4));
BUFX4 BUFX4_746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf3));
BUFX4 BUFX4_747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf2));
BUFX4 BUFX4_748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf1));
BUFX4 BUFX4_749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7564__bF_buf0));
BUFX4 BUFX4_75 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_));
BUFX4 BUFX4_750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7));
BUFX4 BUFX4_751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf6));
BUFX4 BUFX4_752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5));
BUFX4 BUFX4_753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf4));
BUFX4 BUFX4_754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3));
BUFX4 BUFX4_755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf2));
BUFX4 BUFX4_756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1));
BUFX4 BUFX4_757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf0));
BUFX4 BUFX4_758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4));
BUFX4 BUFX4_759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3));
BUFX4 BUFX4_76 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_));
BUFX4 BUFX4_760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2));
BUFX4 BUFX4_761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1));
BUFX4 BUFX4_762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0));
BUFX4 BUFX4_763 ( .A(enable_i), .Y(enable_i_bF_buf7));
BUFX4 BUFX4_764 ( .A(enable_i), .Y(enable_i_bF_buf6));
BUFX4 BUFX4_765 ( .A(enable_i), .Y(enable_i_bF_buf5));
BUFX4 BUFX4_766 ( .A(enable_i), .Y(enable_i_bF_buf4));
BUFX4 BUFX4_767 ( .A(enable_i), .Y(enable_i_bF_buf3));
BUFX4 BUFX4_768 ( .A(enable_i), .Y(enable_i_bF_buf2));
BUFX4 BUFX4_769 ( .A(enable_i), .Y(enable_i_bF_buf1));
BUFX4 BUFX4_77 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_));
BUFX4 BUFX4_770 ( .A(enable_i), .Y(enable_i_bF_buf0));
BUFX4 BUFX4_771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf4));
BUFX4 BUFX4_772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf3));
BUFX4 BUFX4_773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf2));
BUFX4 BUFX4_774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf1));
BUFX4 BUFX4_775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5568__bF_buf0));
BUFX4 BUFX4_776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7));
BUFX4 BUFX4_777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf6));
BUFX4 BUFX4_778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5));
BUFX4 BUFX4_779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf4));
BUFX4 BUFX4_78 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_));
BUFX4 BUFX4_780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3));
BUFX4 BUFX4_781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf2));
BUFX4 BUFX4_782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1));
BUFX4 BUFX4_783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf0));
BUFX4 BUFX4_784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4));
BUFX4 BUFX4_785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3));
BUFX4 BUFX4_786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2));
BUFX4 BUFX4_787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1));
BUFX4 BUFX4_788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0));
BUFX4 BUFX4_789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4));
BUFX4 BUFX4_79 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_));
BUFX4 BUFX4_790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3));
BUFX4 BUFX4_791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2));
BUFX4 BUFX4_792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1));
BUFX4 BUFX4_793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0));
BUFX4 BUFX4_794 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf5_));
BUFX4 BUFX4_795 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf4_));
BUFX4 BUFX4_796 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3_));
BUFX4 BUFX4_797 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2_));
BUFX4 BUFX4_798 ( .A(REGFILE_SIM_reg_bank_rb_i_4_), .Y(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1_));
BUFX4 BUFX4_799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf4));
BUFX4 BUFX4_8 ( .A(clk_i), .Y(clk_i_hier0_bF_buf2));
BUFX4 BUFX4_80 ( .A(_abc_44694_new_n3520_), .Y(_abc_44694_new_n3520__bF_buf4));
BUFX4 BUFX4_800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf3));
BUFX4 BUFX4_801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf2));
BUFX4 BUFX4_802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf1));
BUFX4 BUFX4_803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7558__bF_buf0));
BUFX4 BUFX4_804 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf5_));
BUFX4 BUFX4_805 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf4_));
BUFX4 BUFX4_806 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf3_));
BUFX4 BUFX4_807 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf2_));
BUFX4 BUFX4_808 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf1_));
BUFX4 BUFX4_809 ( .A(alu_b_i_4_), .Y(alu_b_i_4_bF_buf0_));
BUFX4 BUFX4_81 ( .A(_abc_44694_new_n3520_), .Y(_abc_44694_new_n3520__bF_buf3));
BUFX4 BUFX4_810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf4));
BUFX4 BUFX4_811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf3));
BUFX4 BUFX4_812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf2));
BUFX4 BUFX4_813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf1));
BUFX4 BUFX4_814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5565_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5565__bF_buf0));
BUFX4 BUFX4_815 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf6));
BUFX4 BUFX4_816 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf5));
BUFX4 BUFX4_817 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf4));
BUFX4 BUFX4_818 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf3));
BUFX4 BUFX4_819 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf2));
BUFX4 BUFX4_82 ( .A(_abc_44694_new_n3520_), .Y(_abc_44694_new_n3520__bF_buf2));
BUFX4 BUFX4_820 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf1));
BUFX4 BUFX4_821 ( .A(alu__abc_42281_new_n299_), .Y(alu__abc_42281_new_n299__bF_buf0));
BUFX4 BUFX4_822 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_));
BUFX4 BUFX4_823 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_));
BUFX4 BUFX4_824 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_));
BUFX4 BUFX4_825 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_));
BUFX4 BUFX4_826 ( .A(_abc_44694_new_n4297_), .Y(_abc_44694_new_n4297__bF_buf4));
BUFX4 BUFX4_827 ( .A(_abc_44694_new_n4297_), .Y(_abc_44694_new_n4297__bF_buf3));
BUFX4 BUFX4_828 ( .A(_abc_44694_new_n4297_), .Y(_abc_44694_new_n4297__bF_buf2));
BUFX4 BUFX4_829 ( .A(_abc_44694_new_n4297_), .Y(_abc_44694_new_n4297__bF_buf1));
BUFX4 BUFX4_83 ( .A(_abc_44694_new_n3520_), .Y(_abc_44694_new_n3520__bF_buf1));
BUFX4 BUFX4_830 ( .A(_abc_44694_new_n4297_), .Y(_abc_44694_new_n4297__bF_buf0));
BUFX4 BUFX4_831 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf7_));
BUFX4 BUFX4_832 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf6_));
BUFX4 BUFX4_833 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf5_));
BUFX4 BUFX4_834 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf4_));
BUFX4 BUFX4_835 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf3_));
BUFX4 BUFX4_836 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf2_));
BUFX4 BUFX4_837 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf1_));
BUFX4 BUFX4_838 ( .A(alu_b_i_1_), .Y(alu_b_i_1_bF_buf0_));
BUFX4 BUFX4_839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf4));
BUFX4 BUFX4_84 ( .A(_abc_44694_new_n3520_), .Y(_abc_44694_new_n3520__bF_buf0));
BUFX4 BUFX4_840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf3));
BUFX4 BUFX4_841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf2));
BUFX4 BUFX4_842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf1));
BUFX4 BUFX4_843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5621__bF_buf0));
BUFX4 BUFX4_844 ( .A(alu__abc_42281_new_n928_), .Y(alu__abc_42281_new_n928__bF_buf4));
BUFX4 BUFX4_845 ( .A(alu__abc_42281_new_n928_), .Y(alu__abc_42281_new_n928__bF_buf3));
BUFX4 BUFX4_846 ( .A(alu__abc_42281_new_n928_), .Y(alu__abc_42281_new_n928__bF_buf2));
BUFX4 BUFX4_847 ( .A(alu__abc_42281_new_n928_), .Y(alu__abc_42281_new_n928__bF_buf1));
BUFX4 BUFX4_848 ( .A(alu__abc_42281_new_n928_), .Y(alu__abc_42281_new_n928__bF_buf0));
BUFX4 BUFX4_849 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_));
BUFX4 BUFX4_85 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf4));
BUFX4 BUFX4_850 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_));
BUFX4 BUFX4_851 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_));
BUFX4 BUFX4_852 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_));
BUFX4 BUFX4_853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4));
BUFX4 BUFX4_854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3));
BUFX4 BUFX4_855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2));
BUFX4 BUFX4_856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1));
BUFX4 BUFX4_857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0));
BUFX4 BUFX4_858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7));
BUFX4 BUFX4_859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf6));
BUFX4 BUFX4_86 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf3));
BUFX4 BUFX4_860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5));
BUFX4 BUFX4_861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf4));
BUFX4 BUFX4_862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3));
BUFX4 BUFX4_863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf2));
BUFX4 BUFX4_864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1));
BUFX4 BUFX4_865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf0));
BUFX4 BUFX4_866 ( .A(_abc_44694_new_n3527_), .Y(_abc_44694_new_n3527__bF_buf4));
BUFX4 BUFX4_867 ( .A(_abc_44694_new_n3527_), .Y(_abc_44694_new_n3527__bF_buf3));
BUFX4 BUFX4_868 ( .A(_abc_44694_new_n3527_), .Y(_abc_44694_new_n3527__bF_buf2));
BUFX4 BUFX4_869 ( .A(_abc_44694_new_n3527_), .Y(_abc_44694_new_n3527__bF_buf1));
BUFX4 BUFX4_87 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf2));
BUFX4 BUFX4_870 ( .A(_abc_44694_new_n3527_), .Y(_abc_44694_new_n3527__bF_buf0));
BUFX4 BUFX4_871 ( .A(_abc_44694_new_n1114_), .Y(_abc_44694_new_n1114__bF_buf4));
BUFX4 BUFX4_872 ( .A(_abc_44694_new_n1114_), .Y(_abc_44694_new_n1114__bF_buf3));
BUFX4 BUFX4_873 ( .A(_abc_44694_new_n1114_), .Y(_abc_44694_new_n1114__bF_buf2));
BUFX4 BUFX4_874 ( .A(_abc_44694_new_n1114_), .Y(_abc_44694_new_n1114__bF_buf1));
BUFX4 BUFX4_875 ( .A(_abc_44694_new_n1114_), .Y(_abc_44694_new_n1114__bF_buf0));
BUFX4 BUFX4_876 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_));
BUFX4 BUFX4_877 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_));
BUFX4 BUFX4_878 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_));
BUFX4 BUFX4_879 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_));
BUFX4 BUFX4_88 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf1));
BUFX4 BUFX4_880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf4));
BUFX4 BUFX4_881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf3));
BUFX4 BUFX4_882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf2));
BUFX4 BUFX4_883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf1));
BUFX4 BUFX4_884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5615_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5615__bF_buf0));
BUFX4 BUFX4_885 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_));
BUFX4 BUFX4_886 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_));
BUFX4 BUFX4_887 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_));
BUFX4 BUFX4_888 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_));
BUFX4 BUFX4_889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4));
BUFX4 BUFX4_89 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5646__bF_buf0));
BUFX4 BUFX4_890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3));
BUFX4 BUFX4_891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2));
BUFX4 BUFX4_892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1));
BUFX4 BUFX4_893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0));
BUFX4 BUFX4_894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf4));
BUFX4 BUFX4_895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf3));
BUFX4 BUFX4_896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf2));
BUFX4 BUFX4_897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf1));
BUFX4 BUFX4_898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5594__bF_buf0));
BUFX4 BUFX4_899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf4));
BUFX4 BUFX4_9 ( .A(clk_i), .Y(clk_i_hier0_bF_buf1));
BUFX4 BUFX4_90 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_));
BUFX4 BUFX4_900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf3));
BUFX4 BUFX4_901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf2));
BUFX4 BUFX4_902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf1));
BUFX4 BUFX4_903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7643_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7643__bF_buf0));
BUFX4 BUFX4_904 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_));
BUFX4 BUFX4_905 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_));
BUFX4 BUFX4_906 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_));
BUFX4 BUFX4_907 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_));
BUFX4 BUFX4_908 ( .A(_abc_44694_new_n1340_), .Y(_abc_44694_new_n1340__bF_buf4));
BUFX4 BUFX4_909 ( .A(_abc_44694_new_n1340_), .Y(_abc_44694_new_n1340__bF_buf3));
BUFX4 BUFX4_91 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_));
BUFX4 BUFX4_910 ( .A(_abc_44694_new_n1340_), .Y(_abc_44694_new_n1340__bF_buf2));
BUFX4 BUFX4_911 ( .A(_abc_44694_new_n1340_), .Y(_abc_44694_new_n1340__bF_buf1));
BUFX4 BUFX4_912 ( .A(_abc_44694_new_n1340_), .Y(_abc_44694_new_n1340__bF_buf0));
BUFX4 BUFX4_913 ( .A(_abc_44694_new_n2965_), .Y(_abc_44694_new_n2965__bF_buf4));
BUFX4 BUFX4_914 ( .A(_abc_44694_new_n2965_), .Y(_abc_44694_new_n2965__bF_buf3));
BUFX4 BUFX4_915 ( .A(_abc_44694_new_n2965_), .Y(_abc_44694_new_n2965__bF_buf2));
BUFX4 BUFX4_916 ( .A(_abc_44694_new_n2965_), .Y(_abc_44694_new_n2965__bF_buf1));
BUFX4 BUFX4_917 ( .A(_abc_44694_new_n2965_), .Y(_abc_44694_new_n2965__bF_buf0));
BUFX4 BUFX4_918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf4));
BUFX4 BUFX4_919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf3));
BUFX4 BUFX4_92 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_));
BUFX4 BUFX4_920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf2));
BUFX4 BUFX4_921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf1));
BUFX4 BUFX4_922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7584_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7584__bF_buf0));
BUFX4 BUFX4_923 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_));
BUFX4 BUFX4_924 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_));
BUFX4 BUFX4_925 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_));
BUFX4 BUFX4_926 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_));
BUFX4 BUFX4_927 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_));
BUFX4 BUFX4_928 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_));
BUFX4 BUFX4_929 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_));
BUFX4 BUFX4_93 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_));
BUFX4 BUFX4_930 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_));
BUFX4 BUFX4_931 ( .A(_abc_44694_new_n1337_), .Y(_abc_44694_new_n1337__bF_buf4));
BUFX4 BUFX4_932 ( .A(_abc_44694_new_n1337_), .Y(_abc_44694_new_n1337__bF_buf3));
BUFX4 BUFX4_933 ( .A(_abc_44694_new_n1337_), .Y(_abc_44694_new_n1337__bF_buf2));
BUFX4 BUFX4_934 ( .A(_abc_44694_new_n1337_), .Y(_abc_44694_new_n1337__bF_buf1));
BUFX4 BUFX4_935 ( .A(_abc_44694_new_n1337_), .Y(_abc_44694_new_n1337__bF_buf0));
BUFX4 BUFX4_936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf4));
BUFX4 BUFX4_937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf3));
BUFX4 BUFX4_938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf2));
BUFX4 BUFX4_939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf1));
BUFX4 BUFX4_94 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf4));
BUFX4 BUFX4_940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5609_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5609__bF_buf0));
BUFX4 BUFX4_941 ( .A(_abc_44694_new_n3521_), .Y(_abc_44694_new_n3521__bF_buf4));
BUFX4 BUFX4_942 ( .A(_abc_44694_new_n3521_), .Y(_abc_44694_new_n3521__bF_buf3));
BUFX4 BUFX4_943 ( .A(_abc_44694_new_n3521_), .Y(_abc_44694_new_n3521__bF_buf2));
BUFX4 BUFX4_944 ( .A(_abc_44694_new_n3521_), .Y(_abc_44694_new_n3521__bF_buf1));
BUFX4 BUFX4_945 ( .A(_abc_44694_new_n3521_), .Y(_abc_44694_new_n3521__bF_buf0));
BUFX4 BUFX4_946 ( .A(_abc_44694_new_n1278_), .Y(_abc_44694_new_n1278__bF_buf5));
BUFX4 BUFX4_947 ( .A(_abc_44694_new_n1278_), .Y(_abc_44694_new_n1278__bF_buf4));
BUFX4 BUFX4_948 ( .A(_abc_44694_new_n1278_), .Y(_abc_44694_new_n1278__bF_buf3));
BUFX4 BUFX4_949 ( .A(_abc_44694_new_n1278_), .Y(_abc_44694_new_n1278__bF_buf2));
BUFX4 BUFX4_95 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf3));
BUFX4 BUFX4_950 ( .A(_abc_44694_new_n1278_), .Y(_abc_44694_new_n1278__bF_buf1));
BUFX4 BUFX4_951 ( .A(_abc_44694_new_n1278_), .Y(_abc_44694_new_n1278__bF_buf0));
BUFX4 BUFX4_952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4));
BUFX4 BUFX4_953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3));
BUFX4 BUFX4_954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2));
BUFX4 BUFX4_955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1));
BUFX4 BUFX4_956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0));
BUFX4 BUFX4_957 ( .A(_abc_44694_new_n1087_), .Y(_abc_44694_new_n1087__bF_buf3));
BUFX4 BUFX4_958 ( .A(_abc_44694_new_n1087_), .Y(_abc_44694_new_n1087__bF_buf2));
BUFX4 BUFX4_959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4));
BUFX4 BUFX4_96 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf2));
BUFX4 BUFX4_960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3));
BUFX4 BUFX4_961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2));
BUFX4 BUFX4_962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1));
BUFX4 BUFX4_963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0));
BUFX4 BUFX4_964 ( .A(_abc_44694_new_n3518_), .Y(_abc_44694_new_n3518__bF_buf3));
BUFX4 BUFX4_965 ( .A(_abc_44694_new_n3518_), .Y(_abc_44694_new_n3518__bF_buf2));
BUFX4 BUFX4_966 ( .A(_abc_44694_new_n3518_), .Y(_abc_44694_new_n3518__bF_buf1));
BUFX4 BUFX4_967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf4));
BUFX4 BUFX4_968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf3));
BUFX4 BUFX4_969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf2));
BUFX4 BUFX4_97 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf1));
BUFX4 BUFX4_970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf1));
BUFX4 BUFX4_971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5588__bF_buf0));
BUFX4 BUFX4_972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4));
BUFX4 BUFX4_973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3));
BUFX4 BUFX4_974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2));
BUFX4 BUFX4_975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1));
BUFX4 BUFX4_976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0));
BUFX4 BUFX4_977 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_));
BUFX4 BUFX4_978 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_));
BUFX4 BUFX4_979 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_));
BUFX4 BUFX4_98 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7636__bF_buf0));
BUFX4 BUFX4_980 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_));
BUFX4 BUFX4_981 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_));
BUFX4 BUFX4_982 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_));
BUFX4 BUFX4_983 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_));
BUFX4 BUFX4_984 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_));
BUFX4 BUFX4_985 ( .A(_abc_44694_new_n1334_), .Y(_abc_44694_new_n1334__bF_buf4));
BUFX4 BUFX4_986 ( .A(_abc_44694_new_n1334_), .Y(_abc_44694_new_n1334__bF_buf3));
BUFX4 BUFX4_987 ( .A(_abc_44694_new_n1334_), .Y(_abc_44694_new_n1334__bF_buf2));
BUFX4 BUFX4_988 ( .A(_abc_44694_new_n1334_), .Y(_abc_44694_new_n1334__bF_buf1));
BUFX4 BUFX4_989 ( .A(_abc_44694_new_n1334_), .Y(_abc_44694_new_n1334__bF_buf0));
BUFX4 BUFX4_99 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_));
BUFX4 BUFX4_990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf4));
BUFX4 BUFX4_991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf3));
BUFX4 BUFX4_992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf2));
BUFX4 BUFX4_993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf1));
BUFX4 BUFX4_994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7578__bF_buf0));
BUFX4 BUFX4_995 ( .A(_abc_44694_new_n1181_), .Y(_abc_44694_new_n1181__bF_buf3));
BUFX4 BUFX4_996 ( .A(_abc_44694_new_n1181_), .Y(_abc_44694_new_n1181__bF_buf2));
BUFX4 BUFX4_997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf4));
BUFX4 BUFX4_998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf3));
BUFX4 BUFX4_999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5644_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5644__bF_buf2));
DFFSR DFFSR_1 ( .CLK(clk_i_bF_buf114), .D(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2386), .Q(state_q_0_), .R(1'h1), .S(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3));
DFFSR DFFSR_10 ( .CLK(clk_i_bF_buf105), .D(_0pc_q_31_0__1_), .Q(next_pc_r_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk_i_bF_buf15), .D(alu_input_a_r_15_), .Q(alu_a_i_15_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_1000 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r24_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_1001 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r24_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_1002 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r24_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_1003 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r24_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_1004 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r24_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_1005 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r24_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_1006 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r24_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_1007 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r24_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_1008 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r24_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_1009 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r24_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_101 ( .CLK(clk_i_bF_buf14), .D(alu_input_a_r_16_), .Q(alu_a_i_16_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_1010 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r24_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_1011 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r24_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_1012 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r24_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_1013 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r24_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_1014 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r24_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_1015 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r24_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_1016 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r24_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_1017 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r24_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_1018 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r24_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_1019 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r24_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_102 ( .CLK(clk_i_bF_buf13), .D(alu_input_a_r_17_), .Q(alu_a_i_17_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_1020 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r24_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_1021 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r24_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_1022 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r24_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_1023 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r24_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_1024 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r24_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_1025 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r24_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_1026 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r25_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_1027 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r25_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_1028 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r25_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_1029 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r25_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_103 ( .CLK(clk_i_bF_buf12), .D(alu_input_a_r_18_), .Q(alu_a_i_18_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_1030 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r25_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_1031 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r25_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_1032 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r25_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_1033 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r25_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_1034 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r25_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_1035 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r25_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_1036 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r25_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_1037 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r25_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_1038 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r25_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_1039 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r25_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_104 ( .CLK(clk_i_bF_buf11), .D(alu_input_a_r_19_), .Q(alu_a_i_19_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_1040 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r25_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_1041 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r25_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_1042 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r25_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_1043 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r25_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_1044 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r25_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_1045 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r25_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_1046 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r25_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_1047 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r25_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_1048 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r25_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_1049 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r25_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_105 ( .CLK(clk_i_bF_buf10), .D(alu_input_a_r_20_), .Q(alu_a_i_20_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_1050 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r25_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_1051 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r25_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_1052 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r25_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_1053 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r25_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_1054 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r25_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_1055 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r25_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_1056 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r25_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_1057 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r25_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r25_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_1058 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r26_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_1059 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r26_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_106 ( .CLK(clk_i_bF_buf9), .D(alu_input_a_r_21_), .Q(alu_a_i_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_1060 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r26_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_1061 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r26_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_1062 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r26_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_1063 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r26_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_1064 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r26_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_1065 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r26_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_1066 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r26_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_1067 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r26_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_1068 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r26_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_1069 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r26_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_107 ( .CLK(clk_i_bF_buf8), .D(alu_input_a_r_22_), .Q(alu_a_i_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_1070 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r26_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_1071 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r26_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_1072 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r26_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_1073 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r26_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_1074 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r26_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_1075 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r26_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_1076 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r26_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_1077 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r26_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_1078 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r26_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_1079 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r26_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_108 ( .CLK(clk_i_bF_buf7), .D(alu_input_a_r_23_), .Q(alu_a_i_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_1080 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r26_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_1081 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r26_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_1082 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r26_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_1083 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r26_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_1084 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r26_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_1085 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r26_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_1086 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r26_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_1087 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r26_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_1088 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r26_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_1089 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r26_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r26_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_109 ( .CLK(clk_i_bF_buf6), .D(alu_input_a_r_24_), .Q(alu_a_i_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_1090 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r27_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_1091 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r27_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_1092 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r27_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_1093 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r27_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_1094 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r27_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_1095 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r27_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_1096 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r27_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_1097 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r27_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_1098 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r27_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_1099 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r27_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk_i_bF_buf104), .D(_0pc_q_31_0__2_), .Q(pc_q_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk_i_bF_buf5), .D(alu_input_a_r_25_), .Q(alu_a_i_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_1100 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r27_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_1101 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r27_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_1102 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r27_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_1103 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r27_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_1104 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r27_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_1105 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r27_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_1106 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r27_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_1107 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r27_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_1108 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r27_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_1109 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r27_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk_i_bF_buf4), .D(alu_input_a_r_26_), .Q(alu_a_i_26_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_1110 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r27_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_1111 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r27_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_1112 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r27_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_1113 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r27_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_1114 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r27_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_1115 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r27_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_1116 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r27_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_1117 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r27_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_1118 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r27_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_1119 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r27_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk_i_bF_buf3), .D(alu_input_a_r_27_), .Q(alu_a_i_27_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_1120 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r27_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_1121 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r27_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r27_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_1122 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r28_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_1123 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r28_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_1124 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r28_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_1125 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r28_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_1126 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r28_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_1127 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r28_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_1128 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r28_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_1129 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r28_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk_i_bF_buf2), .D(alu_input_a_r_28_), .Q(alu_a_i_28_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf0), .S(1'h1));
DFFSR DFFSR_1130 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r28_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_1131 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r28_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_1132 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r28_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_1133 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r28_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_1134 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r28_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_1135 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r28_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_1136 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r28_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_1137 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r28_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_1138 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r28_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_1139 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r28_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk_i_bF_buf1), .D(alu_input_a_r_29_), .Q(alu_a_i_29_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_1140 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r28_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_1141 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r28_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_1142 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r28_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_1143 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r28_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_1144 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r28_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_1145 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r28_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_1146 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r28_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_1147 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r28_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_1148 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r28_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_1149 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r28_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk_i_bF_buf0), .D(alu_input_a_r_30_), .Q(alu_a_i_30_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_1150 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r28_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_1151 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r28_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_1152 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r28_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_1153 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r28_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r28_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_1154 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r29_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_1155 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r29_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_1156 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r29_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_1157 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r29_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_1158 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r29_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_1159 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r29_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk_i_bF_buf114), .D(alu_input_a_r_31_), .Q(alu_a_i_31_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_1160 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r29_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_1161 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r29_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_1162 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r29_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_1163 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r29_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_1164 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r29_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_1165 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r29_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_1166 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r29_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_1167 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r29_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_1168 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r29_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_1169 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r29_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk_i_bF_buf113), .D(alu_input_b_r_0_), .Q(alu_b_i_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_1170 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r29_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_1171 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r29_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_1172 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r29_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_1173 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r29_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_1174 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r29_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_1175 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r29_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_1176 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r29_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_1177 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r29_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_1178 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r29_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_1179 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r29_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk_i_bF_buf112), .D(alu_input_b_r_1_), .Q(alu_b_i_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_1180 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r29_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_1181 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r29_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_1182 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r29_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_1183 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r29_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_1184 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r29_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_1185 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r29_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r29_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_1186 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r30_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_1187 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r30_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_1188 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r30_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_1189 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r30_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk_i_bF_buf111), .D(alu_input_b_r_2_), .Q(alu_b_i_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_1190 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r30_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_1191 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r30_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_1192 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r30_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_1193 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r30_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_1194 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r30_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_1195 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r30_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_1196 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r30_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_1197 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r30_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_1198 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r30_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_1199 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r30_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk_i_bF_buf103), .D(_0pc_q_31_0__3_), .Q(pc_q_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_120 ( .CLK(clk_i_bF_buf110), .D(alu_input_b_r_3_), .Q(alu_b_i_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_1200 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r30_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_1201 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r30_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_1202 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r30_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_1203 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r30_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_1204 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r30_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_1205 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r30_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_1206 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r30_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_1207 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r30_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_1208 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r30_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_1209 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r30_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk_i_bF_buf109), .D(alu_input_b_r_4_), .Q(alu_b_i_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_1210 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r30_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_1211 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r30_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_1212 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r30_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_1213 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r30_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_1214 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r30_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_1215 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r30_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_1216 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r30_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_1217 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r30_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r30_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_1218 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r31_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_1219 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r31_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk_i_bF_buf108), .D(alu_input_b_r_5_), .Q(alu_b_i_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_1220 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r31_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_1221 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r31_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_1222 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r31_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_1223 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r31_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_1224 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r31_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_1225 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r31_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_1226 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r31_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_1227 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r31_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_1228 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r31_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_1229 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r31_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk_i_bF_buf107), .D(alu_input_b_r_6_), .Q(alu_b_i_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_1230 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r31_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_1231 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r31_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_1232 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r31_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_1233 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r31_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_1234 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r31_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_1235 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r31_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_1236 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r31_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_1237 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r31_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_1238 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r31_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_1239 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r31_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk_i_bF_buf106), .D(alu_input_b_r_7_), .Q(alu_b_i_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_1240 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r31_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_1241 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r31_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_1242 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r31_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_1243 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r31_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_1244 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r31_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_1245 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r31_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_1246 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r31_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_1247 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r31_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_1248 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r31_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_1249 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r31_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r31_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk_i_bF_buf105), .D(alu_input_b_r_8_), .Q(alu_b_i_8_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk_i_bF_buf104), .D(alu_input_b_r_9_), .Q(alu_b_i_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk_i_bF_buf103), .D(alu_input_b_r_10_), .Q(alu_b_i_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk_i_bF_buf102), .D(alu_input_b_r_11_), .Q(alu_b_i_11_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk_i_bF_buf101), .D(alu_input_b_r_12_), .Q(alu_b_i_12_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk_i_bF_buf102), .D(_0pc_q_31_0__4_), .Q(pc_q_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_130 ( .CLK(clk_i_bF_buf100), .D(alu_input_b_r_13_), .Q(alu_b_i_13_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk_i_bF_buf99), .D(alu_input_b_r_14_), .Q(alu_b_i_14_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk_i_bF_buf98), .D(alu_input_b_r_15_), .Q(alu_b_i_15_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk_i_bF_buf97), .D(alu_input_b_r_16_), .Q(alu_b_i_16_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_134 ( .CLK(clk_i_bF_buf96), .D(alu_input_b_r_17_), .Q(alu_b_i_17_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk_i_bF_buf95), .D(alu_input_b_r_18_), .Q(alu_b_i_18_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk_i_bF_buf94), .D(alu_input_b_r_19_), .Q(alu_b_i_19_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk_i_bF_buf93), .D(alu_input_b_r_20_), .Q(alu_b_i_20_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk_i_bF_buf92), .D(alu_input_b_r_21_), .Q(alu_b_i_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk_i_bF_buf91), .D(alu_input_b_r_22_), .Q(alu_b_i_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_14 ( .CLK(clk_i_bF_buf101), .D(_0pc_q_31_0__5_), .Q(pc_q_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_140 ( .CLK(clk_i_bF_buf90), .D(alu_input_b_r_23_), .Q(alu_b_i_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk_i_bF_buf89), .D(alu_input_b_r_24_), .Q(alu_b_i_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk_i_bF_buf88), .D(alu_input_b_r_25_), .Q(alu_b_i_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk_i_bF_buf87), .D(alu_input_b_r_26_), .Q(alu_b_i_26_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk_i_bF_buf86), .D(alu_input_b_r_27_), .Q(alu_b_i_27_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk_i_bF_buf85), .D(alu_input_b_r_28_), .Q(alu_b_i_28_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf2), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk_i_bF_buf84), .D(alu_input_b_r_29_), .Q(alu_b_i_29_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk_i_bF_buf83), .D(alu_input_b_r_30_), .Q(alu_b_i_30_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk_i_bF_buf82), .D(alu_input_b_r_31_), .Q(alu_b_i_31_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_149 ( .CLK(clk_i_bF_buf81), .D(alu_func_r_0_), .Q(alu_op_i_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk_i_bF_buf100), .D(_0pc_q_31_0__6_), .Q(pc_q_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_150 ( .CLK(clk_i_bF_buf80), .D(alu_func_r_1_), .Q(alu_op_i_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk_i_bF_buf79), .D(alu_func_r_2_), .Q(alu_op_i_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk_i_bF_buf78), .D(alu_func_r_3_), .Q(alu_op_i_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_153 ( .CLK(clk_i_bF_buf77), .D(_0mem_addr_o_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_48711_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk_i_bF_buf76), .D(_0mem_addr_o_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_48711_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk_i_bF_buf75), .D(_0mem_addr_o_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_48711_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk_i_bF_buf74), .D(_0mem_addr_o_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_48711_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk_i_bF_buf73), .D(_0mem_addr_o_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_48711_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk_i_bF_buf72), .D(_0mem_addr_o_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_48711_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk_i_bF_buf71), .D(_0mem_addr_o_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_48711_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk_i_bF_buf99), .D(_0pc_q_31_0__7_), .Q(pc_q_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_160 ( .CLK(clk_i_bF_buf70), .D(_0mem_addr_o_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_48711_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk_i_bF_buf69), .D(_0mem_addr_o_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_48711_8_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf1), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk_i_bF_buf68), .D(_0mem_addr_o_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_48711_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk_i_bF_buf67), .D(_0mem_addr_o_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_48711_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk_i_bF_buf66), .D(_0mem_addr_o_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_48711_11_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk_i_bF_buf65), .D(_0mem_addr_o_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_48711_12_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk_i_bF_buf64), .D(_0mem_addr_o_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_48711_13_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk_i_bF_buf63), .D(_0mem_addr_o_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_48711_14_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk_i_bF_buf62), .D(_0mem_addr_o_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_48711_15_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk_i_bF_buf61), .D(_0mem_addr_o_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_48711_16_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk_i_bF_buf98), .D(_0pc_q_31_0__8_), .Q(pc_q_8_), .R(1'h1), .S(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf2));
DFFSR DFFSR_170 ( .CLK(clk_i_bF_buf60), .D(_0mem_addr_o_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_48711_17_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk_i_bF_buf59), .D(_0mem_addr_o_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_48711_18_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk_i_bF_buf58), .D(_0mem_addr_o_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_48711_19_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk_i_bF_buf57), .D(_0mem_addr_o_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_48711_20_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk_i_bF_buf56), .D(_0mem_addr_o_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_48711_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk_i_bF_buf55), .D(_0mem_addr_o_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_48711_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk_i_bF_buf54), .D(_0mem_addr_o_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_48711_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_177 ( .CLK(clk_i_bF_buf53), .D(_0mem_addr_o_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_48711_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf0), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk_i_bF_buf52), .D(_0mem_addr_o_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_48711_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk_i_bF_buf51), .D(_0mem_addr_o_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_48711_26_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk_i_bF_buf97), .D(_0pc_q_31_0__9_), .Q(pc_q_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_180 ( .CLK(clk_i_bF_buf50), .D(_0mem_addr_o_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_48711_27_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk_i_bF_buf49), .D(_0mem_addr_o_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_48711_28_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk_i_bF_buf48), .D(_0mem_addr_o_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_48711_29_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk_i_bF_buf47), .D(_0mem_addr_o_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_48711_30_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk_i_bF_buf46), .D(_0mem_addr_o_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_48711_31_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk_i_bF_buf45), .D(_0mem_dat_o_31_0__0_), .Q(_auto_iopadmap_cc_368_execute_48750_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk_i_bF_buf44), .D(_0mem_dat_o_31_0__1_), .Q(_auto_iopadmap_cc_368_execute_48750_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk_i_bF_buf43), .D(_0mem_dat_o_31_0__2_), .Q(_auto_iopadmap_cc_368_execute_48750_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk_i_bF_buf42), .D(_0mem_dat_o_31_0__3_), .Q(_auto_iopadmap_cc_368_execute_48750_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk_i_bF_buf41), .D(_0mem_dat_o_31_0__4_), .Q(_auto_iopadmap_cc_368_execute_48750_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk_i_bF_buf96), .D(_0pc_q_31_0__10_), .Q(pc_q_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_190 ( .CLK(clk_i_bF_buf40), .D(_0mem_dat_o_31_0__5_), .Q(_auto_iopadmap_cc_368_execute_48750_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk_i_bF_buf39), .D(_0mem_dat_o_31_0__6_), .Q(_auto_iopadmap_cc_368_execute_48750_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk_i_bF_buf38), .D(_0mem_dat_o_31_0__7_), .Q(_auto_iopadmap_cc_368_execute_48750_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk_i_bF_buf37), .D(_0mem_dat_o_31_0__8_), .Q(_auto_iopadmap_cc_368_execute_48750_8_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk_i_bF_buf36), .D(_0mem_dat_o_31_0__9_), .Q(_auto_iopadmap_cc_368_execute_48750_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk_i_bF_buf35), .D(_0mem_dat_o_31_0__10_), .Q(_auto_iopadmap_cc_368_execute_48750_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk_i_bF_buf34), .D(_0mem_dat_o_31_0__11_), .Q(_auto_iopadmap_cc_368_execute_48750_11_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk_i_bF_buf33), .D(_0mem_dat_o_31_0__12_), .Q(_auto_iopadmap_cc_368_execute_48750_12_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk_i_bF_buf32), .D(_0mem_dat_o_31_0__13_), .Q(_auto_iopadmap_cc_368_execute_48750_13_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk_i_bF_buf31), .D(_0mem_dat_o_31_0__14_), .Q(_auto_iopadmap_cc_368_execute_48750_14_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk_i_bF_buf113), .D(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_1_), .Q(state_q_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk_i_bF_buf95), .D(_0pc_q_31_0__11_), .Q(pc_q_11_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_200 ( .CLK(clk_i_bF_buf30), .D(_0mem_dat_o_31_0__15_), .Q(_auto_iopadmap_cc_368_execute_48750_15_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk_i_bF_buf29), .D(_0mem_dat_o_31_0__16_), .Q(_auto_iopadmap_cc_368_execute_48750_16_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk_i_bF_buf28), .D(_0mem_dat_o_31_0__17_), .Q(_auto_iopadmap_cc_368_execute_48750_17_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk_i_bF_buf27), .D(_0mem_dat_o_31_0__18_), .Q(_auto_iopadmap_cc_368_execute_48750_18_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk_i_bF_buf26), .D(_0mem_dat_o_31_0__19_), .Q(_auto_iopadmap_cc_368_execute_48750_19_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk_i_bF_buf25), .D(_0mem_dat_o_31_0__20_), .Q(_auto_iopadmap_cc_368_execute_48750_20_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk_i_bF_buf24), .D(_0mem_dat_o_31_0__21_), .Q(_auto_iopadmap_cc_368_execute_48750_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk_i_bF_buf23), .D(_0mem_dat_o_31_0__22_), .Q(_auto_iopadmap_cc_368_execute_48750_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk_i_bF_buf22), .D(_0mem_dat_o_31_0__23_), .Q(_auto_iopadmap_cc_368_execute_48750_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk_i_bF_buf21), .D(_0mem_dat_o_31_0__24_), .Q(_auto_iopadmap_cc_368_execute_48750_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf2), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk_i_bF_buf94), .D(_0pc_q_31_0__12_), .Q(pc_q_12_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_210 ( .CLK(clk_i_bF_buf20), .D(_0mem_dat_o_31_0__25_), .Q(_auto_iopadmap_cc_368_execute_48750_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk_i_bF_buf19), .D(_0mem_dat_o_31_0__26_), .Q(_auto_iopadmap_cc_368_execute_48750_26_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk_i_bF_buf18), .D(_0mem_dat_o_31_0__27_), .Q(_auto_iopadmap_cc_368_execute_48750_27_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk_i_bF_buf17), .D(_0mem_dat_o_31_0__28_), .Q(_auto_iopadmap_cc_368_execute_48750_28_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk_i_bF_buf16), .D(_0mem_dat_o_31_0__29_), .Q(_auto_iopadmap_cc_368_execute_48750_29_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk_i_bF_buf15), .D(_0mem_dat_o_31_0__30_), .Q(_auto_iopadmap_cc_368_execute_48750_30_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk_i_bF_buf14), .D(_0mem_dat_o_31_0__31_), .Q(_auto_iopadmap_cc_368_execute_48750_31_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk_i_bF_buf13), .D(_0mem_cyc_o_0_0_), .Q(_auto_iopadmap_cc_368_execute_48748), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk_i_bF_buf12), .D(_0mem_stb_o_0_0_), .Q(_auto_iopadmap_cc_368_execute_48788), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk_i_bF_buf11), .D(_0mem_we_o_0_0_), .Q(_auto_iopadmap_cc_368_execute_48790), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk_i_bF_buf93), .D(_0pc_q_31_0__13_), .Q(pc_q_13_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_220 ( .CLK(clk_i_bF_buf10), .D(_0mem_sel_o_3_0__0_), .Q(_auto_iopadmap_cc_368_execute_48783_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk_i_bF_buf9), .D(_0mem_sel_o_3_0__1_), .Q(_auto_iopadmap_cc_368_execute_48783_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk_i_bF_buf8), .D(_0mem_sel_o_3_0__2_), .Q(_auto_iopadmap_cc_368_execute_48783_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk_i_bF_buf7), .D(_0mem_sel_o_3_0__3_), .Q(_auto_iopadmap_cc_368_execute_48783_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk_i_bF_buf6), .D(_0opcode_q_31_0__0_), .Q(alu_op_r_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk_i_bF_buf5), .D(_0opcode_q_31_0__1_), .Q(alu_op_r_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf1), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk_i_bF_buf4), .D(_0opcode_q_31_0__2_), .Q(alu_op_r_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk_i_bF_buf3), .D(_0opcode_q_31_0__3_), .Q(alu_op_r_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk_i_bF_buf2), .D(_0opcode_q_31_0__4_), .Q(int32_r_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk_i_bF_buf1), .D(_0opcode_q_31_0__5_), .Q(int32_r_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk_i_bF_buf92), .D(_0pc_q_31_0__14_), .Q(pc_q_14_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_230 ( .CLK(clk_i_bF_buf0), .D(_0opcode_q_31_0__6_), .Q(alu_op_r_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk_i_bF_buf114), .D(_0opcode_q_31_0__7_), .Q(alu_op_r_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk_i_bF_buf113), .D(_0opcode_q_31_0__8_), .Q(alu_op_r_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk_i_bF_buf112), .D(_0opcode_q_31_0__9_), .Q(alu_op_r_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk_i_bF_buf111), .D(_0opcode_q_31_0__10_), .Q(int32_r_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk_i_bF_buf110), .D(_0opcode_q_31_0__11_), .Q(REGFILE_SIM_reg_bank_rb_i_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk_i_bF_buf109), .D(_0opcode_q_31_0__12_), .Q(REGFILE_SIM_reg_bank_rb_i_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk_i_bF_buf108), .D(_0opcode_q_31_0__13_), .Q(REGFILE_SIM_reg_bank_rb_i_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk_i_bF_buf107), .D(_0opcode_q_31_0__14_), .Q(REGFILE_SIM_reg_bank_rb_i_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk_i_bF_buf106), .D(_0opcode_q_31_0__15_), .Q(REGFILE_SIM_reg_bank_rb_i_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk_i_bF_buf91), .D(_0pc_q_31_0__15_), .Q(pc_q_15_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_240 ( .CLK(clk_i_bF_buf105), .D(_0opcode_q_31_0__16_), .Q(REGFILE_SIM_reg_bank_ra_i_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk_i_bF_buf104), .D(_0opcode_q_31_0__17_), .Q(REGFILE_SIM_reg_bank_ra_i_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf0), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk_i_bF_buf103), .D(_0opcode_q_31_0__18_), .Q(REGFILE_SIM_reg_bank_ra_i_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk_i_bF_buf102), .D(_0opcode_q_31_0__19_), .Q(REGFILE_SIM_reg_bank_ra_i_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk_i_bF_buf101), .D(_0opcode_q_31_0__20_), .Q(REGFILE_SIM_reg_bank_ra_i_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk_i_bF_buf100), .D(_0opcode_q_31_0__21_), .Q(opcode_q_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk_i_bF_buf99), .D(_0opcode_q_31_0__22_), .Q(opcode_q_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk_i_bF_buf98), .D(_0opcode_q_31_0__23_), .Q(opcode_q_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_248 ( .CLK(clk_i_bF_buf97), .D(_0opcode_q_31_0__24_), .Q(opcode_q_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk_i_bF_buf96), .D(_0opcode_q_31_0__25_), .Q(opcode_q_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_25 ( .CLK(clk_i_bF_buf90), .D(_0pc_q_31_0__16_), .Q(pc_q_16_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_250 ( .CLK(clk_i_bF_buf95), .D(_0opcode_q_31_0__26_), .Q(inst_r_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_251 ( .CLK(clk_i_bF_buf94), .D(_0opcode_q_31_0__27_), .Q(inst_r_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_252 ( .CLK(clk_i_bF_buf93), .D(_0opcode_q_31_0__28_), .Q(inst_r_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_253 ( .CLK(clk_i_bF_buf92), .D(_0opcode_q_31_0__29_), .Q(inst_r_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_254 ( .CLK(clk_i_bF_buf91), .D(_0opcode_q_31_0__30_), .Q(inst_r_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk_i_bF_buf90), .D(_0opcode_q_31_0__31_), .Q(inst_r_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk_i_bF_buf89), .D(_0mem_offset_q_1_0__0_), .Q(mem_offset_q_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk_i_bF_buf88), .D(_0mem_offset_q_1_0__1_), .Q(mem_offset_q_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk_i_bF_buf89), .D(_0pc_q_31_0__17_), .Q(pc_q_17_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_260 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk_i_bF_buf88), .D(_0pc_q_31_0__18_), .Q(pc_q_18_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_270 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_273 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_276 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_277 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_278 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_28 ( .CLK(clk_i_bF_buf87), .D(_0pc_q_31_0__19_), .Q(pc_q_19_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_280 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_281 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_282 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_289 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r2_fp_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk_i_bF_buf86), .D(_0pc_q_31_0__20_), .Q(pc_q_20_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_290 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r3_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r3_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r3_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r3_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r3_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r3_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r3_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r3_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r3_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r3_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_3 ( .CLK(clk_i_bF_buf112), .D(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_2_), .Q(state_q_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk_i_bF_buf85), .D(_0pc_q_31_0__21_), .Q(pc_q_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_300 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r3_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_301 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r3_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_302 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r3_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_303 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r3_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_304 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r3_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_305 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r3_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_306 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r3_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_307 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r3_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_308 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r3_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_309 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r3_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk_i_bF_buf84), .D(_0pc_q_31_0__22_), .Q(pc_q_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_310 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r3_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_311 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r3_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_312 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r3_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_313 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r3_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_314 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r3_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_315 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r3_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_316 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r3_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_317 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r3_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_318 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r3_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_319 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r3_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_32 ( .CLK(clk_i_bF_buf83), .D(_0pc_q_31_0__23_), .Q(pc_q_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_320 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r3_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_321 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r3_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r3_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_322 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r4_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_323 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r4_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_324 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r4_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_325 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r4_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_326 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r4_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_327 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r4_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_328 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r4_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_329 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r4_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_33 ( .CLK(clk_i_bF_buf82), .D(_0pc_q_31_0__24_), .Q(pc_q_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf1), .S(1'h1));
DFFSR DFFSR_330 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r4_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_331 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r4_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_332 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r4_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_333 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r4_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_334 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r4_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_335 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r4_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_336 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r4_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_337 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r4_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_338 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r4_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_339 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r4_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_34 ( .CLK(clk_i_bF_buf81), .D(_0pc_q_31_0__25_), .Q(pc_q_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_340 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r4_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_341 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r4_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_342 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r4_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_343 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r4_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_344 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r4_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_345 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r4_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_346 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r4_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_347 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r4_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_348 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r4_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_349 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r4_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_35 ( .CLK(clk_i_bF_buf80), .D(_0pc_q_31_0__26_), .Q(pc_q_26_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_350 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r4_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_351 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r4_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_352 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r4_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_353 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r4_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r4_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_354 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r5_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_355 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r5_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_356 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r5_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_357 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r5_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_358 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r5_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_359 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r5_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_36 ( .CLK(clk_i_bF_buf79), .D(_0pc_q_31_0__27_), .Q(pc_q_27_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_360 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r5_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_361 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r5_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_362 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r5_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_363 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r5_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_364 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r5_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_365 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r5_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_366 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r5_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_367 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r5_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_368 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r5_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_369 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r5_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_37 ( .CLK(clk_i_bF_buf78), .D(_0pc_q_31_0__28_), .Q(pc_q_28_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_370 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r5_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_371 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r5_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_372 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r5_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_373 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r5_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_374 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r5_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_375 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r5_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_376 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r5_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_377 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r5_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_378 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r5_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_379 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r5_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_38 ( .CLK(clk_i_bF_buf77), .D(_0pc_q_31_0__29_), .Q(pc_q_29_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_380 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r5_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_381 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r5_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_382 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r5_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_383 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r5_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_384 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r5_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_385 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r5_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r5_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_386 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r6_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_387 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r6_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_388 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r6_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_389 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r6_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_39 ( .CLK(clk_i_bF_buf76), .D(_0pc_q_31_0__30_), .Q(pc_q_30_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_390 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r6_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_391 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r6_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_392 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r6_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_393 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r6_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_394 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r6_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_395 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r6_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_396 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r6_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_397 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r6_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_398 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r6_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_399 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r6_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_4 ( .CLK(clk_i_bF_buf111), .D(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_3_), .Q(state_q_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk_i_bF_buf75), .D(_0pc_q_31_0__31_), .Q(pc_q_31_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_400 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r6_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_401 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r6_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_402 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r6_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_403 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r6_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_404 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r6_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_405 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r6_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_406 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r6_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_407 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r6_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_408 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r6_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_409 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r6_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk_i_bF_buf74), .D(_0epc_q_31_0__0_), .Q(epc_q_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_410 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r6_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_411 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r6_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_412 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r6_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_413 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r6_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_414 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r6_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_415 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r6_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_416 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r6_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_417 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r6_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r6_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_418 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r7_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_419 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r7_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk_i_bF_buf73), .D(_0epc_q_31_0__1_), .Q(epc_q_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_420 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r7_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_421 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r7_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_422 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r7_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_423 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r7_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_424 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r7_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_425 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r7_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_426 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r7_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_427 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r7_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_428 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r7_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_429 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r7_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk_i_bF_buf72), .D(_0epc_q_31_0__2_), .Q(epc_q_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_430 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r7_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_431 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r7_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_432 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r7_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_433 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r7_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_434 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r7_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_435 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r7_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_436 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r7_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_437 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r7_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_438 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r7_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_439 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r7_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk_i_bF_buf71), .D(_0epc_q_31_0__3_), .Q(epc_q_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_440 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r7_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_441 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r7_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_442 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r7_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_443 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r7_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_444 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r7_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_445 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r7_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_446 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r7_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_447 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r7_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_448 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r7_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_449 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r7_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r7_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk_i_bF_buf70), .D(_0epc_q_31_0__4_), .Q(epc_q_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_450 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r8_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_451 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r8_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_452 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r8_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_453 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r8_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_454 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r8_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_455 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r8_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_456 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r8_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_457 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r8_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_458 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r8_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_459 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r8_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk_i_bF_buf69), .D(_0epc_q_31_0__5_), .Q(epc_q_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_460 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r8_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_461 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r8_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_462 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r8_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_463 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r8_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_464 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r8_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_465 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r8_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_466 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r8_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_467 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r8_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_468 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r8_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_469 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r8_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk_i_bF_buf68), .D(_0epc_q_31_0__6_), .Q(epc_q_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_470 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r8_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_471 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r8_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_472 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r8_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_473 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r8_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_474 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r8_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_475 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r8_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_476 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r8_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_477 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r8_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_478 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r8_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_479 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r8_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk_i_bF_buf67), .D(_0epc_q_31_0__7_), .Q(epc_q_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_480 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r8_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_481 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r8_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r8_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_482 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_483 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_484 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_485 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_486 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_487 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_488 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_489 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk_i_bF_buf66), .D(_0epc_q_31_0__8_), .Q(epc_q_8_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf0), .S(1'h1));
DFFSR DFFSR_490 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_491 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_492 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_493 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_494 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_495 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_496 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_497 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_498 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_499 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_5 ( .CLK(clk_i_bF_buf110), .D(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_4_), .Q(state_q_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk_i_bF_buf65), .D(_0epc_q_31_0__9_), .Q(epc_q_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_500 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_501 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_502 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_503 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_504 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_505 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_506 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_507 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_508 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_509 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_51 ( .CLK(clk_i_bF_buf64), .D(_0epc_q_31_0__10_), .Q(epc_q_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_510 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_511 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_512 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_513 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r9_lr_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_514 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_515 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_516 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_517 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_518 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_519 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_52 ( .CLK(clk_i_bF_buf63), .D(_0epc_q_31_0__11_), .Q(epc_q_11_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_520 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_521 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_522 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_523 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_524 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_525 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_526 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_527 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_528 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_529 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_53 ( .CLK(clk_i_bF_buf62), .D(_0epc_q_31_0__12_), .Q(epc_q_12_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_530 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_531 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_532 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_533 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_534 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_535 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_536 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_537 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_538 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_539 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_54 ( .CLK(clk_i_bF_buf61), .D(_0epc_q_31_0__13_), .Q(epc_q_13_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_540 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_541 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_542 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_543 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_544 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_545 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r1_sp_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_546 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r10_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_547 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r10_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_548 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r10_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_549 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r10_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_55 ( .CLK(clk_i_bF_buf60), .D(_0epc_q_31_0__14_), .Q(epc_q_14_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_550 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r10_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_551 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r10_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_552 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r10_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_553 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r10_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_554 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r10_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_555 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r10_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_556 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r10_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_557 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r10_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_558 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r10_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_559 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r10_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_56 ( .CLK(clk_i_bF_buf59), .D(_0epc_q_31_0__15_), .Q(epc_q_15_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_560 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r10_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_561 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r10_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_562 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r10_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_563 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r10_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_564 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r10_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_565 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r10_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_566 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r10_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_567 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r10_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_568 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r10_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_569 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r10_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_57 ( .CLK(clk_i_bF_buf58), .D(_0epc_q_31_0__16_), .Q(epc_q_16_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_570 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r10_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_571 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r10_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_572 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r10_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_573 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r10_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_574 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r10_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_575 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r10_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_576 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r10_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_577 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r10_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r10_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_578 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r11_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_579 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r11_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_58 ( .CLK(clk_i_bF_buf57), .D(_0epc_q_31_0__17_), .Q(epc_q_17_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_580 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r11_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_581 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r11_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_582 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r11_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_583 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r11_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_584 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r11_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_585 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r11_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_586 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r11_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_587 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r11_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_588 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r11_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_589 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r11_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_59 ( .CLK(clk_i_bF_buf56), .D(_0epc_q_31_0__18_), .Q(epc_q_18_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_590 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r11_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_591 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r11_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_592 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r11_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_593 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r11_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_594 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r11_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_595 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r11_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_596 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r11_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_597 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r11_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_598 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r11_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_599 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r11_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_6 ( .CLK(clk_i_bF_buf109), .D(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .Q(state_q_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk_i_bF_buf55), .D(_0epc_q_31_0__19_), .Q(epc_q_19_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_600 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r11_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_601 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r11_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_602 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r11_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_603 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r11_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_604 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r11_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_605 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r11_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_606 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r11_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_607 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r11_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_608 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r11_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_609 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r11_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r11_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_61 ( .CLK(clk_i_bF_buf54), .D(_0epc_q_31_0__20_), .Q(epc_q_20_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_610 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r12_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_611 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r12_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_612 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r12_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_613 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r12_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_614 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r12_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_615 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r12_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_616 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r12_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_617 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r12_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_618 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r12_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_619 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r12_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_62 ( .CLK(clk_i_bF_buf53), .D(_0epc_q_31_0__21_), .Q(epc_q_21_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_620 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r12_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_621 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r12_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_622 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r12_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_623 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r12_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_624 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r12_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_625 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r12_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_626 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r12_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_627 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r12_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_628 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r12_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_629 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r12_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_63 ( .CLK(clk_i_bF_buf52), .D(_0epc_q_31_0__22_), .Q(epc_q_22_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_630 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r12_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_631 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r12_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_632 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r12_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_633 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r12_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_634 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r12_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_635 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r12_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_636 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r12_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_637 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r12_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_638 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r12_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_639 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r12_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_64 ( .CLK(clk_i_bF_buf51), .D(_0epc_q_31_0__23_), .Q(epc_q_23_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_640 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r12_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_641 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r12_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r12_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_642 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r13_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_643 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r13_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_644 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r13_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_645 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r13_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_646 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r13_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_647 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r13_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_648 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r13_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_649 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r13_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_65 ( .CLK(clk_i_bF_buf50), .D(_0epc_q_31_0__24_), .Q(epc_q_24_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf3), .S(1'h1));
DFFSR DFFSR_650 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r13_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_651 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r13_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_652 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r13_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_653 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r13_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_654 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r13_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_655 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r13_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_656 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r13_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_657 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r13_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_658 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r13_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_659 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r13_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_66 ( .CLK(clk_i_bF_buf49), .D(_0epc_q_31_0__25_), .Q(epc_q_25_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_660 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r13_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_661 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r13_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_662 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r13_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_663 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r13_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_664 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r13_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_665 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r13_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_666 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r13_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_667 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r13_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_668 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r13_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_669 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r13_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_67 ( .CLK(clk_i_bF_buf48), .D(_0epc_q_31_0__26_), .Q(epc_q_26_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_670 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r13_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_671 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r13_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_672 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r13_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_673 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r13_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r13_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_674 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r14_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_675 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r14_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_676 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r14_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_677 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r14_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_678 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r14_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_679 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r14_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_68 ( .CLK(clk_i_bF_buf47), .D(_0epc_q_31_0__27_), .Q(epc_q_27_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_680 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r14_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_681 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r14_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_682 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r14_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_683 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r14_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_684 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r14_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_685 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r14_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_686 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r14_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_687 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r14_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_688 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r14_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_689 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r14_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_69 ( .CLK(clk_i_bF_buf46), .D(_0epc_q_31_0__28_), .Q(epc_q_28_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_690 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r14_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_691 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r14_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_692 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r14_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_693 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r14_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_694 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r14_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_695 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r14_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_696 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r14_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_697 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r14_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_698 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r14_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_699 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r14_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_7 ( .CLK(clk_i_bF_buf108), .D(inst_trap_w), .Q(_auto_iopadmap_cc_368_execute_48707), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk_i_bF_buf45), .D(_0epc_q_31_0__29_), .Q(epc_q_29_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_700 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r14_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_701 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r14_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_702 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r14_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_703 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r14_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_704 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r14_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_705 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r14_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r14_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_706 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r15_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_707 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r15_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_708 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r15_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_709 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r15_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_71 ( .CLK(clk_i_bF_buf44), .D(_0epc_q_31_0__30_), .Q(epc_q_30_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_710 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r15_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_711 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r15_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_712 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r15_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_713 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r15_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_714 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r15_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_715 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r15_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_716 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r15_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_717 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r15_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_718 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r15_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_719 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r15_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_72 ( .CLK(clk_i_bF_buf43), .D(_0epc_q_31_0__31_), .Q(epc_q_31_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_720 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r15_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_721 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r15_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_722 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r15_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_723 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r15_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_724 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r15_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_725 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r15_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_726 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r15_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_727 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r15_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_728 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r15_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_729 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r15_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_73 ( .CLK(clk_i_bF_buf42), .D(_0sr_q_31_0__2_), .Q(sr_q_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_730 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r15_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_731 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r15_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_732 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r15_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_733 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r15_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_734 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r15_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_735 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r15_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_736 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r15_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_737 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r15_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r15_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_738 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r16_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_739 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r16_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_74 ( .CLK(clk_i_bF_buf41), .D(_0sr_q_31_0__9_), .Q(sr_q_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_740 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r16_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_741 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r16_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_742 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r16_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_743 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r16_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_744 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r16_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_745 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r16_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_746 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r16_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_747 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r16_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_748 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r16_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_749 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r16_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_75 ( .CLK(clk_i_bF_buf40), .D(_0sr_q_31_0__10_), .Q(alu_c_i), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_750 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r16_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_751 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r16_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_752 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r16_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_753 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r16_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_754 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r16_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_755 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r16_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_756 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r16_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_757 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r16_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_758 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r16_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_759 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r16_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_76 ( .CLK(clk_i_bF_buf39), .D(_0esr_q_31_0__2_), .Q(esr_q_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_760 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r16_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_761 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r16_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_762 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r16_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_763 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r16_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_764 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r16_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_765 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r16_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_766 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r16_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_767 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r16_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_768 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r16_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_769 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r16_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r16_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_77 ( .CLK(clk_i_bF_buf38), .D(_0esr_q_31_0__9_), .Q(esr_q_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_770 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r17_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_771 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r17_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_772 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r17_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_773 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r17_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_774 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r17_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_775 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r17_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_776 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r17_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_777 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r17_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_778 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r17_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_779 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r17_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk_i_bF_buf37), .D(_0esr_q_31_0__10_), .Q(esr_q_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_780 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r17_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_781 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r17_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_782 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r17_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_783 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r17_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_784 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r17_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_785 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r17_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_786 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r17_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_787 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r17_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_788 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r17_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_789 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r17_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk_i_bF_buf36), .D(_0nmi_q_0_0_), .Q(nmi_q), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_790 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r17_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_791 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r17_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_792 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r17_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_793 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r17_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_794 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r17_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_795 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r17_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_796 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r17_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_797 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r17_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_798 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r17_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_799 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r17_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk_i_bF_buf107), .D(_0fault_o_0_0_), .Q(_auto_iopadmap_cc_368_execute_48709), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk_i_bF_buf35), .D(_0ex_rd_q_4_0__0_), .Q(REGFILE_SIM_reg_bank_rd_i_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_800 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r17_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_801 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r17_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r17_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_802 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r18_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_803 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r18_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_804 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r18_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_805 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r18_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_806 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r18_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_807 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r18_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_808 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r18_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_809 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r18_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk_i_bF_buf34), .D(_0ex_rd_q_4_0__1_), .Q(REGFILE_SIM_reg_bank_rd_i_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf2), .S(1'h1));
DFFSR DFFSR_810 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r18_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_811 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r18_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_812 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r18_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_813 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r18_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_814 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r18_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_815 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r18_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_816 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r18_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_817 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r18_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_818 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r18_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_819 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r18_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_82 ( .CLK(clk_i_bF_buf33), .D(_0ex_rd_q_4_0__2_), .Q(REGFILE_SIM_reg_bank_rd_i_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_820 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r18_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_821 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r18_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_822 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r18_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_823 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r18_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_824 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r18_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_825 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r18_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_826 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r18_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_827 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r18_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_828 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r18_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_829 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r18_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk_i_bF_buf32), .D(_0ex_rd_q_4_0__3_), .Q(REGFILE_SIM_reg_bank_rd_i_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_830 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r18_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_831 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r18_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_832 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r18_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_833 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r18_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r18_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_834 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r19_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_835 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r19_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_836 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r19_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_837 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r19_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_838 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r19_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_839 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r19_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk_i_bF_buf31), .D(_0ex_rd_q_4_0__4_), .Q(REGFILE_SIM_reg_bank_rd_i_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf12), .S(1'h1));
DFFSR DFFSR_840 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r19_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_841 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r19_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_842 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r19_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_843 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r19_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_844 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r19_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_845 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r19_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_846 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r19_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_847 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r19_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_848 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r19_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_849 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r19_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk_i_bF_buf30), .D(alu_input_a_r_0_), .Q(alu_a_i_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf11), .S(1'h1));
DFFSR DFFSR_850 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r19_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_851 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r19_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_852 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r19_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_853 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r19_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_854 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r19_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_855 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r19_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_856 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r19_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_857 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r19_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_858 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r19_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_859 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r19_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk_i_bF_buf29), .D(alu_input_a_r_1_), .Q(alu_a_i_1_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf10), .S(1'h1));
DFFSR DFFSR_860 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r19_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_861 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r19_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_862 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r19_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_863 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r19_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_864 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r19_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_865 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r19_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r19_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_866 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r20_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_867 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r20_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_868 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r20_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_869 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r20_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk_i_bF_buf28), .D(alu_input_a_r_2_), .Q(alu_a_i_2_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf9), .S(1'h1));
DFFSR DFFSR_870 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r20_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_871 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r20_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_872 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r20_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_873 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r20_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_874 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r20_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_875 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r20_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_876 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r20_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_877 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r20_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_878 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r20_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_879 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r20_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk_i_bF_buf27), .D(alu_input_a_r_3_), .Q(alu_a_i_3_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf8), .S(1'h1));
DFFSR DFFSR_880 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r20_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_881 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r20_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_882 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r20_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_883 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r20_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_884 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r20_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_885 ( .CLK(clk_i_bF_buf35), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r20_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_886 ( .CLK(clk_i_bF_buf34), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r20_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_887 ( .CLK(clk_i_bF_buf33), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r20_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_888 ( .CLK(clk_i_bF_buf32), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r20_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_889 ( .CLK(clk_i_bF_buf31), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r20_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk_i_bF_buf26), .D(alu_input_a_r_4_), .Q(alu_a_i_4_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_890 ( .CLK(clk_i_bF_buf30), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r20_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_891 ( .CLK(clk_i_bF_buf29), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r20_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_892 ( .CLK(clk_i_bF_buf28), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r20_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_893 ( .CLK(clk_i_bF_buf27), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r20_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_894 ( .CLK(clk_i_bF_buf26), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r20_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_895 ( .CLK(clk_i_bF_buf25), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r20_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_896 ( .CLK(clk_i_bF_buf24), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r20_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_897 ( .CLK(clk_i_bF_buf23), .D(REGFILE_SIM_reg_bank__0reg_r20_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r20_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_898 ( .CLK(clk_i_bF_buf22), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r21_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_899 ( .CLK(clk_i_bF_buf21), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r21_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk_i_bF_buf106), .D(_0pc_q_31_0__0_), .Q(next_pc_r_0_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf7), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk_i_bF_buf25), .D(alu_input_a_r_5_), .Q(alu_a_i_5_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf6), .S(1'h1));
DFFSR DFFSR_900 ( .CLK(clk_i_bF_buf20), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r21_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
DFFSR DFFSR_901 ( .CLK(clk_i_bF_buf19), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r21_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf49), .S(1'h1));
DFFSR DFFSR_902 ( .CLK(clk_i_bF_buf18), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r21_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf48), .S(1'h1));
DFFSR DFFSR_903 ( .CLK(clk_i_bF_buf17), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r21_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf47), .S(1'h1));
DFFSR DFFSR_904 ( .CLK(clk_i_bF_buf16), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r21_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf46), .S(1'h1));
DFFSR DFFSR_905 ( .CLK(clk_i_bF_buf15), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r21_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf45), .S(1'h1));
DFFSR DFFSR_906 ( .CLK(clk_i_bF_buf14), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r21_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf44), .S(1'h1));
DFFSR DFFSR_907 ( .CLK(clk_i_bF_buf13), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r21_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf43), .S(1'h1));
DFFSR DFFSR_908 ( .CLK(clk_i_bF_buf12), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r21_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf42), .S(1'h1));
DFFSR DFFSR_909 ( .CLK(clk_i_bF_buf11), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r21_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf41), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk_i_bF_buf24), .D(alu_input_a_r_6_), .Q(alu_a_i_6_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf5), .S(1'h1));
DFFSR DFFSR_910 ( .CLK(clk_i_bF_buf10), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r21_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf40), .S(1'h1));
DFFSR DFFSR_911 ( .CLK(clk_i_bF_buf9), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r21_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf39), .S(1'h1));
DFFSR DFFSR_912 ( .CLK(clk_i_bF_buf8), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r21_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf38), .S(1'h1));
DFFSR DFFSR_913 ( .CLK(clk_i_bF_buf7), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r21_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf37), .S(1'h1));
DFFSR DFFSR_914 ( .CLK(clk_i_bF_buf6), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r21_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf36), .S(1'h1));
DFFSR DFFSR_915 ( .CLK(clk_i_bF_buf5), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r21_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf35), .S(1'h1));
DFFSR DFFSR_916 ( .CLK(clk_i_bF_buf4), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r21_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf34), .S(1'h1));
DFFSR DFFSR_917 ( .CLK(clk_i_bF_buf3), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r21_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf33), .S(1'h1));
DFFSR DFFSR_918 ( .CLK(clk_i_bF_buf2), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r21_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf32), .S(1'h1));
DFFSR DFFSR_919 ( .CLK(clk_i_bF_buf1), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r21_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf31), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk_i_bF_buf23), .D(alu_input_a_r_7_), .Q(alu_a_i_7_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf4), .S(1'h1));
DFFSR DFFSR_920 ( .CLK(clk_i_bF_buf0), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r21_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf30), .S(1'h1));
DFFSR DFFSR_921 ( .CLK(clk_i_bF_buf114), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r21_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf29), .S(1'h1));
DFFSR DFFSR_922 ( .CLK(clk_i_bF_buf113), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r21_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf28), .S(1'h1));
DFFSR DFFSR_923 ( .CLK(clk_i_bF_buf112), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r21_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf27), .S(1'h1));
DFFSR DFFSR_924 ( .CLK(clk_i_bF_buf111), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r21_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf26), .S(1'h1));
DFFSR DFFSR_925 ( .CLK(clk_i_bF_buf110), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r21_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf25), .S(1'h1));
DFFSR DFFSR_926 ( .CLK(clk_i_bF_buf109), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r21_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf24), .S(1'h1));
DFFSR DFFSR_927 ( .CLK(clk_i_bF_buf108), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r21_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf23), .S(1'h1));
DFFSR DFFSR_928 ( .CLK(clk_i_bF_buf107), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r21_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf22), .S(1'h1));
DFFSR DFFSR_929 ( .CLK(clk_i_bF_buf106), .D(REGFILE_SIM_reg_bank__0reg_r21_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r21_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf21), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk_i_bF_buf22), .D(alu_input_a_r_8_), .Q(alu_a_i_8_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf3), .S(1'h1));
DFFSR DFFSR_930 ( .CLK(clk_i_bF_buf105), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r22_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf20), .S(1'h1));
DFFSR DFFSR_931 ( .CLK(clk_i_bF_buf104), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r22_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf19), .S(1'h1));
DFFSR DFFSR_932 ( .CLK(clk_i_bF_buf103), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r22_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf18), .S(1'h1));
DFFSR DFFSR_933 ( .CLK(clk_i_bF_buf102), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r22_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf17), .S(1'h1));
DFFSR DFFSR_934 ( .CLK(clk_i_bF_buf101), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r22_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf16), .S(1'h1));
DFFSR DFFSR_935 ( .CLK(clk_i_bF_buf100), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r22_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf15), .S(1'h1));
DFFSR DFFSR_936 ( .CLK(clk_i_bF_buf99), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r22_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf14), .S(1'h1));
DFFSR DFFSR_937 ( .CLK(clk_i_bF_buf98), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r22_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf13), .S(1'h1));
DFFSR DFFSR_938 ( .CLK(clk_i_bF_buf97), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r22_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf12), .S(1'h1));
DFFSR DFFSR_939 ( .CLK(clk_i_bF_buf96), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r22_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf11), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk_i_bF_buf21), .D(alu_input_a_r_9_), .Q(alu_a_i_9_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf2), .S(1'h1));
DFFSR DFFSR_940 ( .CLK(clk_i_bF_buf95), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r22_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf10), .S(1'h1));
DFFSR DFFSR_941 ( .CLK(clk_i_bF_buf94), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r22_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf9), .S(1'h1));
DFFSR DFFSR_942 ( .CLK(clk_i_bF_buf93), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r22_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf8), .S(1'h1));
DFFSR DFFSR_943 ( .CLK(clk_i_bF_buf92), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r22_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf7), .S(1'h1));
DFFSR DFFSR_944 ( .CLK(clk_i_bF_buf91), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r22_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf6), .S(1'h1));
DFFSR DFFSR_945 ( .CLK(clk_i_bF_buf90), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r22_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf5), .S(1'h1));
DFFSR DFFSR_946 ( .CLK(clk_i_bF_buf89), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r22_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf4), .S(1'h1));
DFFSR DFFSR_947 ( .CLK(clk_i_bF_buf88), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r22_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf3), .S(1'h1));
DFFSR DFFSR_948 ( .CLK(clk_i_bF_buf87), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r22_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf2), .S(1'h1));
DFFSR DFFSR_949 ( .CLK(clk_i_bF_buf86), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r22_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf1), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk_i_bF_buf20), .D(alu_input_a_r_10_), .Q(alu_a_i_10_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf1), .S(1'h1));
DFFSR DFFSR_950 ( .CLK(clk_i_bF_buf85), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r22_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf0), .S(1'h1));
DFFSR DFFSR_951 ( .CLK(clk_i_bF_buf84), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r22_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf98), .S(1'h1));
DFFSR DFFSR_952 ( .CLK(clk_i_bF_buf83), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r22_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf97), .S(1'h1));
DFFSR DFFSR_953 ( .CLK(clk_i_bF_buf82), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r22_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf96), .S(1'h1));
DFFSR DFFSR_954 ( .CLK(clk_i_bF_buf81), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r22_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf95), .S(1'h1));
DFFSR DFFSR_955 ( .CLK(clk_i_bF_buf80), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r22_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf94), .S(1'h1));
DFFSR DFFSR_956 ( .CLK(clk_i_bF_buf79), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r22_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf93), .S(1'h1));
DFFSR DFFSR_957 ( .CLK(clk_i_bF_buf78), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r22_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf92), .S(1'h1));
DFFSR DFFSR_958 ( .CLK(clk_i_bF_buf77), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r22_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf91), .S(1'h1));
DFFSR DFFSR_959 ( .CLK(clk_i_bF_buf76), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r22_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf90), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk_i_bF_buf19), .D(alu_input_a_r_11_), .Q(alu_a_i_11_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf0), .S(1'h1));
DFFSR DFFSR_960 ( .CLK(clk_i_bF_buf75), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r22_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf89), .S(1'h1));
DFFSR DFFSR_961 ( .CLK(clk_i_bF_buf74), .D(REGFILE_SIM_reg_bank__0reg_r22_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r22_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf88), .S(1'h1));
DFFSR DFFSR_962 ( .CLK(clk_i_bF_buf73), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r23_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf87), .S(1'h1));
DFFSR DFFSR_963 ( .CLK(clk_i_bF_buf72), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r23_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf86), .S(1'h1));
DFFSR DFFSR_964 ( .CLK(clk_i_bF_buf71), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r23_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf85), .S(1'h1));
DFFSR DFFSR_965 ( .CLK(clk_i_bF_buf70), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r23_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf84), .S(1'h1));
DFFSR DFFSR_966 ( .CLK(clk_i_bF_buf69), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r23_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf83), .S(1'h1));
DFFSR DFFSR_967 ( .CLK(clk_i_bF_buf68), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r23_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf82), .S(1'h1));
DFFSR DFFSR_968 ( .CLK(clk_i_bF_buf67), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__6_), .Q(REGFILE_SIM_reg_bank_reg_r23_6_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf81), .S(1'h1));
DFFSR DFFSR_969 ( .CLK(clk_i_bF_buf66), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__7_), .Q(REGFILE_SIM_reg_bank_reg_r23_7_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf80), .S(1'h1));
DFFSR DFFSR_97 ( .CLK(clk_i_bF_buf18), .D(alu_input_a_r_12_), .Q(alu_a_i_12_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf15_bF_buf1), .S(1'h1));
DFFSR DFFSR_970 ( .CLK(clk_i_bF_buf65), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__8_), .Q(REGFILE_SIM_reg_bank_reg_r23_8_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf79), .S(1'h1));
DFFSR DFFSR_971 ( .CLK(clk_i_bF_buf64), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__9_), .Q(REGFILE_SIM_reg_bank_reg_r23_9_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf78), .S(1'h1));
DFFSR DFFSR_972 ( .CLK(clk_i_bF_buf63), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__10_), .Q(REGFILE_SIM_reg_bank_reg_r23_10_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf77), .S(1'h1));
DFFSR DFFSR_973 ( .CLK(clk_i_bF_buf62), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__11_), .Q(REGFILE_SIM_reg_bank_reg_r23_11_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf76), .S(1'h1));
DFFSR DFFSR_974 ( .CLK(clk_i_bF_buf61), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__12_), .Q(REGFILE_SIM_reg_bank_reg_r23_12_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf75), .S(1'h1));
DFFSR DFFSR_975 ( .CLK(clk_i_bF_buf60), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__13_), .Q(REGFILE_SIM_reg_bank_reg_r23_13_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf74), .S(1'h1));
DFFSR DFFSR_976 ( .CLK(clk_i_bF_buf59), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__14_), .Q(REGFILE_SIM_reg_bank_reg_r23_14_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf73), .S(1'h1));
DFFSR DFFSR_977 ( .CLK(clk_i_bF_buf58), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__15_), .Q(REGFILE_SIM_reg_bank_reg_r23_15_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf72), .S(1'h1));
DFFSR DFFSR_978 ( .CLK(clk_i_bF_buf57), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__16_), .Q(REGFILE_SIM_reg_bank_reg_r23_16_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf71), .S(1'h1));
DFFSR DFFSR_979 ( .CLK(clk_i_bF_buf56), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__17_), .Q(REGFILE_SIM_reg_bank_reg_r23_17_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf70), .S(1'h1));
DFFSR DFFSR_98 ( .CLK(clk_i_bF_buf17), .D(alu_input_a_r_13_), .Q(alu_a_i_13_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf14), .S(1'h1));
DFFSR DFFSR_980 ( .CLK(clk_i_bF_buf55), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__18_), .Q(REGFILE_SIM_reg_bank_reg_r23_18_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf69), .S(1'h1));
DFFSR DFFSR_981 ( .CLK(clk_i_bF_buf54), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__19_), .Q(REGFILE_SIM_reg_bank_reg_r23_19_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf68), .S(1'h1));
DFFSR DFFSR_982 ( .CLK(clk_i_bF_buf53), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__20_), .Q(REGFILE_SIM_reg_bank_reg_r23_20_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf67), .S(1'h1));
DFFSR DFFSR_983 ( .CLK(clk_i_bF_buf52), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__21_), .Q(REGFILE_SIM_reg_bank_reg_r23_21_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf66), .S(1'h1));
DFFSR DFFSR_984 ( .CLK(clk_i_bF_buf51), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__22_), .Q(REGFILE_SIM_reg_bank_reg_r23_22_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf65), .S(1'h1));
DFFSR DFFSR_985 ( .CLK(clk_i_bF_buf50), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__23_), .Q(REGFILE_SIM_reg_bank_reg_r23_23_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf64), .S(1'h1));
DFFSR DFFSR_986 ( .CLK(clk_i_bF_buf49), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__24_), .Q(REGFILE_SIM_reg_bank_reg_r23_24_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf63), .S(1'h1));
DFFSR DFFSR_987 ( .CLK(clk_i_bF_buf48), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__25_), .Q(REGFILE_SIM_reg_bank_reg_r23_25_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf62), .S(1'h1));
DFFSR DFFSR_988 ( .CLK(clk_i_bF_buf47), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__26_), .Q(REGFILE_SIM_reg_bank_reg_r23_26_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf61), .S(1'h1));
DFFSR DFFSR_989 ( .CLK(clk_i_bF_buf46), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__27_), .Q(REGFILE_SIM_reg_bank_reg_r23_27_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf60), .S(1'h1));
DFFSR DFFSR_99 ( .CLK(clk_i_bF_buf16), .D(alu_input_a_r_14_), .Q(alu_a_i_14_), .R(_abc_44694_auto_rtlil_cc_1942_NotGate_34306_bF_buf13), .S(1'h1));
DFFSR DFFSR_990 ( .CLK(clk_i_bF_buf45), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__28_), .Q(REGFILE_SIM_reg_bank_reg_r23_28_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf59), .S(1'h1));
DFFSR DFFSR_991 ( .CLK(clk_i_bF_buf44), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__29_), .Q(REGFILE_SIM_reg_bank_reg_r23_29_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf58), .S(1'h1));
DFFSR DFFSR_992 ( .CLK(clk_i_bF_buf43), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__30_), .Q(REGFILE_SIM_reg_bank_reg_r23_30_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf57), .S(1'h1));
DFFSR DFFSR_993 ( .CLK(clk_i_bF_buf42), .D(REGFILE_SIM_reg_bank__0reg_r23_31_0__31_), .Q(REGFILE_SIM_reg_bank_reg_r23_31_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf56), .S(1'h1));
DFFSR DFFSR_994 ( .CLK(clk_i_bF_buf41), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__0_), .Q(REGFILE_SIM_reg_bank_reg_r24_0_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf55), .S(1'h1));
DFFSR DFFSR_995 ( .CLK(clk_i_bF_buf40), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__1_), .Q(REGFILE_SIM_reg_bank_reg_r24_1_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf54), .S(1'h1));
DFFSR DFFSR_996 ( .CLK(clk_i_bF_buf39), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__2_), .Q(REGFILE_SIM_reg_bank_reg_r24_2_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf53), .S(1'h1));
DFFSR DFFSR_997 ( .CLK(clk_i_bF_buf38), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__3_), .Q(REGFILE_SIM_reg_bank_reg_r24_3_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf52), .S(1'h1));
DFFSR DFFSR_998 ( .CLK(clk_i_bF_buf37), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__4_), .Q(REGFILE_SIM_reg_bank_reg_r24_4_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf51), .S(1'h1));
DFFSR DFFSR_999 ( .CLK(clk_i_bF_buf36), .D(REGFILE_SIM_reg_bank__0reg_r24_31_0__5_), .Q(REGFILE_SIM_reg_bank_reg_r24_5_), .R(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322_bF_buf50), .S(1'h1));
INVX1 INVX1_1 ( .A(inst_r_4_), .Y(_abc_44694_new_n617_));
INVX1 INVX1_10 ( .A(_abc_44694_new_n647_), .Y(_abc_44694_new_n648_));
INVX1 INVX1_100 ( .A(_abc_44694_new_n1446_), .Y(_abc_44694_new_n1447_));
INVX1 INVX1_1000 ( .A(alu__abc_42281_new_n1483_), .Y(alu__abc_42281_new_n1484_));
INVX1 INVX1_1001 ( .A(alu__abc_42281_new_n775_), .Y(alu__abc_42281_new_n1489_));
INVX1 INVX1_1002 ( .A(alu__abc_42281_new_n1528_), .Y(alu__abc_42281_new_n1529_));
INVX1 INVX1_1003 ( .A(alu__abc_42281_new_n1534_), .Y(alu__abc_42281_new_n1535_));
INVX1 INVX1_1004 ( .A(alu__abc_42281_new_n1571_), .Y(alu__abc_42281_new_n1573_));
INVX1 INVX1_1005 ( .A(alu__abc_42281_new_n1577_), .Y(alu__abc_42281_new_n1578_));
INVX1 INVX1_1006 ( .A(alu__abc_42281_new_n1618_), .Y(alu__abc_42281_new_n1619_));
INVX1 INVX1_1007 ( .A(alu__abc_42281_new_n1623_), .Y(alu__abc_42281_new_n1624_));
INVX1 INVX1_1008 ( .A(alu__abc_42281_new_n1660_), .Y(alu__abc_42281_new_n1661_));
INVX1 INVX1_1009 ( .A(alu__abc_42281_new_n1666_), .Y(alu__abc_42281_new_n1667_));
INVX1 INVX1_101 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n1460_));
INVX1 INVX1_1010 ( .A(alu__abc_42281_new_n1707_), .Y(alu__abc_42281_new_n1708_));
INVX1 INVX1_1011 ( .A(alu__abc_42281_new_n1712_), .Y(alu__abc_42281_new_n1713_));
INVX1 INVX1_1012 ( .A(alu__abc_42281_new_n1749_), .Y(alu__abc_42281_new_n1750_));
INVX1 INVX1_1013 ( .A(alu__abc_42281_new_n806_), .Y(alu__abc_42281_new_n1757_));
INVX1 INVX1_1014 ( .A(alu__abc_42281_new_n807_), .Y(alu__abc_42281_new_n1793_));
INVX1 INVX1_1015 ( .A(alu__abc_42281_new_n1797_), .Y(alu__abc_42281_new_n1798_));
INVX1 INVX1_1016 ( .A(alu__abc_42281_new_n1836_), .Y(alu__abc_42281_new_n1837_));
INVX1 INVX1_1017 ( .A(alu__abc_42281_new_n1841_), .Y(alu__abc_42281_new_n1843_));
INVX1 INVX1_1018 ( .A(alu__abc_42281_new_n1876_), .Y(alu__abc_42281_new_n1877_));
INVX1 INVX1_1019 ( .A(alu__abc_42281_new_n1884_), .Y(alu__abc_42281_new_n1885_));
INVX1 INVX1_102 ( .A(_abc_44694_new_n1461_), .Y(_abc_44694_new_n1462_));
INVX1 INVX1_1020 ( .A(alu__abc_42281_new_n1918_), .Y(alu__abc_42281_new_n1919_));
INVX1 INVX1_1021 ( .A(alu__abc_42281_new_n1922_), .Y(alu__abc_42281_new_n1924_));
INVX1 INVX1_1022 ( .A(alu__abc_42281_new_n811_), .Y(alu__abc_42281_new_n1958_));
INVX1 INVX1_1023 ( .A(alu__abc_42281_new_n1963_), .Y(alu__abc_42281_new_n1964_));
INVX1 INVX1_1024 ( .A(alu__abc_42281_new_n1999_), .Y(alu__abc_42281_new_n2000_));
INVX1 INVX1_1025 ( .A(alu__abc_42281_new_n2003_), .Y(alu__abc_42281_new_n2004_));
INVX1 INVX1_1026 ( .A(alu__abc_42281_new_n2041_), .Y(alu__abc_42281_new_n2042_));
INVX1 INVX1_1027 ( .A(alu__abc_42281_new_n2046_), .Y(alu__abc_42281_new_n2047_));
INVX1 INVX1_1028 ( .A(alu__abc_42281_new_n2081_), .Y(alu__abc_42281_new_n2082_));
INVX1 INVX1_1029 ( .A(alu__abc_42281_new_n2085_), .Y(alu__abc_42281_new_n2086_));
INVX1 INVX1_103 ( .A(_abc_44694_new_n1468_), .Y(_abc_44694_new_n1469_));
INVX1 INVX1_1030 ( .A(alu__abc_42281_new_n2122_), .Y(alu__abc_42281_new_n2123_));
INVX1 INVX1_1031 ( .A(alu__abc_42281_new_n477_), .Y(alu__abc_42281_new_n2127_));
INVX1 INVX1_1032 ( .A(alu__abc_42281_new_n2159_), .Y(alu__abc_42281_new_n2160_));
INVX1 INVX1_1033 ( .A(alu__abc_42281_new_n2164_), .Y(alu__abc_42281_new_n2165_));
INVX1 INVX1_1034 ( .A(alu__abc_42281_new_n2201_), .Y(alu__abc_42281_new_n2202_));
INVX1 INVX1_1035 ( .A(alu__abc_42281_new_n2206_), .Y(alu__abc_42281_new_n2208_));
INVX1 INVX1_1036 ( .A(alu__abc_42281_new_n2242_), .Y(alu__abc_42281_new_n2243_));
INVX1 INVX1_1037 ( .A(alu__abc_42281_new_n480_), .Y(alu__abc_42281_new_n2247_));
INVX1 INVX1_1038 ( .A(alu__abc_42281_new_n2248_), .Y(alu__abc_42281_new_n2249_));
INVX1 INVX1_1039 ( .A(alu__abc_42281_new_n2282_), .Y(alu__abc_42281_new_n2283_));
INVX1 INVX1_104 ( .A(_abc_44694_new_n1470_), .Y(_abc_44694_new_n1471_));
INVX1 INVX1_1040 ( .A(alu__abc_42281_new_n2287_), .Y(alu__abc_42281_new_n2288_));
INVX1 INVX1_1041 ( .A(alu__abc_42281_new_n2321_), .Y(alu__abc_42281_new_n2322_));
INVX1 INVX1_1042 ( .A(alu__abc_42281_new_n2325_), .Y(alu__abc_42281_new_n2327_));
INVX1 INVX1_1043 ( .A(alu__abc_42281_new_n2360_), .Y(alu__abc_42281_new_n2361_));
INVX1 INVX1_1044 ( .A(alu__abc_42281_new_n506_), .Y(alu__abc_42281_new_n2366_));
INVX1 INVX1_1045 ( .A(alu__abc_42281_new_n826_), .Y(alu__abc_42281_new_n2398_));
INVX1 INVX1_1046 ( .A(alu_equal_o), .Y(alu__abc_42281_new_n2433_));
INVX1 INVX1_1047 ( .A(alu_less_than_signed_o), .Y(alu__abc_42281_new_n2434_));
INVX1 INVX1_1048 ( .A(alu__abc_42281_new_n2437_), .Y(alu__abc_42281_new_n2438_));
INVX1 INVX1_1049 ( .A(alu__abc_42281_new_n2519_), .Y(alu_greater_than_o));
INVX1 INVX1_105 ( .A(_abc_44694_new_n1466_), .Y(_abc_44694_new_n1473_));
INVX1 INVX1_106 ( .A(_abc_44694_new_n1484_), .Y(_abc_44694_new_n1485_));
INVX1 INVX1_107 ( .A(_abc_44694_new_n1499_), .Y(_abc_44694_new_n1500_));
INVX1 INVX1_108 ( .A(_abc_44694_new_n1505_), .Y(_abc_44694_new_n1506_));
INVX1 INVX1_109 ( .A(_abc_44694_new_n1507_), .Y(_abc_44694_new_n1508_));
INVX1 INVX1_11 ( .A(_abc_44694_new_n649_), .Y(_abc_44694_new_n650_));
INVX1 INVX1_110 ( .A(_abc_44694_new_n1509_), .Y(_abc_44694_new_n1510_));
INVX1 INVX1_111 ( .A(_abc_44694_new_n1537_), .Y(_abc_44694_new_n1538_));
INVX1 INVX1_112 ( .A(_abc_44694_new_n1550_), .Y(_abc_44694_new_n1551_));
INVX1 INVX1_113 ( .A(_abc_44694_new_n1554_), .Y(_abc_44694_new_n1555_));
INVX1 INVX1_114 ( .A(_abc_44694_new_n1576_), .Y(_abc_44694_new_n1577_));
INVX1 INVX1_115 ( .A(_abc_44694_new_n1584_), .Y(_abc_44694_new_n1585_));
INVX1 INVX1_116 ( .A(_abc_44694_new_n1590_), .Y(_abc_44694_new_n1591_));
INVX1 INVX1_117 ( .A(_abc_44694_new_n1592_), .Y(_abc_44694_new_n1593_));
INVX1 INVX1_118 ( .A(_abc_44694_new_n1615_), .Y(_abc_44694_new_n1616_));
INVX1 INVX1_119 ( .A(_abc_44694_new_n1622_), .Y(_abc_44694_new_n1623_));
INVX1 INVX1_12 ( .A(_abc_44694_new_n653_), .Y(_abc_44694_new_n654_));
INVX1 INVX1_120 ( .A(_abc_44694_new_n1626_), .Y(_abc_44694_new_n1627_));
INVX1 INVX1_121 ( .A(_abc_44694_new_n1630_), .Y(_abc_44694_new_n1631_));
INVX1 INVX1_122 ( .A(_abc_44694_new_n1652_), .Y(_abc_44694_new_n1653_));
INVX1 INVX1_123 ( .A(_abc_44694_new_n1048_), .Y(_abc_44694_new_n1659_));
INVX1 INVX1_124 ( .A(_abc_44694_new_n1662_), .Y(_abc_44694_new_n1663_));
INVX1 INVX1_125 ( .A(_abc_44694_new_n1667_), .Y(_abc_44694_new_n1668_));
INVX1 INVX1_126 ( .A(_abc_44694_new_n1670_), .Y(_abc_44694_new_n1671_));
INVX1 INVX1_127 ( .A(_abc_44694_new_n1694_), .Y(_abc_44694_new_n1695_));
INVX1 INVX1_128 ( .A(_abc_44694_new_n1699_), .Y(_abc_44694_new_n1700_));
INVX1 INVX1_129 ( .A(_abc_44694_new_n1701_), .Y(_abc_44694_new_n1702_));
INVX1 INVX1_13 ( .A(enable_i_bF_buf7), .Y(_abc_44694_new_n657_));
INVX1 INVX1_130 ( .A(_abc_44694_new_n1704_), .Y(_abc_44694_new_n1705_));
INVX1 INVX1_131 ( .A(_abc_44694_new_n1707_), .Y(_abc_44694_new_n1708_));
INVX1 INVX1_132 ( .A(_abc_44694_new_n1732_), .Y(_abc_44694_new_n1733_));
INVX1 INVX1_133 ( .A(_abc_44694_new_n1741_), .Y(_abc_44694_new_n1742_));
INVX1 INVX1_134 ( .A(_abc_44694_new_n1739_), .Y(_abc_44694_new_n1745_));
INVX1 INVX1_135 ( .A(_abc_44694_new_n1743_), .Y(_abc_44694_new_n1746_));
INVX1 INVX1_136 ( .A(_abc_44694_new_n1768_), .Y(_abc_44694_new_n1769_));
INVX1 INVX1_137 ( .A(_abc_44694_new_n1784_), .Y(_abc_44694_new_n1785_));
INVX1 INVX1_138 ( .A(_abc_44694_new_n1788_), .Y(_abc_44694_new_n1789_));
INVX1 INVX1_139 ( .A(_abc_44694_new_n1810_), .Y(_abc_44694_new_n1811_));
INVX1 INVX1_14 ( .A(mem_ack_i), .Y(_abc_44694_new_n664_));
INVX1 INVX1_140 ( .A(_abc_44694_new_n1818_), .Y(_abc_44694_new_n1819_));
INVX1 INVX1_141 ( .A(_abc_44694_new_n1824_), .Y(_abc_44694_new_n1825_));
INVX1 INVX1_142 ( .A(_abc_44694_new_n1826_), .Y(_abc_44694_new_n1827_));
INVX1 INVX1_143 ( .A(_abc_44694_new_n1849_), .Y(_abc_44694_new_n1850_));
INVX1 INVX1_144 ( .A(_abc_44694_new_n1857_), .Y(_abc_44694_new_n1858_));
INVX1 INVX1_145 ( .A(_abc_44694_new_n1860_), .Y(_abc_44694_new_n1861_));
INVX1 INVX1_146 ( .A(_abc_44694_new_n1863_), .Y(_abc_44694_new_n1864_));
INVX1 INVX1_147 ( .A(_abc_44694_new_n1886_), .Y(_abc_44694_new_n1887_));
INVX1 INVX1_148 ( .A(_abc_44694_new_n1893_), .Y(_abc_44694_new_n1894_));
INVX1 INVX1_149 ( .A(_abc_44694_new_n1896_), .Y(_abc_44694_new_n1897_));
INVX1 INVX1_15 ( .A(mem_offset_q_0_), .Y(_abc_44694_new_n674_));
INVX1 INVX1_150 ( .A(_abc_44694_new_n1898_), .Y(_abc_44694_new_n1900_));
INVX1 INVX1_151 ( .A(_abc_44694_new_n1922_), .Y(_abc_44694_new_n1923_));
INVX1 INVX1_152 ( .A(_abc_44694_new_n1856_), .Y(_abc_44694_new_n1934_));
INVX1 INVX1_153 ( .A(_abc_44694_new_n1942_), .Y(_abc_44694_new_n1943_));
INVX1 INVX1_154 ( .A(_abc_44694_new_n1946_), .Y(_abc_44694_new_n1947_));
INVX1 INVX1_155 ( .A(_abc_44694_new_n1968_), .Y(_abc_44694_new_n1969_));
INVX1 INVX1_156 ( .A(_abc_44694_new_n1976_), .Y(_abc_44694_new_n1977_));
INVX1 INVX1_157 ( .A(_abc_44694_new_n1979_), .Y(_abc_44694_new_n1980_));
INVX1 INVX1_158 ( .A(_abc_44694_new_n1981_), .Y(_abc_44694_new_n1982_));
INVX1 INVX1_159 ( .A(_abc_44694_new_n2004_), .Y(_abc_44694_new_n2005_));
INVX1 INVX1_16 ( .A(mem_offset_q_1_), .Y(_abc_44694_new_n680_));
INVX1 INVX1_160 ( .A(_abc_44694_new_n2011_), .Y(_abc_44694_new_n2012_));
INVX1 INVX1_161 ( .A(_abc_44694_new_n2014_), .Y(_abc_44694_new_n2015_));
INVX1 INVX1_162 ( .A(_abc_44694_new_n2017_), .Y(_abc_44694_new_n2018_));
INVX1 INVX1_163 ( .A(_abc_44694_new_n2040_), .Y(_abc_44694_new_n2041_));
INVX1 INVX1_164 ( .A(_abc_44694_new_n2049_), .Y(_abc_44694_new_n2050_));
INVX1 INVX1_165 ( .A(_abc_44694_new_n2051_), .Y(_abc_44694_new_n2052_));
INVX1 INVX1_166 ( .A(_abc_44694_new_n2047_), .Y(_abc_44694_new_n2054_));
INVX1 INVX1_167 ( .A(_abc_44694_new_n2076_), .Y(_abc_44694_new_n2077_));
INVX1 INVX1_168 ( .A(_abc_44694_new_n2089_), .Y(_abc_44694_new_n2090_));
INVX1 INVX1_169 ( .A(_abc_44694_new_n1940_), .Y(_abc_44694_new_n2091_));
INVX1 INVX1_17 ( .A(sr_q_2_), .Y(_abc_44694_new_n971_));
INVX1 INVX1_170 ( .A(_abc_44694_new_n2093_), .Y(_abc_44694_new_n2094_));
INVX1 INVX1_171 ( .A(_abc_44694_new_n2096_), .Y(_abc_44694_new_n2097_));
INVX1 INVX1_172 ( .A(_abc_44694_new_n2099_), .Y(_abc_44694_new_n2100_));
INVX1 INVX1_173 ( .A(_abc_44694_new_n2102_), .Y(_abc_44694_new_n2103_));
INVX1 INVX1_174 ( .A(_abc_44694_new_n2125_), .Y(_abc_44694_new_n2126_));
INVX1 INVX1_175 ( .A(_abc_44694_new_n2133_), .Y(_abc_44694_new_n2134_));
INVX1 INVX1_176 ( .A(_abc_44694_new_n2139_), .Y(_abc_44694_new_n2140_));
INVX1 INVX1_177 ( .A(_abc_44694_new_n2141_), .Y(_abc_44694_new_n2142_));
INVX1 INVX1_178 ( .A(_abc_44694_new_n2164_), .Y(_abc_44694_new_n2165_));
INVX1 INVX1_179 ( .A(_abc_44694_new_n2172_), .Y(_abc_44694_new_n2173_));
INVX1 INVX1_18 ( .A(_abc_44694_new_n972_), .Y(_abc_44694_new_n973_));
INVX1 INVX1_180 ( .A(_abc_44694_new_n2175_), .Y(_abc_44694_new_n2176_));
INVX1 INVX1_181 ( .A(_abc_44694_new_n2178_), .Y(_abc_44694_new_n2179_));
INVX1 INVX1_182 ( .A(_abc_44694_new_n2201_), .Y(_abc_44694_new_n2202_));
INVX1 INVX1_183 ( .A(_abc_44694_new_n2208_), .Y(_abc_44694_new_n2209_));
INVX1 INVX1_184 ( .A(_abc_44694_new_n2211_), .Y(_abc_44694_new_n2212_));
INVX1 INVX1_185 ( .A(_abc_44694_new_n2213_), .Y(_abc_44694_new_n2215_));
INVX1 INVX1_186 ( .A(_abc_44694_new_n2237_), .Y(_abc_44694_new_n2238_));
INVX1 INVX1_187 ( .A(_abc_44694_new_n2171_), .Y(_abc_44694_new_n2246_));
INVX1 INVX1_188 ( .A(_abc_44694_new_n2255_), .Y(_abc_44694_new_n2256_));
INVX1 INVX1_189 ( .A(_abc_44694_new_n2259_), .Y(_abc_44694_new_n2260_));
INVX1 INVX1_19 ( .A(_abc_44694_new_n974_), .Y(_abc_44694_new_n975_));
INVX1 INVX1_190 ( .A(_abc_44694_new_n2283_), .Y(_abc_44694_new_n2284_));
INVX1 INVX1_191 ( .A(_abc_44694_new_n2289_), .Y(_abc_44694_new_n2290_));
INVX1 INVX1_192 ( .A(_abc_44694_new_n2295_), .Y(_abc_44694_new_n2296_));
INVX1 INVX1_193 ( .A(_abc_44694_new_n2297_), .Y(_abc_44694_new_n2298_));
INVX1 INVX1_194 ( .A(_abc_44694_new_n2322_), .Y(_abc_44694_new_n2323_));
INVX1 INVX1_195 ( .A(_abc_44694_new_n2327_), .Y(_abc_44694_new_n2328_));
INVX1 INVX1_196 ( .A(_abc_44694_new_n2331_), .Y(_abc_44694_new_n2332_));
INVX1 INVX1_197 ( .A(_abc_44694_new_n2335_), .Y(_abc_44694_new_n2336_));
INVX1 INVX1_198 ( .A(_abc_44694_new_n2359_), .Y(_abc_44694_new_n2360_));
INVX1 INVX1_199 ( .A(_abc_44694_new_n2365_), .Y(_abc_44694_new_n2366_));
INVX1 INVX1_2 ( .A(inst_r_5_), .Y(_abc_44694_new_n618_));
INVX1 INVX1_20 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_44694_new_n977_));
INVX1 INVX1_200 ( .A(_abc_44694_new_n2371_), .Y(_abc_44694_new_n2372_));
INVX1 INVX1_201 ( .A(_abc_44694_new_n2373_), .Y(_abc_44694_new_n2374_));
INVX1 INVX1_202 ( .A(_abc_44694_new_n2398_), .Y(_abc_44694_new_n2399_));
INVX1 INVX1_203 ( .A(_abc_44694_new_n2403_), .Y(_abc_44694_new_n2404_));
INVX1 INVX1_204 ( .A(_abc_44694_new_n2407_), .Y(_abc_44694_new_n2408_));
INVX1 INVX1_205 ( .A(_abc_44694_new_n2411_), .Y(_abc_44694_new_n2412_));
INVX1 INVX1_206 ( .A(_abc_44694_new_n2435_), .Y(_abc_44694_new_n2436_));
INVX1 INVX1_207 ( .A(_abc_44694_new_n2440_), .Y(_abc_44694_new_n2441_));
INVX1 INVX1_208 ( .A(_abc_44694_new_n2443_), .Y(_abc_44694_new_n2444_));
INVX1 INVX1_209 ( .A(_abc_44694_new_n2445_), .Y(_abc_44694_new_n2447_));
INVX1 INVX1_21 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_44694_new_n978_));
INVX1 INVX1_210 ( .A(_abc_44694_new_n2471_), .Y(_abc_44694_new_n2472_));
INVX1 INVX1_211 ( .A(_abc_44694_new_n2477_), .Y(_abc_44694_new_n2478_));
INVX1 INVX1_212 ( .A(_abc_44694_new_n2479_), .Y(_abc_44694_new_n2480_));
INVX1 INVX1_213 ( .A(pc_q_30_), .Y(_abc_44694_new_n2481_));
INVX1 INVX1_214 ( .A(_abc_44694_new_n2482_), .Y(_abc_44694_new_n2483_));
INVX1 INVX1_215 ( .A(_abc_44694_new_n2484_), .Y(_abc_44694_new_n2485_));
INVX1 INVX1_216 ( .A(_abc_44694_new_n2486_), .Y(_abc_44694_new_n2488_));
INVX1 INVX1_217 ( .A(_abc_44694_new_n2512_), .Y(_abc_44694_new_n2513_));
INVX1 INVX1_218 ( .A(pc_q_31_), .Y(_abc_44694_new_n2517_));
INVX1 INVX1_219 ( .A(_abc_44694_new_n2518_), .Y(_abc_44694_new_n2519_));
INVX1 INVX1_22 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_15_), .Y(_abc_44694_new_n979_));
INVX1 INVX1_220 ( .A(_abc_44694_new_n2521_), .Y(_abc_44694_new_n2522_));
INVX1 INVX1_221 ( .A(_abc_44694_new_n1203_), .Y(_abc_44694_new_n2608_));
INVX1 INVX1_222 ( .A(_abc_44694_new_n1191_), .Y(_abc_44694_new_n2716_));
INVX1 INVX1_223 ( .A(_abc_44694_new_n2743_), .Y(_abc_44694_new_n2744_));
INVX1 INVX1_224 ( .A(_abc_44694_new_n2773_), .Y(_abc_44694_new_n2774_));
INVX1 INVX1_225 ( .A(_abc_44694_new_n1181__bF_buf2), .Y(_abc_44694_new_n2831_));
INVX1 INVX1_226 ( .A(REGFILE_SIM_reg_bank_rb_i_4_bF_buf0_), .Y(_abc_44694_new_n2833_));
INVX1 INVX1_227 ( .A(_abc_44694_new_n668__bF_buf3), .Y(_abc_44694_new_n3331_));
INVX1 INVX1_228 ( .A(_abc_44694_new_n3332_), .Y(_abc_44694_new_n3333_));
INVX1 INVX1_229 ( .A(_abc_44694_new_n3339_), .Y(_abc_44694_new_n3340_));
INVX1 INVX1_23 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_44694_new_n982_));
INVX1 INVX1_230 ( .A(_abc_44694_new_n3341_), .Y(_abc_44694_new_n3343_));
INVX1 INVX1_231 ( .A(_abc_44694_new_n3345_), .Y(_abc_44694_new_n3346_));
INVX1 INVX1_232 ( .A(\mem_dat_i[0] ), .Y(_abc_44694_new_n3351_));
INVX1 INVX1_233 ( .A(_abc_44694_new_n3352_), .Y(_abc_44694_new_n3353_));
INVX1 INVX1_234 ( .A(\mem_dat_i[1] ), .Y(_abc_44694_new_n3356_));
INVX1 INVX1_235 ( .A(_abc_44694_new_n3357_), .Y(_abc_44694_new_n3358_));
INVX1 INVX1_236 ( .A(\mem_dat_i[2] ), .Y(_abc_44694_new_n3361_));
INVX1 INVX1_237 ( .A(_abc_44694_new_n3362_), .Y(_abc_44694_new_n3363_));
INVX1 INVX1_238 ( .A(\mem_dat_i[3] ), .Y(_abc_44694_new_n3366_));
INVX1 INVX1_239 ( .A(_abc_44694_new_n3367_), .Y(_abc_44694_new_n3368_));
INVX1 INVX1_24 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_44694_new_n983_));
INVX1 INVX1_240 ( .A(\mem_dat_i[4] ), .Y(_abc_44694_new_n3371_));
INVX1 INVX1_241 ( .A(_abc_44694_new_n3372_), .Y(_abc_44694_new_n3373_));
INVX1 INVX1_242 ( .A(\mem_dat_i[5] ), .Y(_abc_44694_new_n3376_));
INVX1 INVX1_243 ( .A(_abc_44694_new_n3377_), .Y(_abc_44694_new_n3378_));
INVX1 INVX1_244 ( .A(\mem_dat_i[6] ), .Y(_abc_44694_new_n3381_));
INVX1 INVX1_245 ( .A(_abc_44694_new_n3382_), .Y(_abc_44694_new_n3383_));
INVX1 INVX1_246 ( .A(\mem_dat_i[7] ), .Y(_abc_44694_new_n3386_));
INVX1 INVX1_247 ( .A(_abc_44694_new_n3387_), .Y(_abc_44694_new_n3388_));
INVX1 INVX1_248 ( .A(\mem_dat_i[8] ), .Y(_abc_44694_new_n3391_));
INVX1 INVX1_249 ( .A(_abc_44694_new_n3392_), .Y(_abc_44694_new_n3393_));
INVX1 INVX1_25 ( .A(_abc_44694_new_n985_), .Y(_abc_44694_new_n986_));
INVX1 INVX1_250 ( .A(\mem_dat_i[9] ), .Y(_abc_44694_new_n3396_));
INVX1 INVX1_251 ( .A(_abc_44694_new_n3397_), .Y(_abc_44694_new_n3398_));
INVX1 INVX1_252 ( .A(\mem_dat_i[10] ), .Y(_abc_44694_new_n3401_));
INVX1 INVX1_253 ( .A(_abc_44694_new_n3402_), .Y(_abc_44694_new_n3403_));
INVX1 INVX1_254 ( .A(\mem_dat_i[11] ), .Y(_abc_44694_new_n3406_));
INVX1 INVX1_255 ( .A(_abc_44694_new_n3407_), .Y(_abc_44694_new_n3408_));
INVX1 INVX1_256 ( .A(\mem_dat_i[12] ), .Y(_abc_44694_new_n3411_));
INVX1 INVX1_257 ( .A(_abc_44694_new_n3412_), .Y(_abc_44694_new_n3413_));
INVX1 INVX1_258 ( .A(\mem_dat_i[13] ), .Y(_abc_44694_new_n3416_));
INVX1 INVX1_259 ( .A(_abc_44694_new_n3417_), .Y(_abc_44694_new_n3418_));
INVX1 INVX1_26 ( .A(_abc_44694_new_n990_), .Y(_abc_44694_new_n991_));
INVX1 INVX1_260 ( .A(\mem_dat_i[14] ), .Y(_abc_44694_new_n3421_));
INVX1 INVX1_261 ( .A(_abc_44694_new_n3422_), .Y(_abc_44694_new_n3423_));
INVX1 INVX1_262 ( .A(\mem_dat_i[15] ), .Y(_abc_44694_new_n3426_));
INVX1 INVX1_263 ( .A(_abc_44694_new_n3427_), .Y(_abc_44694_new_n3428_));
INVX1 INVX1_264 ( .A(\mem_dat_i[16] ), .Y(_abc_44694_new_n3431_));
INVX1 INVX1_265 ( .A(_abc_44694_new_n3432_), .Y(_abc_44694_new_n3433_));
INVX1 INVX1_266 ( .A(\mem_dat_i[17] ), .Y(_abc_44694_new_n3436_));
INVX1 INVX1_267 ( .A(_abc_44694_new_n3437_), .Y(_abc_44694_new_n3438_));
INVX1 INVX1_268 ( .A(\mem_dat_i[18] ), .Y(_abc_44694_new_n3441_));
INVX1 INVX1_269 ( .A(_abc_44694_new_n3442_), .Y(_abc_44694_new_n3443_));
INVX1 INVX1_27 ( .A(_abc_44694_new_n995_), .Y(_abc_44694_new_n996_));
INVX1 INVX1_270 ( .A(\mem_dat_i[19] ), .Y(_abc_44694_new_n3446_));
INVX1 INVX1_271 ( .A(_abc_44694_new_n3447_), .Y(_abc_44694_new_n3448_));
INVX1 INVX1_272 ( .A(\mem_dat_i[20] ), .Y(_abc_44694_new_n3451_));
INVX1 INVX1_273 ( .A(_abc_44694_new_n3452_), .Y(_abc_44694_new_n3453_));
INVX1 INVX1_274 ( .A(\mem_dat_i[21] ), .Y(_abc_44694_new_n3456_));
INVX1 INVX1_275 ( .A(_abc_44694_new_n3457_), .Y(_abc_44694_new_n3458_));
INVX1 INVX1_276 ( .A(\mem_dat_i[22] ), .Y(_abc_44694_new_n3461_));
INVX1 INVX1_277 ( .A(_abc_44694_new_n3462_), .Y(_abc_44694_new_n3463_));
INVX1 INVX1_278 ( .A(\mem_dat_i[23] ), .Y(_abc_44694_new_n3466_));
INVX1 INVX1_279 ( .A(_abc_44694_new_n3467_), .Y(_abc_44694_new_n3468_));
INVX1 INVX1_28 ( .A(_abc_44694_new_n999_), .Y(_abc_44694_new_n1000_));
INVX1 INVX1_280 ( .A(\mem_dat_i[24] ), .Y(_abc_44694_new_n3471_));
INVX1 INVX1_281 ( .A(_abc_44694_new_n3472_), .Y(_abc_44694_new_n3473_));
INVX1 INVX1_282 ( .A(\mem_dat_i[25] ), .Y(_abc_44694_new_n3476_));
INVX1 INVX1_283 ( .A(_abc_44694_new_n3477_), .Y(_abc_44694_new_n3478_));
INVX1 INVX1_284 ( .A(\mem_dat_i[26] ), .Y(_abc_44694_new_n3481_));
INVX1 INVX1_285 ( .A(_abc_44694_new_n3482_), .Y(_abc_44694_new_n3483_));
INVX1 INVX1_286 ( .A(\mem_dat_i[27] ), .Y(_abc_44694_new_n3486_));
INVX1 INVX1_287 ( .A(_abc_44694_new_n3487_), .Y(_abc_44694_new_n3488_));
INVX1 INVX1_288 ( .A(\mem_dat_i[28] ), .Y(_abc_44694_new_n3491_));
INVX1 INVX1_289 ( .A(_abc_44694_new_n3492_), .Y(_abc_44694_new_n3493_));
INVX1 INVX1_29 ( .A(_abc_44694_new_n1001_), .Y(_abc_44694_new_n1002_));
INVX1 INVX1_290 ( .A(\mem_dat_i[29] ), .Y(_abc_44694_new_n3496_));
INVX1 INVX1_291 ( .A(_abc_44694_new_n3497_), .Y(_abc_44694_new_n3498_));
INVX1 INVX1_292 ( .A(\mem_dat_i[30] ), .Y(_abc_44694_new_n3501_));
INVX1 INVX1_293 ( .A(_abc_44694_new_n3502_), .Y(_abc_44694_new_n3503_));
INVX1 INVX1_294 ( .A(\mem_dat_i[31] ), .Y(_abc_44694_new_n3506_));
INVX1 INVX1_295 ( .A(_abc_44694_new_n3507_), .Y(_abc_44694_new_n3508_));
INVX1 INVX1_296 ( .A(_abc_44694_new_n3334__bF_buf3), .Y(_abc_44694_new_n3514_));
INVX1 INVX1_297 ( .A(_abc_44694_new_n3522_), .Y(_abc_44694_new_n3523_));
INVX1 INVX1_298 ( .A(_abc_44694_new_n3537_), .Y(_abc_44694_new_n3538_));
INVX1 INVX1_299 ( .A(state_q_3_bF_buf4_), .Y(_abc_44694_new_n4046_));
INVX1 INVX1_3 ( .A(inst_r_2_), .Y(_abc_44694_new_n620_));
INVX1 INVX1_30 ( .A(_abc_44694_new_n1004_), .Y(_abc_44694_new_n1005_));
INVX1 INVX1_300 ( .A(state_q_2_), .Y(_abc_44694_new_n4056_));
INVX1 INVX1_301 ( .A(_abc_44694_new_n4073_), .Y(_abc_44694_new_n4074_));
INVX1 INVX1_302 ( .A(_abc_44694_new_n4076_), .Y(_abc_44694_new_n4077_));
INVX1 INVX1_303 ( .A(_abc_44694_new_n4085_), .Y(_abc_44694_new_n4086_));
INVX1 INVX1_304 ( .A(_abc_44694_new_n4087_), .Y(_abc_44694_new_n4088_));
INVX1 INVX1_305 ( .A(_abc_44694_new_n4089_), .Y(_abc_44694_new_n4091_));
INVX1 INVX1_306 ( .A(_abc_44694_new_n4097_), .Y(_abc_44694_new_n4098_));
INVX1 INVX1_307 ( .A(_abc_44694_new_n4101_), .Y(_abc_44694_new_n4102_));
INVX1 INVX1_308 ( .A(_abc_44694_new_n4099_), .Y(_abc_44694_new_n4104_));
INVX1 INVX1_309 ( .A(_abc_44694_new_n4113_), .Y(_abc_44694_new_n4114_));
INVX1 INVX1_31 ( .A(_abc_44694_new_n1006_), .Y(_abc_44694_new_n1007_));
INVX1 INVX1_310 ( .A(_abc_44694_new_n4115_), .Y(_abc_44694_new_n4116_));
INVX1 INVX1_311 ( .A(_abc_44694_new_n4112_), .Y(_abc_44694_new_n4118_));
INVX1 INVX1_312 ( .A(_abc_44694_new_n4126_), .Y(_abc_44694_new_n4127_));
INVX1 INVX1_313 ( .A(_abc_44694_new_n4128_), .Y(_abc_44694_new_n4129_));
INVX1 INVX1_314 ( .A(_abc_44694_new_n4132_), .Y(_abc_44694_new_n4133_));
INVX1 INVX1_315 ( .A(_abc_44694_new_n4142_), .Y(_abc_44694_new_n4143_));
INVX1 INVX1_316 ( .A(_abc_44694_new_n4144_), .Y(_abc_44694_new_n4145_));
INVX1 INVX1_317 ( .A(_abc_44694_new_n4146_), .Y(_abc_44694_new_n4147_));
INVX1 INVX1_318 ( .A(_abc_44694_new_n4158_), .Y(_abc_44694_new_n4159_));
INVX1 INVX1_319 ( .A(_abc_44694_new_n4160_), .Y(_abc_44694_new_n4161_));
INVX1 INVX1_32 ( .A(_abc_44694_new_n1013_), .Y(_abc_44694_new_n1014_));
INVX1 INVX1_320 ( .A(_abc_44694_new_n4163_), .Y(_abc_44694_new_n4164_));
INVX1 INVX1_321 ( .A(_abc_44694_new_n4165_), .Y(_abc_44694_new_n4166_));
INVX1 INVX1_322 ( .A(_abc_44694_new_n4169_), .Y(_abc_44694_new_n4170_));
INVX1 INVX1_323 ( .A(_abc_44694_new_n4177_), .Y(_abc_44694_new_n4178_));
INVX1 INVX1_324 ( .A(_abc_44694_new_n4180_), .Y(_abc_44694_new_n4181_));
INVX1 INVX1_325 ( .A(_abc_44694_new_n4182_), .Y(_abc_44694_new_n4183_));
INVX1 INVX1_326 ( .A(_abc_44694_new_n4191_), .Y(_abc_44694_new_n4192_));
INVX1 INVX1_327 ( .A(_abc_44694_new_n4195_), .Y(_abc_44694_new_n4196_));
INVX1 INVX1_328 ( .A(_abc_44694_new_n4197_), .Y(_abc_44694_new_n4198_));
INVX1 INVX1_329 ( .A(_abc_44694_new_n4199_), .Y(_abc_44694_new_n4200_));
INVX1 INVX1_33 ( .A(_abc_44694_new_n970_), .Y(_abc_44694_new_n1017_));
INVX1 INVX1_330 ( .A(_abc_44694_new_n4202_), .Y(_abc_44694_new_n4203_));
INVX1 INVX1_331 ( .A(_abc_44694_new_n4215_), .Y(_abc_44694_new_n4216_));
INVX1 INVX1_332 ( .A(_abc_44694_new_n4211_), .Y(_abc_44694_new_n4220_));
INVX1 INVX1_333 ( .A(_abc_44694_new_n4218_), .Y(_abc_44694_new_n4221_));
INVX1 INVX1_334 ( .A(_abc_44694_new_n4232_), .Y(_abc_44694_new_n4233_));
INVX1 INVX1_335 ( .A(_abc_44694_new_n4245_), .Y(_abc_44694_new_n4246_));
INVX1 INVX1_336 ( .A(_abc_44694_new_n4256_), .Y(_abc_44694_new_n4257_));
INVX1 INVX1_337 ( .A(_abc_44694_new_n4263_), .Y(_abc_44694_new_n4264_));
INVX1 INVX1_338 ( .A(_abc_44694_new_n4265_), .Y(_abc_44694_new_n4266_));
INVX1 INVX1_339 ( .A(_abc_44694_new_n4275_), .Y(_abc_44694_new_n4276_));
INVX1 INVX1_34 ( .A(_abc_44694_new_n1023_), .Y(_abc_44694_new_n1024_));
INVX1 INVX1_340 ( .A(_abc_44694_new_n4280_), .Y(_abc_44694_new_n4281_));
INVX1 INVX1_341 ( .A(_abc_44694_new_n4285_), .Y(_abc_44694_new_n4286_));
INVX1 INVX1_342 ( .A(_abc_44694_new_n4293_), .Y(_abc_44694_new_n4294_));
INVX1 INVX1_343 ( .A(_abc_44694_new_n4298_), .Y(_abc_44694_new_n4299_));
INVX1 INVX1_344 ( .A(_abc_44694_new_n4301_), .Y(_abc_44694_new_n4302_));
INVX1 INVX1_345 ( .A(_abc_44694_new_n4303_), .Y(_abc_44694_new_n4304_));
INVX1 INVX1_346 ( .A(_abc_44694_new_n4316_), .Y(_abc_44694_new_n4317_));
INVX1 INVX1_347 ( .A(_abc_44694_new_n4321_), .Y(_abc_44694_new_n4322_));
INVX1 INVX1_348 ( .A(_abc_44694_new_n4323_), .Y(_abc_44694_new_n4324_));
INVX1 INVX1_349 ( .A(_abc_44694_new_n4330_), .Y(_abc_44694_new_n4331_));
INVX1 INVX1_35 ( .A(_abc_44694_new_n1026_), .Y(_abc_44694_new_n1027_));
INVX1 INVX1_350 ( .A(_abc_44694_new_n4338_), .Y(_abc_44694_new_n4339_));
INVX1 INVX1_351 ( .A(_abc_44694_new_n4340_), .Y(_abc_44694_new_n4341_));
INVX1 INVX1_352 ( .A(_abc_44694_new_n4343_), .Y(_abc_44694_new_n4344_));
INVX1 INVX1_353 ( .A(_abc_44694_new_n4356_), .Y(_abc_44694_new_n4357_));
INVX1 INVX1_354 ( .A(_abc_44694_new_n4360_), .Y(_abc_44694_new_n4361_));
INVX1 INVX1_355 ( .A(_abc_44694_new_n4366_), .Y(_abc_44694_new_n4367_));
INVX1 INVX1_356 ( .A(_abc_44694_new_n4374_), .Y(_abc_44694_new_n4375_));
INVX1 INVX1_357 ( .A(_abc_44694_new_n4376_), .Y(_abc_44694_new_n4377_));
INVX1 INVX1_358 ( .A(_abc_44694_new_n4379_), .Y(_abc_44694_new_n4380_));
INVX1 INVX1_359 ( .A(_abc_44694_new_n4395_), .Y(_abc_44694_new_n4396_));
INVX1 INVX1_36 ( .A(_abc_44694_new_n992_), .Y(_abc_44694_new_n1029_));
INVX1 INVX1_360 ( .A(_abc_44694_new_n4398_), .Y(_abc_44694_new_n4399_));
INVX1 INVX1_361 ( .A(_abc_44694_new_n4401_), .Y(_abc_44694_new_n4402_));
INVX1 INVX1_362 ( .A(_abc_44694_new_n4406_), .Y(_abc_44694_new_n4407_));
INVX1 INVX1_363 ( .A(_abc_44694_new_n4415_), .Y(_abc_44694_new_n4416_));
INVX1 INVX1_364 ( .A(_abc_44694_new_n4418_), .Y(_abc_44694_new_n4419_));
INVX1 INVX1_365 ( .A(_abc_44694_new_n4414_), .Y(_abc_44694_new_n4421_));
INVX1 INVX1_366 ( .A(_abc_44694_new_n4429_), .Y(_abc_44694_new_n4430_));
INVX1 INVX1_367 ( .A(_abc_44694_new_n4433_), .Y(_abc_44694_new_n4434_));
INVX1 INVX1_368 ( .A(_abc_44694_new_n4439_), .Y(_abc_44694_new_n4440_));
INVX1 INVX1_369 ( .A(_abc_44694_new_n4447_), .Y(_abc_44694_new_n4448_));
INVX1 INVX1_37 ( .A(_abc_44694_new_n994_), .Y(_abc_44694_new_n1032_));
INVX1 INVX1_370 ( .A(_abc_44694_new_n4449_), .Y(_abc_44694_new_n4450_));
INVX1 INVX1_371 ( .A(_abc_44694_new_n4452_), .Y(_abc_44694_new_n4453_));
INVX1 INVX1_372 ( .A(_abc_44694_new_n4466_), .Y(_abc_44694_new_n4467_));
INVX1 INVX1_373 ( .A(_abc_44694_new_n4470_), .Y(_abc_44694_new_n4471_));
INVX1 INVX1_374 ( .A(_abc_44694_new_n4328_), .Y(_abc_44694_new_n4474_));
INVX1 INVX1_375 ( .A(_abc_44694_new_n4475_), .Y(_abc_44694_new_n4476_));
INVX1 INVX1_376 ( .A(_abc_44694_new_n4478_), .Y(_abc_44694_new_n4479_));
INVX1 INVX1_377 ( .A(_abc_44694_new_n4480_), .Y(_abc_44694_new_n4481_));
INVX1 INVX1_378 ( .A(_abc_44694_new_n4485_), .Y(_abc_44694_new_n4486_));
INVX1 INVX1_379 ( .A(_abc_44694_new_n4493_), .Y(_abc_44694_new_n4494_));
INVX1 INVX1_38 ( .A(_abc_44694_new_n1038_), .Y(_abc_44694_new_n1039_));
INVX1 INVX1_380 ( .A(_abc_44694_new_n4495_), .Y(_abc_44694_new_n4496_));
INVX1 INVX1_381 ( .A(_abc_44694_new_n4498_), .Y(_abc_44694_new_n4499_));
INVX1 INVX1_382 ( .A(_abc_44694_new_n4511_), .Y(_abc_44694_new_n4512_));
INVX1 INVX1_383 ( .A(_abc_44694_new_n4515_), .Y(_abc_44694_new_n4516_));
INVX1 INVX1_384 ( .A(_abc_44694_new_n4517_), .Y(_abc_44694_new_n4518_));
INVX1 INVX1_385 ( .A(_abc_44694_new_n4522_), .Y(_abc_44694_new_n4523_));
INVX1 INVX1_386 ( .A(_abc_44694_new_n4530_), .Y(_abc_44694_new_n4531_));
INVX1 INVX1_387 ( .A(_abc_44694_new_n4532_), .Y(_abc_44694_new_n4533_));
INVX1 INVX1_388 ( .A(_abc_44694_new_n4535_), .Y(_abc_44694_new_n4537_));
INVX1 INVX1_389 ( .A(_abc_44694_new_n4547_), .Y(_abc_44694_new_n4548_));
INVX1 INVX1_39 ( .A(_abc_44694_new_n1044_), .Y(_abc_44694_new_n1045_));
INVX1 INVX1_390 ( .A(_abc_44694_new_n4545_), .Y(_abc_44694_new_n4549_));
INVX1 INVX1_391 ( .A(_abc_44694_new_n4553_), .Y(_abc_44694_new_n4554_));
INVX1 INVX1_392 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_28_), .Y(_abc_44694_new_n4556_));
INVX1 INVX1_393 ( .A(_abc_44694_new_n4558_), .Y(_abc_44694_new_n4559_));
INVX1 INVX1_394 ( .A(_abc_44694_new_n4561_), .Y(_abc_44694_new_n4562_));
INVX1 INVX1_395 ( .A(_abc_44694_new_n4569_), .Y(_abc_44694_new_n4570_));
INVX1 INVX1_396 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_29_), .Y(_abc_44694_new_n4572_));
INVX1 INVX1_397 ( .A(_abc_44694_new_n4574_), .Y(_abc_44694_new_n4575_));
INVX1 INVX1_398 ( .A(_abc_44694_new_n4587_), .Y(_abc_44694_new_n4588_));
INVX1 INVX1_399 ( .A(_abc_44694_new_n4593_), .Y(_abc_44694_new_n4594_));
INVX1 INVX1_4 ( .A(opcode_q_25_), .Y(_abc_44694_new_n623_));
INVX1 INVX1_40 ( .A(opcode_q_24_), .Y(_abc_44694_new_n1046_));
INVX1 INVX1_400 ( .A(_abc_44694_new_n4596_), .Y(_abc_44694_new_n4597_));
INVX1 INVX1_401 ( .A(_abc_44694_new_n4590_), .Y(_abc_44694_new_n4599_));
INVX1 INVX1_402 ( .A(_abc_44694_new_n4607_), .Y(_abc_44694_new_n4608_));
INVX1 INVX1_403 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_44694_new_n4609_));
INVX1 INVX1_404 ( .A(_abc_44694_new_n4612_), .Y(_abc_44694_new_n4613_));
INVX1 INVX1_405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2106_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2107_));
INVX1 INVX1_406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2111_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2112_));
INVX1 INVX1_407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2117_));
INVX1 INVX1_408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2121_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2122_));
INVX1 INVX1_409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2126_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2127_));
INVX1 INVX1_41 ( .A(_abc_44694_new_n1049_), .Y(_abc_44694_new_n1050_));
INVX1 INVX1_410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2131_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2132_));
INVX1 INVX1_411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2136_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2137_));
INVX1 INVX1_412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2141_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2142_));
INVX1 INVX1_413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2146_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2147_));
INVX1 INVX1_414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2151_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2152_));
INVX1 INVX1_415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2156_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2157_));
INVX1 INVX1_416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2161_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2162_));
INVX1 INVX1_417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2166_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2167_));
INVX1 INVX1_418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2171_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2172_));
INVX1 INVX1_419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2176_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2177_));
INVX1 INVX1_42 ( .A(alu_op_r_2_), .Y(_abc_44694_new_n1053_));
INVX1 INVX1_420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2181_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2182_));
INVX1 INVX1_421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2186_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2187_));
INVX1 INVX1_422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2191_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2192_));
INVX1 INVX1_423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2196_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2197_));
INVX1 INVX1_424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2201_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2202_));
INVX1 INVX1_425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2206_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2207_));
INVX1 INVX1_426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2211_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2212_));
INVX1 INVX1_427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2216_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2217_));
INVX1 INVX1_428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2221_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2222_));
INVX1 INVX1_429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2226_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2227_));
INVX1 INVX1_43 ( .A(alu_op_r_3_), .Y(_abc_44694_new_n1054_));
INVX1 INVX1_430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2231_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2232_));
INVX1 INVX1_431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2236_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2237_));
INVX1 INVX1_432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2242_));
INVX1 INVX1_433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2246_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2247_));
INVX1 INVX1_434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2251_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2252_));
INVX1 INVX1_435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2256_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2257_));
INVX1 INVX1_436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2261_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2262_));
INVX1 INVX1_437 ( .A(REGFILE_SIM_reg_bank_rd_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2264_));
INVX1 INVX1_438 ( .A(REGFILE_SIM_reg_bank_rd_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2365_));
INVX1 INVX1_439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2470_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2471_));
INVX1 INVX1_44 ( .A(alu_op_r_4_), .Y(_abc_44694_new_n1056_));
INVX1 INVX1_440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2474_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2475_));
INVX1 INVX1_441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2478_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2479_));
INVX1 INVX1_442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2482_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2483_));
INVX1 INVX1_443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2486_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2487_));
INVX1 INVX1_444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2490_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2491_));
INVX1 INVX1_445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2494_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2495_));
INVX1 INVX1_446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2498_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2499_));
INVX1 INVX1_447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2502_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2503_));
INVX1 INVX1_448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2506_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2507_));
INVX1 INVX1_449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2510_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2511_));
INVX1 INVX1_45 ( .A(alu_op_r_5_), .Y(_abc_44694_new_n1057_));
INVX1 INVX1_450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2514_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2515_));
INVX1 INVX1_451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2518_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2519_));
INVX1 INVX1_452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2522_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2523_));
INVX1 INVX1_453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2526_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2527_));
INVX1 INVX1_454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2530_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2531_));
INVX1 INVX1_455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2534_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2535_));
INVX1 INVX1_456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2538_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2539_));
INVX1 INVX1_457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2542_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2543_));
INVX1 INVX1_458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2546_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2547_));
INVX1 INVX1_459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2550_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2551_));
INVX1 INVX1_46 ( .A(alu_op_r_6_), .Y(_abc_44694_new_n1059_));
INVX1 INVX1_460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2555_));
INVX1 INVX1_461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2558_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2559_));
INVX1 INVX1_462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2562_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2563_));
INVX1 INVX1_463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2566_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2567_));
INVX1 INVX1_464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2570_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2571_));
INVX1 INVX1_465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2575_));
INVX1 INVX1_466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2579_));
INVX1 INVX1_467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2583_));
INVX1 INVX1_468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2586_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2587_));
INVX1 INVX1_469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2590_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2591_));
INVX1 INVX1_47 ( .A(alu_op_r_7_), .Y(_abc_44694_new_n1060_));
INVX1 INVX1_470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2595_));
INVX1 INVX1_471 ( .A(REGFILE_SIM_reg_bank_rd_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2597_));
INVX1 INVX1_472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2701_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2702_));
INVX1 INVX1_473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2705_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2706_));
INVX1 INVX1_474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2709_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2710_));
INVX1 INVX1_475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2713_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2714_));
INVX1 INVX1_476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2718_));
INVX1 INVX1_477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2721_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2722_));
INVX1 INVX1_478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2725_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2726_));
INVX1 INVX1_479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2729_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2730_));
INVX1 INVX1_48 ( .A(alu_op_r_0_), .Y(_abc_44694_new_n1063_));
INVX1 INVX1_480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2733_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2734_));
INVX1 INVX1_481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2737_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2738_));
INVX1 INVX1_482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2741_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2742_));
INVX1 INVX1_483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2745_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2746_));
INVX1 INVX1_484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2749_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2750_));
INVX1 INVX1_485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2753_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2754_));
INVX1 INVX1_486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2757_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2758_));
INVX1 INVX1_487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2761_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2762_));
INVX1 INVX1_488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2765_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2766_));
INVX1 INVX1_489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2769_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2770_));
INVX1 INVX1_49 ( .A(alu_op_r_1_), .Y(_abc_44694_new_n1064_));
INVX1 INVX1_490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2773_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2774_));
INVX1 INVX1_491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2777_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2778_));
INVX1 INVX1_492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2781_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2782_));
INVX1 INVX1_493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2785_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2786_));
INVX1 INVX1_494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2789_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2790_));
INVX1 INVX1_495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2794_));
INVX1 INVX1_496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2797_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2798_));
INVX1 INVX1_497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2801_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2802_));
INVX1 INVX1_498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2805_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2806_));
INVX1 INVX1_499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2809_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2810_));
INVX1 INVX1_5 ( .A(inst_r_1_), .Y(_abc_44694_new_n624_));
INVX1 INVX1_50 ( .A(_abc_44694_new_n1080_), .Y(_abc_44694_new_n1081_));
INVX1 INVX1_500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2814_));
INVX1 INVX1_501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2817_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2818_));
INVX1 INVX1_502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2821_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2822_));
INVX1 INVX1_503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2825_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2826_));
INVX1 INVX1_504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2831_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2832_));
INVX1 INVX1_505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2835_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2836_));
INVX1 INVX1_506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2839_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2840_));
INVX1 INVX1_507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2843_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2844_));
INVX1 INVX1_508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2847_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2848_));
INVX1 INVX1_509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2851_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2852_));
INVX1 INVX1_51 ( .A(_abc_44694_new_n1084__bF_buf3), .Y(_abc_44694_new_n1085_));
INVX1 INVX1_510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2855_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2856_));
INVX1 INVX1_511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2859_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2860_));
INVX1 INVX1_512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2863_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2864_));
INVX1 INVX1_513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2867_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2868_));
INVX1 INVX1_514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2871_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2872_));
INVX1 INVX1_515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2875_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2876_));
INVX1 INVX1_516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2879_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2880_));
INVX1 INVX1_517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2883_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2884_));
INVX1 INVX1_518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2887_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2888_));
INVX1 INVX1_519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2892_));
INVX1 INVX1_52 ( .A(opcode_q_22_), .Y(_abc_44694_new_n1094_));
INVX1 INVX1_520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2895_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2896_));
INVX1 INVX1_521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2899_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2900_));
INVX1 INVX1_522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2903_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2904_));
INVX1 INVX1_523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2907_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2908_));
INVX1 INVX1_524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2911_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2912_));
INVX1 INVX1_525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2915_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2916_));
INVX1 INVX1_526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2919_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2920_));
INVX1 INVX1_527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2923_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2924_));
INVX1 INVX1_528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2927_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2928_));
INVX1 INVX1_529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2931_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2932_));
INVX1 INVX1_53 ( .A(opcode_q_21_), .Y(_abc_44694_new_n1095_));
INVX1 INVX1_530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2935_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2936_));
INVX1 INVX1_531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2939_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2940_));
INVX1 INVX1_532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2943_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2944_));
INVX1 INVX1_533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2947_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2948_));
INVX1 INVX1_534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2951_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2952_));
INVX1 INVX1_535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2955_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2956_));
INVX1 INVX1_536 ( .A(REGFILE_SIM_reg_bank_rd_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3056_));
INVX1 INVX1_537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3161_));
INVX1 INVX1_538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3164_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3165_));
INVX1 INVX1_539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3168_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3169_));
INVX1 INVX1_54 ( .A(opcode_q_23_), .Y(_abc_44694_new_n1106_));
INVX1 INVX1_540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3172_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3173_));
INVX1 INVX1_541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3176_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3177_));
INVX1 INVX1_542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3181_));
INVX1 INVX1_543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3184_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3185_));
INVX1 INVX1_544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3188_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3189_));
INVX1 INVX1_545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3192_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3193_));
INVX1 INVX1_546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3196_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3197_));
INVX1 INVX1_547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3201_));
INVX1 INVX1_548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3204_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3205_));
INVX1 INVX1_549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3208_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3209_));
INVX1 INVX1_55 ( .A(_abc_44694_new_n1112_), .Y(_abc_44694_new_n1113_));
INVX1 INVX1_550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3212_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3213_));
INVX1 INVX1_551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3216_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3217_));
INVX1 INVX1_552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3221_));
INVX1 INVX1_553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3224_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3225_));
INVX1 INVX1_554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3228_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3229_));
INVX1 INVX1_555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3232_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3233_));
INVX1 INVX1_556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3236_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3237_));
INVX1 INVX1_557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3241_));
INVX1 INVX1_558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3244_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3245_));
INVX1 INVX1_559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3248_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3249_));
INVX1 INVX1_56 ( .A(_abc_44694_new_n1125_), .Y(_abc_44694_new_n1126_));
INVX1 INVX1_560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3252_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3253_));
INVX1 INVX1_561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3256_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3257_));
INVX1 INVX1_562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3261_));
INVX1 INVX1_563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3264_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3265_));
INVX1 INVX1_564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3268_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3269_));
INVX1 INVX1_565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3272_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3273_));
INVX1 INVX1_566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3276_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3277_));
INVX1 INVX1_567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3280_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3281_));
INVX1 INVX1_568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3284_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3285_));
INVX1 INVX1_569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3290_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3291_));
INVX1 INVX1_57 ( .A(_abc_44694_new_n1128_), .Y(_abc_44694_new_n1129_));
INVX1 INVX1_570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3294_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3295_));
INVX1 INVX1_571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3298_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3299_));
INVX1 INVX1_572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3302_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3303_));
INVX1 INVX1_573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3306_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3307_));
INVX1 INVX1_574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3310_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3311_));
INVX1 INVX1_575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3314_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3315_));
INVX1 INVX1_576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3318_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3319_));
INVX1 INVX1_577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3322_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3323_));
INVX1 INVX1_578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3326_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3327_));
INVX1 INVX1_579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3330_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3331_));
INVX1 INVX1_58 ( .A(_abc_44694_new_n1132_), .Y(_abc_44694_new_n1133_));
INVX1 INVX1_580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3334_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3335_));
INVX1 INVX1_581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3338_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3339_));
INVX1 INVX1_582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3342_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3343_));
INVX1 INVX1_583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3346_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3347_));
INVX1 INVX1_584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3350_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3351_));
INVX1 INVX1_585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3354_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3355_));
INVX1 INVX1_586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3358_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3359_));
INVX1 INVX1_587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3362_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3363_));
INVX1 INVX1_588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3366_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3367_));
INVX1 INVX1_589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3371_));
INVX1 INVX1_59 ( .A(_abc_44694_new_n1136_), .Y(_abc_44694_new_n1137_));
INVX1 INVX1_590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3374_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3375_));
INVX1 INVX1_591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3378_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3379_));
INVX1 INVX1_592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3382_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3383_));
INVX1 INVX1_593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3386_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3387_));
INVX1 INVX1_594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3390_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3391_));
INVX1 INVX1_595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3394_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3395_));
INVX1 INVX1_596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3398_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3399_));
INVX1 INVX1_597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3402_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3403_));
INVX1 INVX1_598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3406_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3407_));
INVX1 INVX1_599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3410_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3411_));
INVX1 INVX1_6 ( .A(inst_r_0_), .Y(_abc_44694_new_n625_));
INVX1 INVX1_60 ( .A(_abc_44694_new_n1162_), .Y(_abc_44694_new_n1163_));
INVX1 INVX1_600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3414_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3415_));
INVX1 INVX1_601 ( .A(REGFILE_SIM_reg_bank_rd_i_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3911_));
INVX1 INVX1_602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3915_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3916_));
INVX1 INVX1_603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3919_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3920_));
INVX1 INVX1_604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3923_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3924_));
INVX1 INVX1_605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3927_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3928_));
INVX1 INVX1_606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3931_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3932_));
INVX1 INVX1_607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3935_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3936_));
INVX1 INVX1_608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3939_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3940_));
INVX1 INVX1_609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3943_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3944_));
INVX1 INVX1_61 ( .A(_abc_44694_new_n1171_), .Y(_abc_44694_new_n1172_));
INVX1 INVX1_610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3947_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3948_));
INVX1 INVX1_611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3951_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3952_));
INVX1 INVX1_612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3955_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3956_));
INVX1 INVX1_613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3959_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3960_));
INVX1 INVX1_614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3963_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3964_));
INVX1 INVX1_615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3967_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3968_));
INVX1 INVX1_616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3971_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3972_));
INVX1 INVX1_617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3975_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3976_));
INVX1 INVX1_618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3979_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3980_));
INVX1 INVX1_619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3983_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3984_));
INVX1 INVX1_62 ( .A(_abc_44694_new_n1173_), .Y(_abc_44694_new_n1174_));
INVX1 INVX1_620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3988_));
INVX1 INVX1_621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3991_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3992_));
INVX1 INVX1_622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3995_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3996_));
INVX1 INVX1_623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3999_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4000_));
INVX1 INVX1_624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4003_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4004_));
INVX1 INVX1_625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4007_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4008_));
INVX1 INVX1_626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4011_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4012_));
INVX1 INVX1_627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4015_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4016_));
INVX1 INVX1_628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4019_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4020_));
INVX1 INVX1_629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4023_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4024_));
INVX1 INVX1_63 ( .A(_abc_44694_new_n1183_), .Y(_abc_44694_new_n1184_));
INVX1 INVX1_630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4027_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4028_));
INVX1 INVX1_631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4031_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4032_));
INVX1 INVX1_632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4035_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4036_));
INVX1 INVX1_633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4039_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4040_));
INVX1 INVX1_634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4437_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4438_));
INVX1 INVX1_635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4442_));
INVX1 INVX1_636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4445_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4446_));
INVX1 INVX1_637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4449_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4450_));
INVX1 INVX1_638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4453_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4454_));
INVX1 INVX1_639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4457_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4458_));
INVX1 INVX1_64 ( .A(_abc_44694_new_n1187_), .Y(_abc_44694_new_n1188_));
INVX1 INVX1_640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4461_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4462_));
INVX1 INVX1_641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4465_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4466_));
INVX1 INVX1_642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4469_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4470_));
INVX1 INVX1_643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4473_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4474_));
INVX1 INVX1_644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4477_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4478_));
INVX1 INVX1_645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4481_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4482_));
INVX1 INVX1_646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4485_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4486_));
INVX1 INVX1_647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4489_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4490_));
INVX1 INVX1_648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4493_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4494_));
INVX1 INVX1_649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4497_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4498_));
INVX1 INVX1_65 ( .A(_abc_44694_new_n1198_), .Y(_abc_44694_new_n1199_));
INVX1 INVX1_650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4501_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4502_));
INVX1 INVX1_651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4505_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4506_));
INVX1 INVX1_652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4509_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4510_));
INVX1 INVX1_653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4513_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4514_));
INVX1 INVX1_654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4518_));
INVX1 INVX1_655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4521_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4522_));
INVX1 INVX1_656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4525_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4526_));
INVX1 INVX1_657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4529_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4530_));
INVX1 INVX1_658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4533_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4534_));
INVX1 INVX1_659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4537_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4538_));
INVX1 INVX1_66 ( .A(_abc_44694_new_n1205_), .Y(_abc_44694_new_n1206_));
INVX1 INVX1_660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4542_));
INVX1 INVX1_661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4545_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4546_));
INVX1 INVX1_662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4550_));
INVX1 INVX1_663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4554_));
INVX1 INVX1_664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4557_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4558_));
INVX1 INVX1_665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4561_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4562_));
INVX1 INVX1_666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4664_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4665_));
INVX1 INVX1_667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4668_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4669_));
INVX1 INVX1_668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4672_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4673_));
INVX1 INVX1_669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4676_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4677_));
INVX1 INVX1_67 ( .A(_abc_44694_new_n1208_), .Y(_abc_44694_new_n1211_));
INVX1 INVX1_670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4680_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4681_));
INVX1 INVX1_671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4684_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4685_));
INVX1 INVX1_672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4688_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4689_));
INVX1 INVX1_673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4692_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4693_));
INVX1 INVX1_674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4696_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4697_));
INVX1 INVX1_675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4700_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4701_));
INVX1 INVX1_676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4704_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4705_));
INVX1 INVX1_677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4708_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4709_));
INVX1 INVX1_678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4712_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4713_));
INVX1 INVX1_679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4716_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4717_));
INVX1 INVX1_68 ( .A(alu_flag_update_o), .Y(_abc_44694_new_n1218_));
INVX1 INVX1_680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4720_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4721_));
INVX1 INVX1_681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4724_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4725_));
INVX1 INVX1_682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4728_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4729_));
INVX1 INVX1_683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4732_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4733_));
INVX1 INVX1_684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4736_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4737_));
INVX1 INVX1_685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4740_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4741_));
INVX1 INVX1_686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4744_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4745_));
INVX1 INVX1_687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4748_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4749_));
INVX1 INVX1_688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4752_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4753_));
INVX1 INVX1_689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4756_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4757_));
INVX1 INVX1_69 ( .A(_abc_44694_new_n1222_), .Y(_abc_44694_new_n1223_));
INVX1 INVX1_690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4760_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4761_));
INVX1 INVX1_691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4764_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4765_));
INVX1 INVX1_692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4768_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4769_));
INVX1 INVX1_693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4772_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4773_));
INVX1 INVX1_694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4776_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4777_));
INVX1 INVX1_695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4780_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4781_));
INVX1 INVX1_696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4784_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4785_));
INVX1 INVX1_697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4788_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4789_));
INVX1 INVX1_698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4989_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4990_));
INVX1 INVX1_699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4993_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4994_));
INVX1 INVX1_7 ( .A(_abc_44694_new_n626_), .Y(_abc_44694_new_n630_));
INVX1 INVX1_70 ( .A(_abc_44694_new_n1099_), .Y(_abc_44694_new_n1226_));
INVX1 INVX1_700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4997_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4998_));
INVX1 INVX1_701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5001_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5002_));
INVX1 INVX1_702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5005_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5006_));
INVX1 INVX1_703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5009_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5010_));
INVX1 INVX1_704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5013_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5014_));
INVX1 INVX1_705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5017_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5018_));
INVX1 INVX1_706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5021_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5022_));
INVX1 INVX1_707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5025_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5026_));
INVX1 INVX1_708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5029_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5030_));
INVX1 INVX1_709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5033_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5034_));
INVX1 INVX1_71 ( .A(alu_less_than_signed_o), .Y(_abc_44694_new_n1230_));
INVX1 INVX1_710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5037_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5038_));
INVX1 INVX1_711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5041_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5042_));
INVX1 INVX1_712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5045_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5046_));
INVX1 INVX1_713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5049_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5050_));
INVX1 INVX1_714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5053_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5054_));
INVX1 INVX1_715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5058_));
INVX1 INVX1_716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5062_));
INVX1 INVX1_717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5065_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5066_));
INVX1 INVX1_718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5069_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5070_));
INVX1 INVX1_719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5073_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5074_));
INVX1 INVX1_72 ( .A(_abc_44694_new_n1231_), .Y(_abc_44694_new_n1232_));
INVX1 INVX1_720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5077_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5078_));
INVX1 INVX1_721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5081_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5082_));
INVX1 INVX1_722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5085_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5086_));
INVX1 INVX1_723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5089_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5090_));
INVX1 INVX1_724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5093_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5094_));
INVX1 INVX1_725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5097_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5098_));
INVX1 INVX1_726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5101_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5102_));
INVX1 INVX1_727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5105_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5106_));
INVX1 INVX1_728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5109_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5110_));
INVX1 INVX1_729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5113_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5114_));
INVX1 INVX1_73 ( .A(alu_equal_o), .Y(_abc_44694_new_n1239_));
INVX1 INVX1_730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5118_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5119_));
INVX1 INVX1_731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5122_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5123_));
INVX1 INVX1_732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5126_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5127_));
INVX1 INVX1_733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5131_));
INVX1 INVX1_734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5134_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5135_));
INVX1 INVX1_735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5138_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5139_));
INVX1 INVX1_736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5143_));
INVX1 INVX1_737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5146_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5147_));
INVX1 INVX1_738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5151_));
INVX1 INVX1_739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5154_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5155_));
INVX1 INVX1_74 ( .A(_abc_44694_new_n1241_), .Y(_abc_44694_new_n1242_));
INVX1 INVX1_740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5159_));
INVX1 INVX1_741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5162_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5163_));
INVX1 INVX1_742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5166_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5167_));
INVX1 INVX1_743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5171_));
INVX1 INVX1_744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5174_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5175_));
INVX1 INVX1_745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5178_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5179_));
INVX1 INVX1_746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5182_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5183_));
INVX1 INVX1_747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5186_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5187_));
INVX1 INVX1_748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5190_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5191_));
INVX1 INVX1_749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5194_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5195_));
INVX1 INVX1_75 ( .A(_abc_44694_new_n1110_), .Y(_abc_44694_new_n1245_));
INVX1 INVX1_750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5198_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5199_));
INVX1 INVX1_751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5202_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5203_));
INVX1 INVX1_752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5206_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5207_));
INVX1 INVX1_753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5211_));
INVX1 INVX1_754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5214_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5215_));
INVX1 INVX1_755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5218_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5219_));
INVX1 INVX1_756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5222_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5223_));
INVX1 INVX1_757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5226_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5227_));
INVX1 INVX1_758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5231_));
INVX1 INVX1_759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5234_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5235_));
INVX1 INVX1_76 ( .A(alu_greater_than_o), .Y(_abc_44694_new_n1246_));
INVX1 INVX1_760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5238_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5239_));
INVX1 INVX1_761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5242_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5243_));
INVX1 INVX1_762 ( .A(REGFILE_SIM_reg_bank_rb_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5545_));
INVX1 INVX1_763 ( .A(REGFILE_SIM_reg_bank_rb_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5551_));
INVX1 INVX1_764 ( .A(REGFILE_SIM_reg_bank_rb_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5562_));
INVX1 INVX1_765 ( .A(REGFILE_SIM_reg_bank_rb_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5579_));
INVX1 INVX1_766 ( .A(REGFILE_SIM_reg_bank_ra_i_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7555_));
INVX1 INVX1_767 ( .A(REGFILE_SIM_reg_bank_ra_i_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7561_));
INVX1 INVX1_768 ( .A(REGFILE_SIM_reg_bank_ra_i_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7572_));
INVX1 INVX1_769 ( .A(REGFILE_SIM_reg_bank_ra_i_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7589_));
INVX1 INVX1_77 ( .A(_abc_44694_new_n1247_), .Y(_abc_44694_new_n1248_));
INVX1 INVX1_770 ( .A(alu__abc_42281_new_n110_), .Y(alu__abc_42281_new_n111_));
INVX1 INVX1_771 ( .A(alu_b_i_20_), .Y(alu__abc_42281_new_n112_));
INVX1 INVX1_772 ( .A(alu_a_i_20_), .Y(alu__abc_42281_new_n113_));
INVX1 INVX1_773 ( .A(alu__abc_42281_new_n114_), .Y(alu__abc_42281_new_n115_));
INVX1 INVX1_774 ( .A(alu__abc_42281_new_n116_), .Y(alu__abc_42281_new_n117_));
INVX1 INVX1_775 ( .A(alu__abc_42281_new_n118_), .Y(alu__abc_42281_new_n119_));
INVX1 INVX1_776 ( .A(alu_b_i_21_), .Y(alu__abc_42281_new_n120_));
INVX1 INVX1_777 ( .A(alu_a_i_21_), .Y(alu__abc_42281_new_n121_));
INVX1 INVX1_778 ( .A(alu__abc_42281_new_n122_), .Y(alu__abc_42281_new_n123_));
INVX1 INVX1_779 ( .A(alu__abc_42281_new_n124_), .Y(alu__abc_42281_new_n125_));
INVX1 INVX1_78 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_9_), .Y(_abc_44694_new_n1271_));
INVX1 INVX1_780 ( .A(alu__abc_42281_new_n127_), .Y(alu__abc_42281_new_n128_));
INVX1 INVX1_781 ( .A(alu_b_i_22_), .Y(alu__abc_42281_new_n129_));
INVX1 INVX1_782 ( .A(alu_a_i_22_), .Y(alu__abc_42281_new_n130_));
INVX1 INVX1_783 ( .A(alu__abc_42281_new_n131_), .Y(alu__abc_42281_new_n132_));
INVX1 INVX1_784 ( .A(alu__abc_42281_new_n133_), .Y(alu__abc_42281_new_n134_));
INVX1 INVX1_785 ( .A(alu__abc_42281_new_n135_), .Y(alu__abc_42281_new_n136_));
INVX1 INVX1_786 ( .A(alu_b_i_23_), .Y(alu__abc_42281_new_n137_));
INVX1 INVX1_787 ( .A(alu_a_i_23_), .Y(alu__abc_42281_new_n138_));
INVX1 INVX1_788 ( .A(alu__abc_42281_new_n139_), .Y(alu__abc_42281_new_n140_));
INVX1 INVX1_789 ( .A(alu__abc_42281_new_n145_), .Y(alu__abc_42281_new_n146_));
INVX1 INVX1_79 ( .A(_abc_44694_new_n1272_), .Y(_abc_44694_new_n1273_));
INVX1 INVX1_790 ( .A(alu_b_i_18_), .Y(alu__abc_42281_new_n147_));
INVX1 INVX1_791 ( .A(alu_a_i_18_), .Y(alu__abc_42281_new_n148_));
INVX1 INVX1_792 ( .A(alu__abc_42281_new_n149_), .Y(alu__abc_42281_new_n150_));
INVX1 INVX1_793 ( .A(alu__abc_42281_new_n151_), .Y(alu__abc_42281_new_n152_));
INVX1 INVX1_794 ( .A(alu__abc_42281_new_n153_), .Y(alu__abc_42281_new_n154_));
INVX1 INVX1_795 ( .A(alu_b_i_19_), .Y(alu__abc_42281_new_n155_));
INVX1 INVX1_796 ( .A(alu_a_i_19_), .Y(alu__abc_42281_new_n156_));
INVX1 INVX1_797 ( .A(alu__abc_42281_new_n157_), .Y(alu__abc_42281_new_n158_));
INVX1 INVX1_798 ( .A(alu__abc_42281_new_n162_), .Y(alu__abc_42281_new_n163_));
INVX1 INVX1_799 ( .A(alu_b_i_16_), .Y(alu__abc_42281_new_n164_));
INVX1 INVX1_8 ( .A(inst_r_3_), .Y(_abc_44694_new_n631_));
INVX1 INVX1_80 ( .A(_abc_44694_new_n1028_), .Y(_abc_44694_new_n1277_));
INVX1 INVX1_800 ( .A(alu_a_i_16_), .Y(alu__abc_42281_new_n165_));
INVX1 INVX1_801 ( .A(alu__abc_42281_new_n166_), .Y(alu__abc_42281_new_n167_));
INVX1 INVX1_802 ( .A(alu__abc_42281_new_n168_), .Y(alu__abc_42281_new_n169_));
INVX1 INVX1_803 ( .A(alu__abc_42281_new_n170_), .Y(alu__abc_42281_new_n171_));
INVX1 INVX1_804 ( .A(alu_b_i_17_), .Y(alu__abc_42281_new_n172_));
INVX1 INVX1_805 ( .A(alu_a_i_17_), .Y(alu__abc_42281_new_n173_));
INVX1 INVX1_806 ( .A(alu__abc_42281_new_n174_), .Y(alu__abc_42281_new_n175_));
INVX1 INVX1_807 ( .A(alu__abc_42281_new_n176_), .Y(alu__abc_42281_new_n177_));
INVX1 INVX1_808 ( .A(alu__abc_42281_new_n181_), .Y(alu__abc_42281_new_n182_));
INVX1 INVX1_809 ( .A(alu_b_i_25_), .Y(alu__abc_42281_new_n183_));
INVX1 INVX1_81 ( .A(_abc_44694_new_n1279_), .Y(_abc_44694_new_n1280_));
INVX1 INVX1_810 ( .A(alu_a_i_25_), .Y(alu__abc_42281_new_n184_));
INVX1 INVX1_811 ( .A(alu__abc_42281_new_n185_), .Y(alu__abc_42281_new_n186_));
INVX1 INVX1_812 ( .A(alu__abc_42281_new_n187_), .Y(alu__abc_42281_new_n188_));
INVX1 INVX1_813 ( .A(alu__abc_42281_new_n189_), .Y(alu__abc_42281_new_n190_));
INVX1 INVX1_814 ( .A(alu_b_i_24_), .Y(alu__abc_42281_new_n191_));
INVX1 INVX1_815 ( .A(alu_a_i_24_), .Y(alu__abc_42281_new_n192_));
INVX1 INVX1_816 ( .A(alu__abc_42281_new_n193_), .Y(alu__abc_42281_new_n194_));
INVX1 INVX1_817 ( .A(alu__abc_42281_new_n195_), .Y(alu__abc_42281_new_n196_));
INVX1 INVX1_818 ( .A(alu__abc_42281_new_n198_), .Y(alu__abc_42281_new_n199_));
INVX1 INVX1_819 ( .A(alu_b_i_26_), .Y(alu__abc_42281_new_n200_));
INVX1 INVX1_82 ( .A(alu_c_update_o), .Y(_abc_44694_new_n1296_));
INVX1 INVX1_820 ( .A(alu_a_i_26_), .Y(alu__abc_42281_new_n201_));
INVX1 INVX1_821 ( .A(alu__abc_42281_new_n202_), .Y(alu__abc_42281_new_n203_));
INVX1 INVX1_822 ( .A(alu__abc_42281_new_n204_), .Y(alu__abc_42281_new_n205_));
INVX1 INVX1_823 ( .A(alu__abc_42281_new_n206_), .Y(alu__abc_42281_new_n207_));
INVX1 INVX1_824 ( .A(alu_b_i_27_), .Y(alu__abc_42281_new_n208_));
INVX1 INVX1_825 ( .A(alu_a_i_27_), .Y(alu__abc_42281_new_n209_));
INVX1 INVX1_826 ( .A(alu__abc_42281_new_n210_), .Y(alu__abc_42281_new_n211_));
INVX1 INVX1_827 ( .A(alu__abc_42281_new_n216_), .Y(alu__abc_42281_new_n217_));
INVX1 INVX1_828 ( .A(alu_b_i_28_), .Y(alu__abc_42281_new_n218_));
INVX1 INVX1_829 ( .A(alu_a_i_28_), .Y(alu__abc_42281_new_n219_));
INVX1 INVX1_83 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_10_), .Y(_abc_44694_new_n1304_));
INVX1 INVX1_830 ( .A(alu__abc_42281_new_n220_), .Y(alu__abc_42281_new_n221_));
INVX1 INVX1_831 ( .A(alu__abc_42281_new_n222_), .Y(alu__abc_42281_new_n223_));
INVX1 INVX1_832 ( .A(alu__abc_42281_new_n224_), .Y(alu__abc_42281_new_n225_));
INVX1 INVX1_833 ( .A(alu_b_i_29_), .Y(alu__abc_42281_new_n226_));
INVX1 INVX1_834 ( .A(alu_a_i_29_), .Y(alu__abc_42281_new_n227_));
INVX1 INVX1_835 ( .A(alu__abc_42281_new_n228_), .Y(alu__abc_42281_new_n229_));
INVX1 INVX1_836 ( .A(alu__abc_42281_new_n230_), .Y(alu__abc_42281_new_n231_));
INVX1 INVX1_837 ( .A(alu__abc_42281_new_n233_), .Y(alu__abc_42281_new_n234_));
INVX1 INVX1_838 ( .A(alu_b_i_30_), .Y(alu__abc_42281_new_n235_));
INVX1 INVX1_839 ( .A(alu_a_i_30_), .Y(alu__abc_42281_new_n236_));
INVX1 INVX1_84 ( .A(_abc_44694_new_n1305_), .Y(_abc_44694_new_n1306_));
INVX1 INVX1_840 ( .A(alu__abc_42281_new_n237_), .Y(alu__abc_42281_new_n238_));
INVX1 INVX1_841 ( .A(alu__abc_42281_new_n239_), .Y(alu__abc_42281_new_n240_));
INVX1 INVX1_842 ( .A(alu_b_i_31_), .Y(alu__abc_42281_new_n242_));
INVX1 INVX1_843 ( .A(alu_a_i_31_), .Y(alu__abc_42281_new_n243_));
INVX1 INVX1_844 ( .A(alu__abc_42281_new_n250_), .Y(alu__abc_42281_new_n251_));
INVX1 INVX1_845 ( .A(alu_b_i_6_), .Y(alu__abc_42281_new_n252_));
INVX1 INVX1_846 ( .A(alu_a_i_6_), .Y(alu__abc_42281_new_n253_));
INVX1 INVX1_847 ( .A(alu__abc_42281_new_n254_), .Y(alu__abc_42281_new_n255_));
INVX1 INVX1_848 ( .A(alu__abc_42281_new_n256_), .Y(alu__abc_42281_new_n257_));
INVX1 INVX1_849 ( .A(alu_b_i_7_), .Y(alu__abc_42281_new_n259_));
INVX1 INVX1_85 ( .A(intr_i), .Y(_abc_44694_new_n1316_));
INVX1 INVX1_850 ( .A(alu_a_i_7_), .Y(alu__abc_42281_new_n260_));
INVX1 INVX1_851 ( .A(alu_b_i_5_), .Y(alu__abc_42281_new_n265_));
INVX1 INVX1_852 ( .A(alu_a_i_5_), .Y(alu__abc_42281_new_n266_));
INVX1 INVX1_853 ( .A(alu__abc_42281_new_n269_), .Y(alu__abc_42281_new_n270_));
INVX1 INVX1_854 ( .A(alu_a_i_4_), .Y(alu__abc_42281_new_n272_));
INVX1 INVX1_855 ( .A(alu__abc_42281_new_n273_), .Y(alu__abc_42281_new_n274_));
INVX1 INVX1_856 ( .A(alu__abc_42281_new_n275_), .Y(alu__abc_42281_new_n276_));
INVX1 INVX1_857 ( .A(alu_a_i_1_), .Y(alu__abc_42281_new_n280_));
INVX1 INVX1_858 ( .A(alu_a_i_0_), .Y(alu__abc_42281_new_n284_));
INVX1 INVX1_859 ( .A(alu__abc_42281_new_n285_), .Y(alu__abc_42281_new_n286_));
INVX1 INVX1_86 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n1350_));
INVX1 INVX1_860 ( .A(alu__abc_42281_new_n289_), .Y(alu__abc_42281_new_n290_));
INVX1 INVX1_861 ( .A(alu_a_i_2_), .Y(alu__abc_42281_new_n293_));
INVX1 INVX1_862 ( .A(alu_a_i_3_), .Y(alu__abc_42281_new_n298_));
INVX1 INVX1_863 ( .A(alu__abc_42281_new_n305_), .Y(alu__abc_42281_new_n306_));
INVX1 INVX1_864 ( .A(alu_b_i_12_), .Y(alu__abc_42281_new_n307_));
INVX1 INVX1_865 ( .A(alu_a_i_12_), .Y(alu__abc_42281_new_n308_));
INVX1 INVX1_866 ( .A(alu__abc_42281_new_n309_), .Y(alu__abc_42281_new_n310_));
INVX1 INVX1_867 ( .A(alu__abc_42281_new_n311_), .Y(alu__abc_42281_new_n312_));
INVX1 INVX1_868 ( .A(alu__abc_42281_new_n313_), .Y(alu__abc_42281_new_n314_));
INVX1 INVX1_869 ( .A(alu_b_i_13_), .Y(alu__abc_42281_new_n315_));
INVX1 INVX1_87 ( .A(_abc_44694_new_n1351_), .Y(_abc_44694_new_n1352_));
INVX1 INVX1_870 ( .A(alu_a_i_13_), .Y(alu__abc_42281_new_n316_));
INVX1 INVX1_871 ( .A(alu__abc_42281_new_n317_), .Y(alu__abc_42281_new_n318_));
INVX1 INVX1_872 ( .A(alu__abc_42281_new_n319_), .Y(alu__abc_42281_new_n320_));
INVX1 INVX1_873 ( .A(alu__abc_42281_new_n322_), .Y(alu__abc_42281_new_n323_));
INVX1 INVX1_874 ( .A(alu_b_i_14_), .Y(alu__abc_42281_new_n324_));
INVX1 INVX1_875 ( .A(alu_a_i_14_), .Y(alu__abc_42281_new_n325_));
INVX1 INVX1_876 ( .A(alu__abc_42281_new_n326_), .Y(alu__abc_42281_new_n327_));
INVX1 INVX1_877 ( .A(alu__abc_42281_new_n328_), .Y(alu__abc_42281_new_n329_));
INVX1 INVX1_878 ( .A(alu__abc_42281_new_n330_), .Y(alu__abc_42281_new_n331_));
INVX1 INVX1_879 ( .A(alu_b_i_15_), .Y(alu__abc_42281_new_n332_));
INVX1 INVX1_88 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n1370_));
INVX1 INVX1_880 ( .A(alu_a_i_15_), .Y(alu__abc_42281_new_n333_));
INVX1 INVX1_881 ( .A(alu__abc_42281_new_n334_), .Y(alu__abc_42281_new_n335_));
INVX1 INVX1_882 ( .A(alu__abc_42281_new_n340_), .Y(alu__abc_42281_new_n341_));
INVX1 INVX1_883 ( .A(alu_b_i_10_), .Y(alu__abc_42281_new_n342_));
INVX1 INVX1_884 ( .A(alu_a_i_10_), .Y(alu__abc_42281_new_n343_));
INVX1 INVX1_885 ( .A(alu__abc_42281_new_n344_), .Y(alu__abc_42281_new_n345_));
INVX1 INVX1_886 ( .A(alu__abc_42281_new_n346_), .Y(alu__abc_42281_new_n347_));
INVX1 INVX1_887 ( .A(alu__abc_42281_new_n348_), .Y(alu__abc_42281_new_n349_));
INVX1 INVX1_888 ( .A(alu_b_i_11_), .Y(alu__abc_42281_new_n350_));
INVX1 INVX1_889 ( .A(alu_a_i_11_), .Y(alu__abc_42281_new_n351_));
INVX1 INVX1_89 ( .A(_abc_44694_new_n1371_), .Y(_abc_44694_new_n1372_));
INVX1 INVX1_890 ( .A(alu__abc_42281_new_n352_), .Y(alu__abc_42281_new_n353_));
INVX1 INVX1_891 ( .A(alu__abc_42281_new_n357_), .Y(alu__abc_42281_new_n358_));
INVX1 INVX1_892 ( .A(alu_b_i_8_), .Y(alu__abc_42281_new_n359_));
INVX1 INVX1_893 ( .A(alu_a_i_8_), .Y(alu__abc_42281_new_n360_));
INVX1 INVX1_894 ( .A(alu__abc_42281_new_n361_), .Y(alu__abc_42281_new_n362_));
INVX1 INVX1_895 ( .A(alu__abc_42281_new_n363_), .Y(alu__abc_42281_new_n364_));
INVX1 INVX1_896 ( .A(alu__abc_42281_new_n365_), .Y(alu__abc_42281_new_n366_));
INVX1 INVX1_897 ( .A(alu_b_i_9_), .Y(alu__abc_42281_new_n367_));
INVX1 INVX1_898 ( .A(alu_a_i_9_), .Y(alu__abc_42281_new_n368_));
INVX1 INVX1_899 ( .A(alu__abc_42281_new_n369_), .Y(alu__abc_42281_new_n370_));
INVX1 INVX1_9 ( .A(_abc_44694_new_n645_), .Y(_abc_44694_new_n646_));
INVX1 INVX1_90 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n1383_));
INVX1 INVX1_900 ( .A(alu__abc_42281_new_n371_), .Y(alu__abc_42281_new_n372_));
INVX1 INVX1_901 ( .A(alu_op_i_1_), .Y(alu__abc_42281_new_n378_));
INVX1 INVX1_902 ( .A(alu_op_i_3_), .Y(alu__abc_42281_new_n379_));
INVX1 INVX1_903 ( .A(alu_op_i_0_), .Y(alu__abc_42281_new_n382_));
INVX1 INVX1_904 ( .A(alu_op_i_2_), .Y(alu__abc_42281_new_n384_));
INVX1 INVX1_905 ( .A(alu__abc_42281_new_n389_), .Y(alu__abc_42281_new_n390_));
INVX1 INVX1_906 ( .A(alu__abc_42281_new_n393_), .Y(alu__abc_42281_new_n394_));
INVX1 INVX1_907 ( .A(alu__abc_42281_new_n397_), .Y(alu__abc_42281_new_n398_));
INVX1 INVX1_908 ( .A(alu__abc_42281_new_n415_), .Y(alu__abc_42281_new_n416_));
INVX1 INVX1_909 ( .A(alu__abc_42281_new_n417_), .Y(alu__abc_42281_new_n418_));
INVX1 INVX1_91 ( .A(_abc_44694_new_n1384_), .Y(_abc_44694_new_n1385_));
INVX1 INVX1_910 ( .A(alu__abc_42281_new_n421_), .Y(alu__abc_42281_new_n422_));
INVX1 INVX1_911 ( .A(alu__abc_42281_new_n430_), .Y(alu__abc_42281_new_n431_));
INVX1 INVX1_912 ( .A(alu__abc_42281_new_n432_), .Y(alu__abc_42281_new_n433_));
INVX1 INVX1_913 ( .A(alu__abc_42281_new_n436_), .Y(alu__abc_42281_new_n437_));
INVX1 INVX1_914 ( .A(alu__abc_42281_new_n447_), .Y(alu__abc_42281_new_n448_));
INVX1 INVX1_915 ( .A(alu__abc_42281_new_n449_), .Y(alu__abc_42281_new_n450_));
INVX1 INVX1_916 ( .A(alu__abc_42281_new_n453_), .Y(alu__abc_42281_new_n454_));
INVX1 INVX1_917 ( .A(alu__abc_42281_new_n462_), .Y(alu__abc_42281_new_n463_));
INVX1 INVX1_918 ( .A(alu__abc_42281_new_n464_), .Y(alu__abc_42281_new_n465_));
INVX1 INVX1_919 ( .A(alu__abc_42281_new_n468_), .Y(alu__abc_42281_new_n469_));
INVX1 INVX1_92 ( .A(_abc_44694_new_n1194__bF_buf1), .Y(_abc_44694_new_n1389_));
INVX1 INVX1_920 ( .A(alu__abc_42281_new_n482_), .Y(alu__abc_42281_new_n483_));
INVX1 INVX1_921 ( .A(alu__abc_42281_new_n214_), .Y(alu__abc_42281_new_n484_));
INVX1 INVX1_922 ( .A(alu__abc_42281_new_n486_), .Y(alu__abc_42281_new_n487_));
INVX1 INVX1_923 ( .A(alu__abc_42281_new_n488_), .Y(alu__abc_42281_new_n489_));
INVX1 INVX1_924 ( .A(alu__abc_42281_new_n493_), .Y(alu__abc_42281_new_n494_));
INVX1 INVX1_925 ( .A(alu__abc_42281_new_n498_), .Y(alu__abc_42281_new_n499_));
INVX1 INVX1_926 ( .A(alu__abc_42281_new_n500_), .Y(alu__abc_42281_new_n501_));
INVX1 INVX1_927 ( .A(alu__abc_42281_new_n503_), .Y(alu__abc_42281_new_n504_));
INVX1 INVX1_928 ( .A(alu__abc_42281_new_n508_), .Y(alu__abc_42281_new_n509_));
INVX1 INVX1_929 ( .A(alu__abc_42281_new_n245_), .Y(alu__abc_42281_new_n512_));
INVX1 INVX1_93 ( .A(_abc_44694_new_n1394_), .Y(_abc_44694_new_n1395_));
INVX1 INVX1_930 ( .A(alu__abc_42281_new_n517_), .Y(alu__abc_42281_new_n518_));
INVX1 INVX1_931 ( .A(alu__abc_42281_new_n521_), .Y(alu__abc_42281_new_n522_));
INVX1 INVX1_932 ( .A(alu__abc_42281_new_n527_), .Y(alu__abc_42281_new_n528_));
INVX1 INVX1_933 ( .A(alu__abc_42281_new_n244_), .Y(alu__abc_42281_new_n530_));
INVX1 INVX1_934 ( .A(alu__abc_42281_new_n540_), .Y(alu__abc_42281_new_n541_));
INVX1 INVX1_935 ( .A(alu__abc_42281_new_n548_), .Y(alu__abc_42281_new_n549_));
INVX1 INVX1_936 ( .A(alu__abc_42281_new_n564_), .Y(alu__abc_42281_new_n565_));
INVX1 INVX1_937 ( .A(alu__abc_42281_new_n279_), .Y(alu__abc_42281_new_n574_));
INVX1 INVX1_938 ( .A(alu__abc_42281_new_n580_), .Y(alu__abc_42281_new_n581_));
INVX1 INVX1_939 ( .A(alu__abc_42281_new_n300_), .Y(alu__abc_42281_new_n583_));
INVX1 INVX1_94 ( .A(_abc_44694_new_n1403_), .Y(_abc_44694_new_n1404_));
INVX1 INVX1_940 ( .A(alu__abc_42281_new_n262_), .Y(alu__abc_42281_new_n587_));
INVX1 INVX1_941 ( .A(alu__abc_42281_new_n268_), .Y(alu__abc_42281_new_n589_));
INVX1 INVX1_942 ( .A(alu__abc_42281_new_n267_), .Y(alu__abc_42281_new_n593_));
INVX1 INVX1_943 ( .A(alu__abc_42281_new_n261_), .Y(alu__abc_42281_new_n597_));
INVX1 INVX1_944 ( .A(alu__abc_42281_new_n622_), .Y(alu__abc_42281_new_n623_));
INVX1 INVX1_945 ( .A(alu__abc_42281_new_n624_), .Y(alu__abc_42281_new_n625_));
INVX1 INVX1_946 ( .A(alu__abc_42281_new_n631_), .Y(alu__abc_42281_new_n632_));
INVX1 INVX1_947 ( .A(alu__abc_42281_new_n633_), .Y(alu__abc_42281_new_n634_));
INVX1 INVX1_948 ( .A(alu__abc_42281_new_n640_), .Y(alu__abc_42281_new_n641_));
INVX1 INVX1_949 ( .A(alu__abc_42281_new_n642_), .Y(alu__abc_42281_new_n643_));
INVX1 INVX1_95 ( .A(pc_q_2_), .Y(_abc_44694_new_n1412_));
INVX1 INVX1_950 ( .A(alu__abc_42281_new_n612_), .Y(alu__abc_42281_new_n648_));
INVX1 INVX1_951 ( .A(alu__abc_42281_new_n652_), .Y(alu__abc_42281_new_n653_));
INVX1 INVX1_952 ( .A(alu__abc_42281_new_n654_), .Y(alu__abc_42281_new_n655_));
INVX1 INVX1_953 ( .A(alu__abc_42281_new_n661_), .Y(alu__abc_42281_new_n662_));
INVX1 INVX1_954 ( .A(alu__abc_42281_new_n667_), .Y(alu__abc_42281_new_n668_));
INVX1 INVX1_955 ( .A(alu__abc_42281_new_n675_), .Y(alu__abc_42281_new_n676_));
INVX1 INVX1_956 ( .A(alu__abc_42281_new_n677_), .Y(alu__abc_42281_new_n678_));
INVX1 INVX1_957 ( .A(alu__abc_42281_new_n684_), .Y(alu__abc_42281_new_n685_));
INVX1 INVX1_958 ( .A(alu__abc_42281_new_n687_), .Y(alu__abc_42281_new_n688_));
INVX1 INVX1_959 ( .A(alu__abc_42281_new_n558_), .Y(alu__abc_42281_new_n693_));
INVX1 INVX1_96 ( .A(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n1424_));
INVX1 INVX1_960 ( .A(alu__abc_42281_new_n570_), .Y(alu__abc_42281_new_n694_));
INVX1 INVX1_961 ( .A(alu__abc_42281_new_n569_), .Y(alu__abc_42281_new_n695_));
INVX1 INVX1_962 ( .A(alu__abc_42281_new_n577_), .Y(alu__abc_42281_new_n696_));
INVX1 INVX1_963 ( .A(alu__abc_42281_new_n585_), .Y(alu__abc_42281_new_n700_));
INVX1 INVX1_964 ( .A(alu__abc_42281_new_n591_), .Y(alu__abc_42281_new_n702_));
INVX1 INVX1_965 ( .A(alu__abc_42281_new_n600_), .Y(alu__abc_42281_new_n704_));
INVX1 INVX1_966 ( .A(alu__abc_42281_new_n603_), .Y(alu__abc_42281_new_n706_));
INVX1 INVX1_967 ( .A(alu__abc_42281_new_n722_), .Y(alu__abc_42281_new_n723_));
INVX1 INVX1_968 ( .A(alu__abc_42281_new_n724_), .Y(alu__abc_42281_new_n725_));
INVX1 INVX1_969 ( .A(alu__abc_42281_new_n730_), .Y(alu__abc_42281_new_n731_));
INVX1 INVX1_97 ( .A(_abc_44694_new_n1425_), .Y(_abc_44694_new_n1426_));
INVX1 INVX1_970 ( .A(alu__abc_42281_new_n734_), .Y(alu__abc_42281_new_n735_));
INVX1 INVX1_971 ( .A(alu__abc_42281_new_n736_), .Y(alu__abc_42281_new_n737_));
INVX1 INVX1_972 ( .A(alu__abc_42281_new_n743_), .Y(alu__abc_42281_new_n744_));
INVX1 INVX1_973 ( .A(alu__abc_42281_new_n745_), .Y(alu__abc_42281_new_n746_));
INVX1 INVX1_974 ( .A(alu__abc_42281_new_n301_), .Y(alu__abc_42281_new_n750_));
INVX1 INVX1_975 ( .A(alu__abc_42281_new_n296_), .Y(alu__abc_42281_new_n751_));
INVX1 INVX1_976 ( .A(alu__abc_42281_new_n753_), .Y(alu__abc_42281_new_n755_));
INVX1 INVX1_977 ( .A(alu__abc_42281_new_n758_), .Y(alu__abc_42281_new_n759_));
INVX1 INVX1_978 ( .A(alu__abc_42281_new_n764_), .Y(alu__abc_42281_new_n765_));
INVX1 INVX1_979 ( .A(alu__abc_42281_new_n602_), .Y(alu__abc_42281_new_n783_));
INVX1 INVX1_98 ( .A(_abc_44694_new_n1431_), .Y(_abc_44694_new_n1432_));
INVX1 INVX1_980 ( .A(alu__abc_42281_new_n816_), .Y(alu__abc_42281_new_n817_));
INVX1 INVX1_981 ( .A(alu__abc_42281_new_n761_), .Y(alu__abc_42281_new_n953_));
INVX1 INVX1_982 ( .A(alu__abc_42281_new_n287_), .Y(alu__abc_42281_new_n1057_));
INVX1 INVX1_983 ( .A(alu__abc_42281_new_n762_), .Y(alu__abc_42281_new_n1069_));
INVX1 INVX1_984 ( .A(alu__abc_42281_new_n766_), .Y(alu__abc_42281_new_n1129_));
INVX1 INVX1_985 ( .A(alu__abc_42281_new_n1135_), .Y(alu__abc_42281_new_n1136_));
INVX1 INVX1_986 ( .A(alu__abc_42281_new_n295_), .Y(alu__abc_42281_new_n1142_));
INVX1 INVX1_987 ( .A(alu__abc_42281_new_n402_), .Y(alu__abc_42281_new_n1152_));
INVX1 INVX1_988 ( .A(alu__abc_42281_new_n767_), .Y(alu__abc_42281_new_n1204_));
INVX1 INVX1_989 ( .A(alu__abc_42281_new_n403_), .Y(alu__abc_42281_new_n1224_));
INVX1 INVX1_99 ( .A(_abc_44694_new_n1435_), .Y(_abc_44694_new_n1436_));
INVX1 INVX1_990 ( .A(alu__abc_42281_new_n770_), .Y(alu__abc_42281_new_n1233_));
INVX1 INVX1_991 ( .A(alu__abc_42281_new_n406_), .Y(alu__abc_42281_new_n1238_));
INVX1 INVX1_992 ( .A(alu__abc_42281_new_n771_), .Y(alu__abc_42281_new_n1286_));
INVX1 INVX1_993 ( .A(alu__abc_42281_new_n407_), .Y(alu__abc_42281_new_n1291_));
INVX1 INVX1_994 ( .A(alu__abc_42281_new_n410_), .Y(alu__abc_42281_new_n1338_));
INVX1 INVX1_995 ( .A(alu__abc_42281_new_n772_), .Y(alu__abc_42281_new_n1341_));
INVX1 INVX1_996 ( .A(alu__abc_42281_new_n411_), .Y(alu__abc_42281_new_n1389_));
INVX1 INVX1_997 ( .A(alu__abc_42281_new_n773_), .Y(alu__abc_42281_new_n1393_));
INVX1 INVX1_998 ( .A(alu__abc_42281_new_n1440_), .Y(alu__abc_42281_new_n1441_));
INVX1 INVX1_999 ( .A(alu__abc_42281_new_n774_), .Y(alu__abc_42281_new_n1445_));
INVX2 INVX2_1 ( .A(_abc_44694_new_n635_), .Y(_abc_44694_new_n636_));
INVX2 INVX2_10 ( .A(alu__abc_42281_new_n212_), .Y(alu__abc_42281_new_n213_));
INVX2 INVX2_11 ( .A(alu__abc_42281_new_n336_), .Y(alu__abc_42281_new_n337_));
INVX2 INVX2_12 ( .A(alu__abc_42281_new_n354_), .Y(alu__abc_42281_new_n355_));
INVX2 INVX2_2 ( .A(_abc_44694_new_n655_), .Y(_abc_44694_new_n667_));
INVX2 INVX2_3 ( .A(_abc_44694_new_n1019__bF_buf3), .Y(_abc_44694_new_n1021_));
INVX2 INVX2_4 ( .A(_abc_44694_new_n1088_), .Y(_abc_44694_new_n1089_));
INVX2 INVX2_5 ( .A(_abc_44694_new_n1114__bF_buf4), .Y(_abc_44694_new_n1115_));
INVX2 INVX2_6 ( .A(_abc_44694_new_n3527__bF_buf4), .Y(_abc_44694_new_n3528_));
INVX2 INVX2_7 ( .A(_abc_44694_new_n4297__bF_buf3), .Y(_abc_44694_new_n4300_));
INVX2 INVX2_8 ( .A(alu__abc_42281_new_n141_), .Y(alu__abc_42281_new_n142_));
INVX2 INVX2_9 ( .A(alu__abc_42281_new_n159_), .Y(alu__abc_42281_new_n160_));
INVX4 INVX4_1 ( .A(state_q_1_bF_buf2_), .Y(_abc_44694_new_n671_));
INVX4 INVX4_10 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2125_));
INVX4 INVX4_11 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2130_));
INVX4 INVX4_12 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2135_));
INVX4 INVX4_13 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2140_));
INVX4 INVX4_14 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2145_));
INVX4 INVX4_15 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2150_));
INVX4 INVX4_16 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2155_));
INVX4 INVX4_17 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2160_));
INVX4 INVX4_18 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2165_));
INVX4 INVX4_19 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2170_));
INVX4 INVX4_2 ( .A(_abc_44694_new_n1185__bF_buf3), .Y(_abc_44694_new_n1186_));
INVX4 INVX4_20 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2175_));
INVX4 INVX4_21 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2180_));
INVX4 INVX4_22 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2185_));
INVX4 INVX4_23 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2190_));
INVX4 INVX4_24 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2195_));
INVX4 INVX4_25 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2200_));
INVX4 INVX4_26 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2205_));
INVX4 INVX4_27 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2210_));
INVX4 INVX4_28 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2215_));
INVX4 INVX4_29 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2220_));
INVX4 INVX4_3 ( .A(_abc_44694_new_n1207__bF_buf0), .Y(_abc_44694_new_n1382_));
INVX4 INVX4_30 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2225_));
INVX4 INVX4_31 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2230_));
INVX4 INVX4_32 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2235_));
INVX4 INVX4_33 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2240_));
INVX4 INVX4_34 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2245_));
INVX4 INVX4_35 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2250_));
INVX4 INVX4_36 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2255_));
INVX4 INVX4_37 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2260_));
INVX4 INVX4_38 ( .A(REGFILE_SIM_reg_bank_rb_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5539_));
INVX4 INVX4_39 ( .A(REGFILE_SIM_reg_bank_ra_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7549_));
INVX4 INVX4_4 ( .A(_abc_44694_new_n1330_), .Y(_abc_44694_new_n1535_));
INVX4 INVX4_5 ( .A(_abc_44694_new_n2834_), .Y(_abc_44694_new_n2835_));
INVX4 INVX4_6 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2105_));
INVX4 INVX4_7 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2110_));
INVX4 INVX4_8 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2115_));
INVX4 INVX4_9 ( .A(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2120_));
INVX8 INVX8_1 ( .A(_abc_44694_new_n644_), .Y(_abc_44694_new_n673_));
INVX8 INVX8_10 ( .A(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3513_));
INVX8 INVX8_11 ( .A(_abc_44694_new_n3518__bF_buf3), .Y(_abc_44694_new_n3519_));
INVX8 INVX8_12 ( .A(_abc_44694_new_n3520__bF_buf4), .Y(_abc_44694_new_n3521_));
INVX8 INVX8_13 ( .A(state_q_5_bF_buf0_), .Y(_abc_44694_new_n3563_));
INVX8 INVX8_14 ( .A(rst_i), .Y(_abc_44694_auto_rtlil_cc_1942_NotGate_34306));
INVX8 INVX8_15 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2269_));
INVX8 INVX8_16 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2370_));
INVX8 INVX8_17 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2602_));
INVX8 INVX8_18 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2960_));
INVX8 INVX8_19 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3061_));
INVX8 INVX8_2 ( .A(_abc_44694_new_n676_), .Y(_abc_44694_new_n677_));
INVX8 INVX8_20 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3419_));
INVX8 INVX8_21 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3519_));
INVX8 INVX8_22 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3618_));
INVX8 INVX8_23 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3717_));
INVX8 INVX8_24 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3815_));
INVX8 INVX8_25 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4044_));
INVX8 INVX8_26 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4142_));
INVX8 INVX8_27 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4241_));
INVX8 INVX8_28 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4339_));
INVX8 INVX8_29 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4566_));
INVX8 INVX8_3 ( .A(_abc_44694_new_n1086_), .Y(_abc_44694_new_n1087_));
INVX8 INVX8_30 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4793_));
INVX8 INVX8_31 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4891_));
INVX8 INVX8_32 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5247_));
INVX8 INVX8_33 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5345_));
INVX8 INVX8_34 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5443_));
INVX8 INVX8_35 ( .A(rst_i), .Y(REGFILE_SIM_reg_bank__abc_34819_auto_rtlil_cc_1942_NotGate_32322));
INVX8 INVX8_36 ( .A(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n271_));
INVX8 INVX8_37 ( .A(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n281_));
INVX8 INVX8_38 ( .A(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n288_));
INVX8 INVX8_39 ( .A(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n294_));
INVX8 INVX8_4 ( .A(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n1179_));
INVX8 INVX8_40 ( .A(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n299_));
INVX8 INVX8_5 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .Y(_abc_44694_new_n1210_));
INVX8 INVX8_6 ( .A(_abc_44694_new_n1278__bF_buf3), .Y(_abc_44694_new_n1334_));
INVX8 INVX8_7 ( .A(_abc_44694_new_n1337__bF_buf3), .Y(_abc_44694_new_n1340_));
INVX8 INVX8_8 ( .A(_abc_44694_new_n1399__bF_buf4), .Y(_abc_44694_new_n1400_));
INVX8 INVX8_9 ( .A(_abc_44694_new_n1348__bF_buf1), .Y(_abc_44694_new_n1522_));
OR2X2 OR2X2_1 ( .A(_abc_44694_new_n641_), .B(_abc_44694_new_n643_), .Y(_abc_44694_new_n644_));
OR2X2 OR2X2_10 ( .A(_abc_44694_new_n686_), .B(_abc_44694_new_n687_), .Y(_abc_44694_new_n688_));
OR2X2 OR2X2_100 ( .A(state_q_1_bF_buf3_), .B(alu_p_o_18_), .Y(_abc_44694_new_n888_));
OR2X2 OR2X2_1000 ( .A(_abc_44694_new_n3310_), .B(_abc_44694_new_n3307_), .Y(alu_func_r_0_));
OR2X2 OR2X2_1001 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1144_), .Y(_abc_44694_new_n3318_));
OR2X2 OR2X2_1002 ( .A(_abc_44694_new_n3318_), .B(_abc_44694_new_n2748_), .Y(_abc_44694_new_n3319_));
OR2X2 OR2X2_1003 ( .A(_abc_44694_new_n3319_), .B(_abc_44694_new_n1182_), .Y(_abc_44694_new_n3320_));
OR2X2 OR2X2_1004 ( .A(_abc_44694_new_n3320_), .B(_abc_44694_new_n1159_), .Y(_abc_44694_new_n3321_));
OR2X2 OR2X2_1005 ( .A(_abc_44694_new_n3321_), .B(_abc_44694_new_n1152_), .Y(_abc_44694_new_n3322_));
OR2X2 OR2X2_1006 ( .A(_abc_44694_new_n3322_), .B(_abc_44694_new_n3317_), .Y(_abc_44694_new_n3323_));
OR2X2 OR2X2_1007 ( .A(_abc_44694_new_n3323_), .B(_abc_44694_new_n3314_), .Y(alu_func_r_1_));
OR2X2 OR2X2_1008 ( .A(_abc_44694_new_n1183_), .B(_abc_44694_new_n1159_), .Y(_abc_44694_new_n3325_));
OR2X2 OR2X2_1009 ( .A(_abc_44694_new_n3325_), .B(_abc_44694_new_n3314_), .Y(_abc_44694_new_n3326_));
OR2X2 OR2X2_101 ( .A(_abc_44694_new_n890_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n891_));
OR2X2 OR2X2_1010 ( .A(_abc_44694_new_n3326_), .B(_abc_44694_new_n1072_), .Y(alu_func_r_2_));
OR2X2 OR2X2_1011 ( .A(_abc_44694_new_n1155_), .B(_abc_44694_new_n1187_), .Y(_abc_44694_new_n3328_));
OR2X2 OR2X2_1012 ( .A(_abc_44694_new_n3328_), .B(_abc_44694_new_n1075_), .Y(_abc_44694_new_n3329_));
OR2X2 OR2X2_1013 ( .A(_abc_44694_new_n2964_), .B(_abc_44694_new_n3329_), .Y(alu_func_r_3_));
OR2X2 OR2X2_1014 ( .A(_abc_44694_new_n3331_), .B(_abc_44694_new_n3334__bF_buf5), .Y(_abc_44694_new_n3335_));
OR2X2 OR2X2_1015 ( .A(_abc_44694_new_n668__bF_buf2), .B(mem_offset_q_0_), .Y(_abc_44694_new_n3336_));
OR2X2 OR2X2_1016 ( .A(_abc_44694_new_n668__bF_buf1), .B(mem_offset_q_1_), .Y(_abc_44694_new_n3338_));
OR2X2 OR2X2_1017 ( .A(_abc_44694_new_n3344_), .B(_abc_44694_new_n3342_), .Y(_abc_44694_new_n3345_));
OR2X2 OR2X2_1018 ( .A(_abc_44694_new_n3331_), .B(_abc_44694_new_n3346_), .Y(_abc_44694_new_n3347_));
OR2X2 OR2X2_1019 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(alu_op_r_0_), .Y(_abc_44694_new_n3350_));
OR2X2 OR2X2_102 ( .A(_abc_44694_new_n892_), .B(_abc_44694_new_n817__bF_buf0), .Y(_abc_44694_new_n893_));
OR2X2 OR2X2_1020 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(alu_op_r_1_), .Y(_abc_44694_new_n3355_));
OR2X2 OR2X2_1021 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(alu_op_r_2_), .Y(_abc_44694_new_n3360_));
OR2X2 OR2X2_1022 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(alu_op_r_3_), .Y(_abc_44694_new_n3365_));
OR2X2 OR2X2_1023 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(int32_r_4_), .Y(_abc_44694_new_n3370_));
OR2X2 OR2X2_1024 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(int32_r_5_), .Y(_abc_44694_new_n3375_));
OR2X2 OR2X2_1025 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(alu_op_r_4_), .Y(_abc_44694_new_n3380_));
OR2X2 OR2X2_1026 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(alu_op_r_5_), .Y(_abc_44694_new_n3385_));
OR2X2 OR2X2_1027 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(alu_op_r_6_), .Y(_abc_44694_new_n3390_));
OR2X2 OR2X2_1028 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(alu_op_r_7_), .Y(_abc_44694_new_n3395_));
OR2X2 OR2X2_1029 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(int32_r_10_), .Y(_abc_44694_new_n3400_));
OR2X2 OR2X2_103 ( .A(state_q_1_bF_buf2_), .B(alu_p_o_19_), .Y(_abc_44694_new_n894_));
OR2X2 OR2X2_1030 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_44694_new_n3405_));
OR2X2 OR2X2_1031 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_44694_new_n3410_));
OR2X2 OR2X2_1032 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_44694_new_n3415_));
OR2X2 OR2X2_1033 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_44694_new_n3420_));
OR2X2 OR2X2_1034 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf4_), .Y(_abc_44694_new_n3425_));
OR2X2 OR2X2_1035 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_44694_new_n3430_));
OR2X2 OR2X2_1036 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_44694_new_n3435_));
OR2X2 OR2X2_1037 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_44694_new_n3440_));
OR2X2 OR2X2_1038 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_44694_new_n3445_));
OR2X2 OR2X2_1039 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf1_), .Y(_abc_44694_new_n3450_));
OR2X2 OR2X2_104 ( .A(_abc_44694_new_n896_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n897_));
OR2X2 OR2X2_1040 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(opcode_q_21_), .Y(_abc_44694_new_n3455_));
OR2X2 OR2X2_1041 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(opcode_q_22_), .Y(_abc_44694_new_n3460_));
OR2X2 OR2X2_1042 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(opcode_q_23_), .Y(_abc_44694_new_n3465_));
OR2X2 OR2X2_1043 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(opcode_q_24_), .Y(_abc_44694_new_n3470_));
OR2X2 OR2X2_1044 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(opcode_q_25_), .Y(_abc_44694_new_n3475_));
OR2X2 OR2X2_1045 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(inst_r_0_), .Y(_abc_44694_new_n3480_));
OR2X2 OR2X2_1046 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(inst_r_1_), .Y(_abc_44694_new_n3485_));
OR2X2 OR2X2_1047 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf7), .B(inst_r_2_), .Y(_abc_44694_new_n3490_));
OR2X2 OR2X2_1048 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf5), .B(inst_r_3_), .Y(_abc_44694_new_n3495_));
OR2X2 OR2X2_1049 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf3), .B(inst_r_4_), .Y(_abc_44694_new_n3500_));
OR2X2 OR2X2_105 ( .A(_abc_44694_new_n898_), .B(_abc_44694_new_n817__bF_buf3), .Y(_abc_44694_new_n899_));
OR2X2 OR2X2_1050 ( .A(_abc_28031_auto_fsm_map_cc_118_implement_pattern_cache_2424_bF_buf1), .B(inst_r_5_), .Y(_abc_44694_new_n3505_));
OR2X2 OR2X2_1051 ( .A(state_q_5_bF_buf1_), .B(_auto_iopadmap_cc_368_execute_48783_0_), .Y(_abc_44694_new_n3510_));
OR2X2 OR2X2_1052 ( .A(_abc_44694_new_n3515__bF_buf3), .B(_abc_44694_new_n3513__bF_buf4), .Y(_abc_44694_new_n3516_));
OR2X2 OR2X2_1053 ( .A(_abc_44694_new_n3516_), .B(_abc_44694_new_n3511_), .Y(_abc_44694_new_n3517_));
OR2X2 OR2X2_1054 ( .A(_abc_44694_new_n3523_), .B(_auto_iopadmap_cc_368_execute_48783_0_), .Y(_abc_44694_new_n3524_));
OR2X2 OR2X2_1055 ( .A(_abc_44694_new_n3528_), .B(_abc_44694_new_n3530_), .Y(_abc_44694_new_n3531_));
OR2X2 OR2X2_1056 ( .A(_abc_44694_new_n3526_), .B(_abc_44694_new_n3531_), .Y(_abc_44694_new_n3532_));
OR2X2 OR2X2_1057 ( .A(_abc_44694_new_n3534_), .B(_auto_iopadmap_cc_368_execute_48783_1_), .Y(_abc_44694_new_n3535_));
OR2X2 OR2X2_1058 ( .A(_abc_44694_new_n3536_), .B(_abc_44694_new_n3518__bF_buf1), .Y(_abc_44694_new_n3537_));
OR2X2 OR2X2_1059 ( .A(_abc_44694_new_n3515__bF_buf2), .B(_abc_44694_new_n3538_), .Y(_abc_44694_new_n3539_));
OR2X2 OR2X2_106 ( .A(state_q_1_bF_buf1_), .B(alu_p_o_20_), .Y(_abc_44694_new_n900_));
OR2X2 OR2X2_1060 ( .A(_abc_44694_new_n3540_), .B(_abc_44694_new_n3528_), .Y(_abc_44694_new_n3541_));
OR2X2 OR2X2_1061 ( .A(state_q_5_bF_buf3_), .B(_auto_iopadmap_cc_368_execute_48783_1_), .Y(_abc_44694_new_n3542_));
OR2X2 OR2X2_1062 ( .A(state_q_5_bF_buf2_), .B(_auto_iopadmap_cc_368_execute_48783_2_), .Y(_abc_44694_new_n3544_));
OR2X2 OR2X2_1063 ( .A(_abc_44694_new_n3546__bF_buf3), .B(_abc_44694_new_n3513__bF_buf2), .Y(_abc_44694_new_n3547_));
OR2X2 OR2X2_1064 ( .A(_abc_44694_new_n3547_), .B(_abc_44694_new_n3545_), .Y(_abc_44694_new_n3548_));
OR2X2 OR2X2_1065 ( .A(_abc_44694_new_n3523_), .B(_auto_iopadmap_cc_368_execute_48783_2_), .Y(_abc_44694_new_n3549_));
OR2X2 OR2X2_1066 ( .A(_abc_44694_new_n3528_), .B(_abc_44694_new_n3552_), .Y(_abc_44694_new_n3553_));
OR2X2 OR2X2_1067 ( .A(_abc_44694_new_n3551_), .B(_abc_44694_new_n3553_), .Y(_abc_44694_new_n3554_));
OR2X2 OR2X2_1068 ( .A(_abc_44694_new_n3556_), .B(_auto_iopadmap_cc_368_execute_48783_3_), .Y(_abc_44694_new_n3557_));
OR2X2 OR2X2_1069 ( .A(_abc_44694_new_n3546__bF_buf2), .B(_abc_44694_new_n3538_), .Y(_abc_44694_new_n3558_));
OR2X2 OR2X2_107 ( .A(_abc_44694_new_n902_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n903_));
OR2X2 OR2X2_1070 ( .A(_abc_44694_new_n3559_), .B(_abc_44694_new_n3528_), .Y(_abc_44694_new_n3560_));
OR2X2 OR2X2_1071 ( .A(state_q_5_bF_buf1_), .B(_auto_iopadmap_cc_368_execute_48783_3_), .Y(_abc_44694_new_n3561_));
OR2X2 OR2X2_1072 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n3567_), .Y(_abc_44694_new_n3568_));
OR2X2 OR2X2_1073 ( .A(_abc_44694_new_n3566_), .B(_abc_44694_new_n3568_), .Y(_abc_44694_new_n3569_));
OR2X2 OR2X2_1074 ( .A(_abc_44694_new_n3571_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n3572_));
OR2X2 OR2X2_1075 ( .A(_abc_44694_new_n3572_), .B(_abc_44694_new_n3570_), .Y(_abc_44694_new_n3573_));
OR2X2 OR2X2_1076 ( .A(_abc_44694_new_n3575_), .B(_abc_44694_new_n3565_), .Y(_abc_44694_new_n3576_));
OR2X2 OR2X2_1077 ( .A(_abc_44694_new_n3577_), .B(_abc_44694_new_n3564_), .Y(_0mem_dat_o_31_0__0_));
OR2X2 OR2X2_1078 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n3582_), .Y(_abc_44694_new_n3583_));
OR2X2 OR2X2_1079 ( .A(_abc_44694_new_n3581_), .B(_abc_44694_new_n3583_), .Y(_abc_44694_new_n3584_));
OR2X2 OR2X2_108 ( .A(_abc_44694_new_n904_), .B(_abc_44694_new_n817__bF_buf2), .Y(_abc_44694_new_n905_));
OR2X2 OR2X2_1080 ( .A(_abc_44694_new_n3586_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n3587_));
OR2X2 OR2X2_1081 ( .A(_abc_44694_new_n3587_), .B(_abc_44694_new_n3585_), .Y(_abc_44694_new_n3588_));
OR2X2 OR2X2_1082 ( .A(_abc_44694_new_n3590_), .B(_abc_44694_new_n3580_), .Y(_abc_44694_new_n3591_));
OR2X2 OR2X2_1083 ( .A(_abc_44694_new_n3592_), .B(_abc_44694_new_n3579_), .Y(_0mem_dat_o_31_0__1_));
OR2X2 OR2X2_1084 ( .A(_abc_44694_new_n3513__bF_buf4), .B(_abc_44694_new_n3597_), .Y(_abc_44694_new_n3598_));
OR2X2 OR2X2_1085 ( .A(_abc_44694_new_n3596_), .B(_abc_44694_new_n3598_), .Y(_abc_44694_new_n3599_));
OR2X2 OR2X2_1086 ( .A(_abc_44694_new_n3601_), .B(_abc_44694_new_n3512__bF_buf0), .Y(_abc_44694_new_n3602_));
OR2X2 OR2X2_1087 ( .A(_abc_44694_new_n3602_), .B(_abc_44694_new_n3600_), .Y(_abc_44694_new_n3603_));
OR2X2 OR2X2_1088 ( .A(_abc_44694_new_n3605_), .B(_abc_44694_new_n3595_), .Y(_abc_44694_new_n3606_));
OR2X2 OR2X2_1089 ( .A(_abc_44694_new_n3607_), .B(_abc_44694_new_n3594_), .Y(_0mem_dat_o_31_0__2_));
OR2X2 OR2X2_109 ( .A(state_q_1_bF_buf0_), .B(alu_p_o_21_), .Y(_abc_44694_new_n906_));
OR2X2 OR2X2_1090 ( .A(_abc_44694_new_n3513__bF_buf3), .B(_abc_44694_new_n3612_), .Y(_abc_44694_new_n3613_));
OR2X2 OR2X2_1091 ( .A(_abc_44694_new_n3611_), .B(_abc_44694_new_n3613_), .Y(_abc_44694_new_n3614_));
OR2X2 OR2X2_1092 ( .A(_abc_44694_new_n3616_), .B(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3617_));
OR2X2 OR2X2_1093 ( .A(_abc_44694_new_n3617_), .B(_abc_44694_new_n3615_), .Y(_abc_44694_new_n3618_));
OR2X2 OR2X2_1094 ( .A(_abc_44694_new_n3620_), .B(_abc_44694_new_n3610_), .Y(_abc_44694_new_n3621_));
OR2X2 OR2X2_1095 ( .A(_abc_44694_new_n3622_), .B(_abc_44694_new_n3609_), .Y(_0mem_dat_o_31_0__3_));
OR2X2 OR2X2_1096 ( .A(_abc_44694_new_n3513__bF_buf2), .B(_abc_44694_new_n3627_), .Y(_abc_44694_new_n3628_));
OR2X2 OR2X2_1097 ( .A(_abc_44694_new_n3626_), .B(_abc_44694_new_n3628_), .Y(_abc_44694_new_n3629_));
OR2X2 OR2X2_1098 ( .A(_abc_44694_new_n3631_), .B(_abc_44694_new_n3512__bF_buf3), .Y(_abc_44694_new_n3632_));
OR2X2 OR2X2_1099 ( .A(_abc_44694_new_n3632_), .B(_abc_44694_new_n3630_), .Y(_abc_44694_new_n3633_));
OR2X2 OR2X2_11 ( .A(_abc_44694_new_n690_), .B(_abc_44694_new_n692_), .Y(_abc_44694_new_n693_));
OR2X2 OR2X2_110 ( .A(_abc_44694_new_n908_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n909_));
OR2X2 OR2X2_1100 ( .A(_abc_44694_new_n3635_), .B(_abc_44694_new_n3625_), .Y(_abc_44694_new_n3636_));
OR2X2 OR2X2_1101 ( .A(_abc_44694_new_n3637_), .B(_abc_44694_new_n3624_), .Y(_0mem_dat_o_31_0__4_));
OR2X2 OR2X2_1102 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n3642_), .Y(_abc_44694_new_n3643_));
OR2X2 OR2X2_1103 ( .A(_abc_44694_new_n3641_), .B(_abc_44694_new_n3643_), .Y(_abc_44694_new_n3644_));
OR2X2 OR2X2_1104 ( .A(_abc_44694_new_n3646_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n3647_));
OR2X2 OR2X2_1105 ( .A(_abc_44694_new_n3647_), .B(_abc_44694_new_n3645_), .Y(_abc_44694_new_n3648_));
OR2X2 OR2X2_1106 ( .A(_abc_44694_new_n3650_), .B(_abc_44694_new_n3640_), .Y(_abc_44694_new_n3651_));
OR2X2 OR2X2_1107 ( .A(_abc_44694_new_n3652_), .B(_abc_44694_new_n3639_), .Y(_0mem_dat_o_31_0__5_));
OR2X2 OR2X2_1108 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n3657_), .Y(_abc_44694_new_n3658_));
OR2X2 OR2X2_1109 ( .A(_abc_44694_new_n3656_), .B(_abc_44694_new_n3658_), .Y(_abc_44694_new_n3659_));
OR2X2 OR2X2_111 ( .A(_abc_44694_new_n910_), .B(_abc_44694_new_n817__bF_buf1), .Y(_abc_44694_new_n911_));
OR2X2 OR2X2_1110 ( .A(_abc_44694_new_n3661_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n3662_));
OR2X2 OR2X2_1111 ( .A(_abc_44694_new_n3662_), .B(_abc_44694_new_n3660_), .Y(_abc_44694_new_n3663_));
OR2X2 OR2X2_1112 ( .A(_abc_44694_new_n3665_), .B(_abc_44694_new_n3655_), .Y(_abc_44694_new_n3666_));
OR2X2 OR2X2_1113 ( .A(_abc_44694_new_n3667_), .B(_abc_44694_new_n3654_), .Y(_0mem_dat_o_31_0__6_));
OR2X2 OR2X2_1114 ( .A(_abc_44694_new_n3513__bF_buf4), .B(_abc_44694_new_n3672_), .Y(_abc_44694_new_n3673_));
OR2X2 OR2X2_1115 ( .A(_abc_44694_new_n3671_), .B(_abc_44694_new_n3673_), .Y(_abc_44694_new_n3674_));
OR2X2 OR2X2_1116 ( .A(_abc_44694_new_n3676_), .B(_abc_44694_new_n3512__bF_buf0), .Y(_abc_44694_new_n3677_));
OR2X2 OR2X2_1117 ( .A(_abc_44694_new_n3677_), .B(_abc_44694_new_n3675_), .Y(_abc_44694_new_n3678_));
OR2X2 OR2X2_1118 ( .A(_abc_44694_new_n3680_), .B(_abc_44694_new_n3670_), .Y(_abc_44694_new_n3681_));
OR2X2 OR2X2_1119 ( .A(_abc_44694_new_n3682_), .B(_abc_44694_new_n3669_), .Y(_0mem_dat_o_31_0__7_));
OR2X2 OR2X2_112 ( .A(state_q_1_bF_buf4_), .B(alu_p_o_22_), .Y(_abc_44694_new_n912_));
OR2X2 OR2X2_1120 ( .A(_abc_44694_new_n3685_), .B(_abc_44694_new_n3686_), .Y(_abc_44694_new_n3687_));
OR2X2 OR2X2_1121 ( .A(_abc_44694_new_n3687_), .B(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3688_));
OR2X2 OR2X2_1122 ( .A(_abc_44694_new_n3513__bF_buf3), .B(_abc_44694_new_n3690_), .Y(_abc_44694_new_n3691_));
OR2X2 OR2X2_1123 ( .A(_abc_44694_new_n3689_), .B(_abc_44694_new_n3691_), .Y(_abc_44694_new_n3692_));
OR2X2 OR2X2_1124 ( .A(_abc_44694_new_n3693_), .B(_abc_44694_new_n3518__bF_buf0), .Y(_abc_44694_new_n3694_));
OR2X2 OR2X2_1125 ( .A(_abc_44694_new_n3566_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3695_));
OR2X2 OR2X2_1126 ( .A(_abc_44694_new_n3697_), .B(_abc_44694_new_n3684_), .Y(_0mem_dat_o_31_0__8_));
OR2X2 OR2X2_1127 ( .A(_abc_44694_new_n3700_), .B(_abc_44694_new_n3701_), .Y(_abc_44694_new_n3702_));
OR2X2 OR2X2_1128 ( .A(_abc_44694_new_n3702_), .B(_abc_44694_new_n3512__bF_buf3), .Y(_abc_44694_new_n3703_));
OR2X2 OR2X2_1129 ( .A(_abc_44694_new_n3513__bF_buf2), .B(_abc_44694_new_n3705_), .Y(_abc_44694_new_n3706_));
OR2X2 OR2X2_113 ( .A(_abc_44694_new_n914_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n915_));
OR2X2 OR2X2_1130 ( .A(_abc_44694_new_n3704_), .B(_abc_44694_new_n3706_), .Y(_abc_44694_new_n3707_));
OR2X2 OR2X2_1131 ( .A(_abc_44694_new_n3708_), .B(_abc_44694_new_n3518__bF_buf3), .Y(_abc_44694_new_n3709_));
OR2X2 OR2X2_1132 ( .A(_abc_44694_new_n3581_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n3710_));
OR2X2 OR2X2_1133 ( .A(_abc_44694_new_n3712_), .B(_abc_44694_new_n3699_), .Y(_0mem_dat_o_31_0__9_));
OR2X2 OR2X2_1134 ( .A(_abc_44694_new_n3715_), .B(_abc_44694_new_n3716_), .Y(_abc_44694_new_n3717_));
OR2X2 OR2X2_1135 ( .A(_abc_44694_new_n3717_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n3718_));
OR2X2 OR2X2_1136 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n3720_), .Y(_abc_44694_new_n3721_));
OR2X2 OR2X2_1137 ( .A(_abc_44694_new_n3719_), .B(_abc_44694_new_n3721_), .Y(_abc_44694_new_n3722_));
OR2X2 OR2X2_1138 ( .A(_abc_44694_new_n3723_), .B(_abc_44694_new_n3518__bF_buf2), .Y(_abc_44694_new_n3724_));
OR2X2 OR2X2_1139 ( .A(_abc_44694_new_n3596_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n3725_));
OR2X2 OR2X2_114 ( .A(_abc_44694_new_n916_), .B(_abc_44694_new_n817__bF_buf0), .Y(_abc_44694_new_n917_));
OR2X2 OR2X2_1140 ( .A(_abc_44694_new_n3727_), .B(_abc_44694_new_n3714_), .Y(_0mem_dat_o_31_0__10_));
OR2X2 OR2X2_1141 ( .A(_abc_44694_new_n3730_), .B(_abc_44694_new_n3731_), .Y(_abc_44694_new_n3732_));
OR2X2 OR2X2_1142 ( .A(_abc_44694_new_n3732_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n3733_));
OR2X2 OR2X2_1143 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n3735_), .Y(_abc_44694_new_n3736_));
OR2X2 OR2X2_1144 ( .A(_abc_44694_new_n3734_), .B(_abc_44694_new_n3736_), .Y(_abc_44694_new_n3737_));
OR2X2 OR2X2_1145 ( .A(_abc_44694_new_n3738_), .B(_abc_44694_new_n3518__bF_buf1), .Y(_abc_44694_new_n3739_));
OR2X2 OR2X2_1146 ( .A(_abc_44694_new_n3611_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n3740_));
OR2X2 OR2X2_1147 ( .A(_abc_44694_new_n3742_), .B(_abc_44694_new_n3729_), .Y(_0mem_dat_o_31_0__11_));
OR2X2 OR2X2_1148 ( .A(_abc_44694_new_n3745_), .B(_abc_44694_new_n3746_), .Y(_abc_44694_new_n3747_));
OR2X2 OR2X2_1149 ( .A(_abc_44694_new_n3747_), .B(_abc_44694_new_n3512__bF_buf0), .Y(_abc_44694_new_n3748_));
OR2X2 OR2X2_115 ( .A(state_q_1_bF_buf3_), .B(alu_p_o_23_), .Y(_abc_44694_new_n918_));
OR2X2 OR2X2_1150 ( .A(_abc_44694_new_n3513__bF_buf4), .B(_abc_44694_new_n3750_), .Y(_abc_44694_new_n3751_));
OR2X2 OR2X2_1151 ( .A(_abc_44694_new_n3749_), .B(_abc_44694_new_n3751_), .Y(_abc_44694_new_n3752_));
OR2X2 OR2X2_1152 ( .A(_abc_44694_new_n3753_), .B(_abc_44694_new_n3518__bF_buf0), .Y(_abc_44694_new_n3754_));
OR2X2 OR2X2_1153 ( .A(_abc_44694_new_n3626_), .B(_abc_44694_new_n3519__bF_buf0), .Y(_abc_44694_new_n3755_));
OR2X2 OR2X2_1154 ( .A(_abc_44694_new_n3757_), .B(_abc_44694_new_n3744_), .Y(_0mem_dat_o_31_0__12_));
OR2X2 OR2X2_1155 ( .A(_abc_44694_new_n3760_), .B(_abc_44694_new_n3761_), .Y(_abc_44694_new_n3762_));
OR2X2 OR2X2_1156 ( .A(_abc_44694_new_n3762_), .B(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3763_));
OR2X2 OR2X2_1157 ( .A(_abc_44694_new_n3513__bF_buf3), .B(_abc_44694_new_n3765_), .Y(_abc_44694_new_n3766_));
OR2X2 OR2X2_1158 ( .A(_abc_44694_new_n3764_), .B(_abc_44694_new_n3766_), .Y(_abc_44694_new_n3767_));
OR2X2 OR2X2_1159 ( .A(_abc_44694_new_n3768_), .B(_abc_44694_new_n3518__bF_buf3), .Y(_abc_44694_new_n3769_));
OR2X2 OR2X2_116 ( .A(_abc_44694_new_n920_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n921_));
OR2X2 OR2X2_1160 ( .A(_abc_44694_new_n3641_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3770_));
OR2X2 OR2X2_1161 ( .A(_abc_44694_new_n3772_), .B(_abc_44694_new_n3759_), .Y(_0mem_dat_o_31_0__13_));
OR2X2 OR2X2_1162 ( .A(_abc_44694_new_n3775_), .B(_abc_44694_new_n3776_), .Y(_abc_44694_new_n3777_));
OR2X2 OR2X2_1163 ( .A(_abc_44694_new_n3777_), .B(_abc_44694_new_n3512__bF_buf3), .Y(_abc_44694_new_n3778_));
OR2X2 OR2X2_1164 ( .A(_abc_44694_new_n3513__bF_buf2), .B(_abc_44694_new_n3780_), .Y(_abc_44694_new_n3781_));
OR2X2 OR2X2_1165 ( .A(_abc_44694_new_n3779_), .B(_abc_44694_new_n3781_), .Y(_abc_44694_new_n3782_));
OR2X2 OR2X2_1166 ( .A(_abc_44694_new_n3783_), .B(_abc_44694_new_n3518__bF_buf2), .Y(_abc_44694_new_n3784_));
OR2X2 OR2X2_1167 ( .A(_abc_44694_new_n3656_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n3785_));
OR2X2 OR2X2_1168 ( .A(_abc_44694_new_n3787_), .B(_abc_44694_new_n3774_), .Y(_0mem_dat_o_31_0__14_));
OR2X2 OR2X2_1169 ( .A(_abc_44694_new_n3790_), .B(_abc_44694_new_n3791_), .Y(_abc_44694_new_n3792_));
OR2X2 OR2X2_117 ( .A(_abc_44694_new_n922_), .B(_abc_44694_new_n817__bF_buf3), .Y(_abc_44694_new_n923_));
OR2X2 OR2X2_1170 ( .A(_abc_44694_new_n3792_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n3793_));
OR2X2 OR2X2_1171 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n3795_), .Y(_abc_44694_new_n3796_));
OR2X2 OR2X2_1172 ( .A(_abc_44694_new_n3794_), .B(_abc_44694_new_n3796_), .Y(_abc_44694_new_n3797_));
OR2X2 OR2X2_1173 ( .A(_abc_44694_new_n3798_), .B(_abc_44694_new_n3518__bF_buf1), .Y(_abc_44694_new_n3799_));
OR2X2 OR2X2_1174 ( .A(_abc_44694_new_n3671_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n3800_));
OR2X2 OR2X2_1175 ( .A(_abc_44694_new_n3802_), .B(_abc_44694_new_n3789_), .Y(_0mem_dat_o_31_0__15_));
OR2X2 OR2X2_1176 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n3807_), .Y(_abc_44694_new_n3808_));
OR2X2 OR2X2_1177 ( .A(_abc_44694_new_n3806_), .B(_abc_44694_new_n3808_), .Y(_abc_44694_new_n3809_));
OR2X2 OR2X2_1178 ( .A(_abc_44694_new_n3811_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n3812_));
OR2X2 OR2X2_1179 ( .A(_abc_44694_new_n3812_), .B(_abc_44694_new_n3810_), .Y(_abc_44694_new_n3813_));
OR2X2 OR2X2_118 ( .A(state_q_1_bF_buf2_), .B(alu_p_o_24_), .Y(_abc_44694_new_n924_));
OR2X2 OR2X2_1180 ( .A(_abc_44694_new_n3815_), .B(_abc_44694_new_n3805_), .Y(_abc_44694_new_n3816_));
OR2X2 OR2X2_1181 ( .A(_abc_44694_new_n3817_), .B(_abc_44694_new_n3804_), .Y(_0mem_dat_o_31_0__16_));
OR2X2 OR2X2_1182 ( .A(_abc_44694_new_n3513__bF_buf4), .B(_abc_44694_new_n3822_), .Y(_abc_44694_new_n3823_));
OR2X2 OR2X2_1183 ( .A(_abc_44694_new_n3821_), .B(_abc_44694_new_n3823_), .Y(_abc_44694_new_n3824_));
OR2X2 OR2X2_1184 ( .A(_abc_44694_new_n3826_), .B(_abc_44694_new_n3512__bF_buf0), .Y(_abc_44694_new_n3827_));
OR2X2 OR2X2_1185 ( .A(_abc_44694_new_n3827_), .B(_abc_44694_new_n3825_), .Y(_abc_44694_new_n3828_));
OR2X2 OR2X2_1186 ( .A(_abc_44694_new_n3830_), .B(_abc_44694_new_n3820_), .Y(_abc_44694_new_n3831_));
OR2X2 OR2X2_1187 ( .A(_abc_44694_new_n3832_), .B(_abc_44694_new_n3819_), .Y(_0mem_dat_o_31_0__17_));
OR2X2 OR2X2_1188 ( .A(_abc_44694_new_n3513__bF_buf3), .B(_abc_44694_new_n3837_), .Y(_abc_44694_new_n3838_));
OR2X2 OR2X2_1189 ( .A(_abc_44694_new_n3836_), .B(_abc_44694_new_n3838_), .Y(_abc_44694_new_n3839_));
OR2X2 OR2X2_119 ( .A(_abc_44694_new_n926_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n927_));
OR2X2 OR2X2_1190 ( .A(_abc_44694_new_n3841_), .B(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3842_));
OR2X2 OR2X2_1191 ( .A(_abc_44694_new_n3842_), .B(_abc_44694_new_n3840_), .Y(_abc_44694_new_n3843_));
OR2X2 OR2X2_1192 ( .A(_abc_44694_new_n3845_), .B(_abc_44694_new_n3835_), .Y(_abc_44694_new_n3846_));
OR2X2 OR2X2_1193 ( .A(_abc_44694_new_n3847_), .B(_abc_44694_new_n3834_), .Y(_0mem_dat_o_31_0__18_));
OR2X2 OR2X2_1194 ( .A(_abc_44694_new_n3513__bF_buf2), .B(_abc_44694_new_n3852_), .Y(_abc_44694_new_n3853_));
OR2X2 OR2X2_1195 ( .A(_abc_44694_new_n3851_), .B(_abc_44694_new_n3853_), .Y(_abc_44694_new_n3854_));
OR2X2 OR2X2_1196 ( .A(_abc_44694_new_n3856_), .B(_abc_44694_new_n3512__bF_buf3), .Y(_abc_44694_new_n3857_));
OR2X2 OR2X2_1197 ( .A(_abc_44694_new_n3857_), .B(_abc_44694_new_n3855_), .Y(_abc_44694_new_n3858_));
OR2X2 OR2X2_1198 ( .A(_abc_44694_new_n3860_), .B(_abc_44694_new_n3850_), .Y(_abc_44694_new_n3861_));
OR2X2 OR2X2_1199 ( .A(_abc_44694_new_n3862_), .B(_abc_44694_new_n3849_), .Y(_0mem_dat_o_31_0__19_));
OR2X2 OR2X2_12 ( .A(_abc_44694_new_n688_), .B(_abc_44694_new_n693_), .Y(_abc_44694_new_n694_));
OR2X2 OR2X2_120 ( .A(_abc_44694_new_n928_), .B(_abc_44694_new_n817__bF_buf2), .Y(_abc_44694_new_n929_));
OR2X2 OR2X2_1200 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n3867_), .Y(_abc_44694_new_n3868_));
OR2X2 OR2X2_1201 ( .A(_abc_44694_new_n3866_), .B(_abc_44694_new_n3868_), .Y(_abc_44694_new_n3869_));
OR2X2 OR2X2_1202 ( .A(_abc_44694_new_n3871_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n3872_));
OR2X2 OR2X2_1203 ( .A(_abc_44694_new_n3872_), .B(_abc_44694_new_n3870_), .Y(_abc_44694_new_n3873_));
OR2X2 OR2X2_1204 ( .A(_abc_44694_new_n3875_), .B(_abc_44694_new_n3865_), .Y(_abc_44694_new_n3876_));
OR2X2 OR2X2_1205 ( .A(_abc_44694_new_n3877_), .B(_abc_44694_new_n3864_), .Y(_0mem_dat_o_31_0__20_));
OR2X2 OR2X2_1206 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n3882_), .Y(_abc_44694_new_n3883_));
OR2X2 OR2X2_1207 ( .A(_abc_44694_new_n3881_), .B(_abc_44694_new_n3883_), .Y(_abc_44694_new_n3884_));
OR2X2 OR2X2_1208 ( .A(_abc_44694_new_n3886_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n3887_));
OR2X2 OR2X2_1209 ( .A(_abc_44694_new_n3887_), .B(_abc_44694_new_n3885_), .Y(_abc_44694_new_n3888_));
OR2X2 OR2X2_121 ( .A(state_q_1_bF_buf1_), .B(alu_p_o_25_), .Y(_abc_44694_new_n930_));
OR2X2 OR2X2_1210 ( .A(_abc_44694_new_n3890_), .B(_abc_44694_new_n3880_), .Y(_abc_44694_new_n3891_));
OR2X2 OR2X2_1211 ( .A(_abc_44694_new_n3892_), .B(_abc_44694_new_n3879_), .Y(_0mem_dat_o_31_0__21_));
OR2X2 OR2X2_1212 ( .A(_abc_44694_new_n3513__bF_buf4), .B(_abc_44694_new_n3897_), .Y(_abc_44694_new_n3898_));
OR2X2 OR2X2_1213 ( .A(_abc_44694_new_n3896_), .B(_abc_44694_new_n3898_), .Y(_abc_44694_new_n3899_));
OR2X2 OR2X2_1214 ( .A(_abc_44694_new_n3901_), .B(_abc_44694_new_n3512__bF_buf0), .Y(_abc_44694_new_n3902_));
OR2X2 OR2X2_1215 ( .A(_abc_44694_new_n3902_), .B(_abc_44694_new_n3900_), .Y(_abc_44694_new_n3903_));
OR2X2 OR2X2_1216 ( .A(_abc_44694_new_n3905_), .B(_abc_44694_new_n3895_), .Y(_abc_44694_new_n3906_));
OR2X2 OR2X2_1217 ( .A(_abc_44694_new_n3907_), .B(_abc_44694_new_n3894_), .Y(_0mem_dat_o_31_0__22_));
OR2X2 OR2X2_1218 ( .A(_abc_44694_new_n3513__bF_buf3), .B(_abc_44694_new_n3912_), .Y(_abc_44694_new_n3913_));
OR2X2 OR2X2_1219 ( .A(_abc_44694_new_n3911_), .B(_abc_44694_new_n3913_), .Y(_abc_44694_new_n3914_));
OR2X2 OR2X2_122 ( .A(_abc_44694_new_n932_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n933_));
OR2X2 OR2X2_1220 ( .A(_abc_44694_new_n3916_), .B(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3917_));
OR2X2 OR2X2_1221 ( .A(_abc_44694_new_n3917_), .B(_abc_44694_new_n3915_), .Y(_abc_44694_new_n3918_));
OR2X2 OR2X2_1222 ( .A(_abc_44694_new_n3920_), .B(_abc_44694_new_n3910_), .Y(_abc_44694_new_n3921_));
OR2X2 OR2X2_1223 ( .A(_abc_44694_new_n3922_), .B(_abc_44694_new_n3909_), .Y(_0mem_dat_o_31_0__23_));
OR2X2 OR2X2_1224 ( .A(_abc_44694_new_n3925_), .B(_abc_44694_new_n3926_), .Y(_abc_44694_new_n3927_));
OR2X2 OR2X2_1225 ( .A(_abc_44694_new_n3927_), .B(_abc_44694_new_n3512__bF_buf3), .Y(_abc_44694_new_n3928_));
OR2X2 OR2X2_1226 ( .A(_abc_44694_new_n3513__bF_buf2), .B(_abc_44694_new_n3930_), .Y(_abc_44694_new_n3931_));
OR2X2 OR2X2_1227 ( .A(_abc_44694_new_n3929_), .B(_abc_44694_new_n3931_), .Y(_abc_44694_new_n3932_));
OR2X2 OR2X2_1228 ( .A(_abc_44694_new_n3933_), .B(_abc_44694_new_n3518__bF_buf0), .Y(_abc_44694_new_n3934_));
OR2X2 OR2X2_1229 ( .A(_abc_44694_new_n3806_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n3935_));
OR2X2 OR2X2_123 ( .A(_abc_44694_new_n934_), .B(_abc_44694_new_n817__bF_buf1), .Y(_abc_44694_new_n935_));
OR2X2 OR2X2_1230 ( .A(_abc_44694_new_n3937_), .B(_abc_44694_new_n3924_), .Y(_0mem_dat_o_31_0__24_));
OR2X2 OR2X2_1231 ( .A(_abc_44694_new_n3940_), .B(_abc_44694_new_n3941_), .Y(_abc_44694_new_n3942_));
OR2X2 OR2X2_1232 ( .A(_abc_44694_new_n3942_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n3943_));
OR2X2 OR2X2_1233 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n3945_), .Y(_abc_44694_new_n3946_));
OR2X2 OR2X2_1234 ( .A(_abc_44694_new_n3944_), .B(_abc_44694_new_n3946_), .Y(_abc_44694_new_n3947_));
OR2X2 OR2X2_1235 ( .A(_abc_44694_new_n3948_), .B(_abc_44694_new_n3518__bF_buf3), .Y(_abc_44694_new_n3949_));
OR2X2 OR2X2_1236 ( .A(_abc_44694_new_n3821_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n3950_));
OR2X2 OR2X2_1237 ( .A(_abc_44694_new_n3952_), .B(_abc_44694_new_n3939_), .Y(_0mem_dat_o_31_0__25_));
OR2X2 OR2X2_1238 ( .A(_abc_44694_new_n3955_), .B(_abc_44694_new_n3956_), .Y(_abc_44694_new_n3957_));
OR2X2 OR2X2_1239 ( .A(_abc_44694_new_n3957_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n3958_));
OR2X2 OR2X2_124 ( .A(state_q_1_bF_buf0_), .B(alu_p_o_26_), .Y(_abc_44694_new_n936_));
OR2X2 OR2X2_1240 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n3960_), .Y(_abc_44694_new_n3961_));
OR2X2 OR2X2_1241 ( .A(_abc_44694_new_n3959_), .B(_abc_44694_new_n3961_), .Y(_abc_44694_new_n3962_));
OR2X2 OR2X2_1242 ( .A(_abc_44694_new_n3963_), .B(_abc_44694_new_n3518__bF_buf2), .Y(_abc_44694_new_n3964_));
OR2X2 OR2X2_1243 ( .A(_abc_44694_new_n3836_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n3965_));
OR2X2 OR2X2_1244 ( .A(_abc_44694_new_n3967_), .B(_abc_44694_new_n3954_), .Y(_0mem_dat_o_31_0__26_));
OR2X2 OR2X2_1245 ( .A(_abc_44694_new_n3970_), .B(_abc_44694_new_n3971_), .Y(_abc_44694_new_n3972_));
OR2X2 OR2X2_1246 ( .A(_abc_44694_new_n3972_), .B(_abc_44694_new_n3512__bF_buf0), .Y(_abc_44694_new_n3973_));
OR2X2 OR2X2_1247 ( .A(_abc_44694_new_n3513__bF_buf4), .B(_abc_44694_new_n3975_), .Y(_abc_44694_new_n3976_));
OR2X2 OR2X2_1248 ( .A(_abc_44694_new_n3974_), .B(_abc_44694_new_n3976_), .Y(_abc_44694_new_n3977_));
OR2X2 OR2X2_1249 ( .A(_abc_44694_new_n3978_), .B(_abc_44694_new_n3518__bF_buf1), .Y(_abc_44694_new_n3979_));
OR2X2 OR2X2_125 ( .A(_abc_44694_new_n938_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n939_));
OR2X2 OR2X2_1250 ( .A(_abc_44694_new_n3851_), .B(_abc_44694_new_n3519__bF_buf0), .Y(_abc_44694_new_n3980_));
OR2X2 OR2X2_1251 ( .A(_abc_44694_new_n3982_), .B(_abc_44694_new_n3969_), .Y(_0mem_dat_o_31_0__27_));
OR2X2 OR2X2_1252 ( .A(_abc_44694_new_n3985_), .B(_abc_44694_new_n3986_), .Y(_abc_44694_new_n3987_));
OR2X2 OR2X2_1253 ( .A(_abc_44694_new_n3987_), .B(_abc_44694_new_n3512__bF_buf4), .Y(_abc_44694_new_n3988_));
OR2X2 OR2X2_1254 ( .A(_abc_44694_new_n3513__bF_buf3), .B(_abc_44694_new_n3990_), .Y(_abc_44694_new_n3991_));
OR2X2 OR2X2_1255 ( .A(_abc_44694_new_n3989_), .B(_abc_44694_new_n3991_), .Y(_abc_44694_new_n3992_));
OR2X2 OR2X2_1256 ( .A(_abc_44694_new_n3993_), .B(_abc_44694_new_n3518__bF_buf0), .Y(_abc_44694_new_n3994_));
OR2X2 OR2X2_1257 ( .A(_abc_44694_new_n3866_), .B(_abc_44694_new_n3519__bF_buf4), .Y(_abc_44694_new_n3995_));
OR2X2 OR2X2_1258 ( .A(_abc_44694_new_n3997_), .B(_abc_44694_new_n3984_), .Y(_0mem_dat_o_31_0__28_));
OR2X2 OR2X2_1259 ( .A(_abc_44694_new_n4000_), .B(_abc_44694_new_n4001_), .Y(_abc_44694_new_n4002_));
OR2X2 OR2X2_126 ( .A(_abc_44694_new_n940_), .B(_abc_44694_new_n817__bF_buf0), .Y(_abc_44694_new_n941_));
OR2X2 OR2X2_1260 ( .A(_abc_44694_new_n4002_), .B(_abc_44694_new_n3512__bF_buf3), .Y(_abc_44694_new_n4003_));
OR2X2 OR2X2_1261 ( .A(_abc_44694_new_n3513__bF_buf2), .B(_abc_44694_new_n4005_), .Y(_abc_44694_new_n4006_));
OR2X2 OR2X2_1262 ( .A(_abc_44694_new_n4004_), .B(_abc_44694_new_n4006_), .Y(_abc_44694_new_n4007_));
OR2X2 OR2X2_1263 ( .A(_abc_44694_new_n4008_), .B(_abc_44694_new_n3518__bF_buf3), .Y(_abc_44694_new_n4009_));
OR2X2 OR2X2_1264 ( .A(_abc_44694_new_n3881_), .B(_abc_44694_new_n3519__bF_buf3), .Y(_abc_44694_new_n4010_));
OR2X2 OR2X2_1265 ( .A(_abc_44694_new_n4012_), .B(_abc_44694_new_n3999_), .Y(_0mem_dat_o_31_0__29_));
OR2X2 OR2X2_1266 ( .A(_abc_44694_new_n4015_), .B(_abc_44694_new_n4016_), .Y(_abc_44694_new_n4017_));
OR2X2 OR2X2_1267 ( .A(_abc_44694_new_n4017_), .B(_abc_44694_new_n3512__bF_buf2), .Y(_abc_44694_new_n4018_));
OR2X2 OR2X2_1268 ( .A(_abc_44694_new_n3513__bF_buf1), .B(_abc_44694_new_n4020_), .Y(_abc_44694_new_n4021_));
OR2X2 OR2X2_1269 ( .A(_abc_44694_new_n4019_), .B(_abc_44694_new_n4021_), .Y(_abc_44694_new_n4022_));
OR2X2 OR2X2_127 ( .A(state_q_1_bF_buf4_), .B(alu_p_o_27_), .Y(_abc_44694_new_n942_));
OR2X2 OR2X2_1270 ( .A(_abc_44694_new_n4023_), .B(_abc_44694_new_n3518__bF_buf2), .Y(_abc_44694_new_n4024_));
OR2X2 OR2X2_1271 ( .A(_abc_44694_new_n3896_), .B(_abc_44694_new_n3519__bF_buf2), .Y(_abc_44694_new_n4025_));
OR2X2 OR2X2_1272 ( .A(_abc_44694_new_n4027_), .B(_abc_44694_new_n4014_), .Y(_0mem_dat_o_31_0__30_));
OR2X2 OR2X2_1273 ( .A(_abc_44694_new_n4030_), .B(_abc_44694_new_n4031_), .Y(_abc_44694_new_n4032_));
OR2X2 OR2X2_1274 ( .A(_abc_44694_new_n4032_), .B(_abc_44694_new_n3512__bF_buf1), .Y(_abc_44694_new_n4033_));
OR2X2 OR2X2_1275 ( .A(_abc_44694_new_n3513__bF_buf0), .B(_abc_44694_new_n4035_), .Y(_abc_44694_new_n4036_));
OR2X2 OR2X2_1276 ( .A(_abc_44694_new_n4034_), .B(_abc_44694_new_n4036_), .Y(_abc_44694_new_n4037_));
OR2X2 OR2X2_1277 ( .A(_abc_44694_new_n4038_), .B(_abc_44694_new_n3518__bF_buf1), .Y(_abc_44694_new_n4039_));
OR2X2 OR2X2_1278 ( .A(_abc_44694_new_n3911_), .B(_abc_44694_new_n3519__bF_buf1), .Y(_abc_44694_new_n4040_));
OR2X2 OR2X2_1279 ( .A(_abc_44694_new_n4042_), .B(_abc_44694_new_n4029_), .Y(_0mem_dat_o_31_0__31_));
OR2X2 OR2X2_128 ( .A(_abc_44694_new_n944_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n945_));
OR2X2 OR2X2_1280 ( .A(_abc_44694_new_n3537_), .B(_abc_44694_new_n3520__bF_buf1), .Y(_abc_44694_new_n4044_));
OR2X2 OR2X2_1281 ( .A(_abc_44694_new_n4044_), .B(_auto_iopadmap_cc_368_execute_48790), .Y(_abc_44694_new_n4045_));
OR2X2 OR2X2_1282 ( .A(_abc_44694_new_n3527__bF_buf1), .B(_abc_44694_new_n4048_), .Y(_abc_44694_new_n4049_));
OR2X2 OR2X2_1283 ( .A(_abc_44694_new_n4044_), .B(_abc_44694_new_n653_), .Y(_abc_44694_new_n4051_));
OR2X2 OR2X2_1284 ( .A(_abc_44694_new_n4053_), .B(state_q_3_bF_buf3_), .Y(_abc_44694_new_n4054_));
OR2X2 OR2X2_1285 ( .A(_abc_44694_new_n4052_), .B(_abc_44694_new_n4054_), .Y(_0mem_stb_o_0_0_));
OR2X2 OR2X2_1286 ( .A(_abc_44694_new_n664_), .B(state_q_5_bF_buf2_), .Y(_abc_44694_new_n4058_));
OR2X2 OR2X2_1287 ( .A(_abc_44694_new_n4058_), .B(_abc_44694_new_n4057_), .Y(_abc_44694_new_n4059_));
OR2X2 OR2X2_1288 ( .A(_abc_44694_new_n4060_), .B(state_q_3_bF_buf2_), .Y(_abc_44694_new_n4061_));
OR2X2 OR2X2_1289 ( .A(_abc_44694_new_n4052_), .B(_abc_44694_new_n4061_), .Y(_0mem_cyc_o_0_0_));
OR2X2 OR2X2_129 ( .A(_abc_44694_new_n946_), .B(_abc_44694_new_n817__bF_buf3), .Y(_abc_44694_new_n947_));
OR2X2 OR2X2_1290 ( .A(_abc_44694_new_n656_), .B(_abc_44694_new_n4047_), .Y(_abc_44694_new_n4064_));
OR2X2 OR2X2_1291 ( .A(_abc_44694_new_n4065_), .B(_abc_44694_new_n4063_), .Y(_0mem_addr_o_31_0__0_));
OR2X2 OR2X2_1292 ( .A(_abc_44694_new_n4068_), .B(_abc_44694_new_n4067_), .Y(_0mem_addr_o_31_0__1_));
OR2X2 OR2X2_1293 ( .A(_abc_44694_new_n3342_), .B(_abc_44694_new_n3339_), .Y(_abc_44694_new_n4072_));
OR2X2 OR2X2_1294 ( .A(_abc_44694_new_n4072_), .B(_abc_44694_new_n4075_), .Y(_abc_44694_new_n4078_));
OR2X2 OR2X2_1295 ( .A(_abc_44694_new_n4080_), .B(_abc_44694_new_n4071_), .Y(_abc_44694_new_n4081_));
OR2X2 OR2X2_1296 ( .A(_abc_44694_new_n4081_), .B(_abc_44694_new_n4070_), .Y(_0mem_addr_o_31_0__2_));
OR2X2 OR2X2_1297 ( .A(_abc_44694_new_n4086_), .B(_abc_44694_new_n4089_), .Y(_abc_44694_new_n4090_));
OR2X2 OR2X2_1298 ( .A(_abc_44694_new_n4085_), .B(_abc_44694_new_n4091_), .Y(_abc_44694_new_n4092_));
OR2X2 OR2X2_1299 ( .A(_abc_44694_new_n4094_), .B(_abc_44694_new_n4084_), .Y(_abc_44694_new_n4095_));
OR2X2 OR2X2_13 ( .A(_abc_44694_new_n685_), .B(_abc_44694_new_n695_), .Y(_abc_44694_new_n696_));
OR2X2 OR2X2_130 ( .A(state_q_1_bF_buf3_), .B(alu_p_o_28_), .Y(_abc_44694_new_n948_));
OR2X2 OR2X2_1300 ( .A(_abc_44694_new_n4095_), .B(_abc_44694_new_n4083_), .Y(_0mem_addr_o_31_0__3_));
OR2X2 OR2X2_1301 ( .A(_abc_44694_new_n4085_), .B(_abc_44694_new_n1005_), .Y(_abc_44694_new_n4100_));
OR2X2 OR2X2_1302 ( .A(_abc_44694_new_n4102_), .B(_abc_44694_new_n4099_), .Y(_abc_44694_new_n4103_));
OR2X2 OR2X2_1303 ( .A(_abc_44694_new_n4101_), .B(_abc_44694_new_n4104_), .Y(_abc_44694_new_n4105_));
OR2X2 OR2X2_1304 ( .A(_abc_44694_new_n4109_), .B(_abc_44694_new_n4108_), .Y(_abc_44694_new_n4110_));
OR2X2 OR2X2_1305 ( .A(_abc_44694_new_n4107_), .B(_abc_44694_new_n4110_), .Y(_0mem_addr_o_31_0__4_));
OR2X2 OR2X2_1306 ( .A(_abc_44694_new_n4112_), .B(_abc_44694_new_n4116_), .Y(_abc_44694_new_n4117_));
OR2X2 OR2X2_1307 ( .A(_abc_44694_new_n4118_), .B(_abc_44694_new_n4115_), .Y(_abc_44694_new_n4119_));
OR2X2 OR2X2_1308 ( .A(_abc_44694_new_n4123_), .B(_abc_44694_new_n4122_), .Y(_abc_44694_new_n4124_));
OR2X2 OR2X2_1309 ( .A(_abc_44694_new_n4121_), .B(_abc_44694_new_n4124_), .Y(_0mem_addr_o_31_0__5_));
OR2X2 OR2X2_131 ( .A(_abc_44694_new_n950_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n951_));
OR2X2 OR2X2_1310 ( .A(_abc_44694_new_n4127_), .B(_abc_44694_new_n4130_), .Y(_abc_44694_new_n4131_));
OR2X2 OR2X2_1311 ( .A(_abc_44694_new_n4137_), .B(_abc_44694_new_n4136_), .Y(_abc_44694_new_n4138_));
OR2X2 OR2X2_1312 ( .A(_abc_44694_new_n4135_), .B(_abc_44694_new_n4138_), .Y(_0mem_addr_o_31_0__6_));
OR2X2 OR2X2_1313 ( .A(_abc_44694_new_n668__bF_buf0), .B(_abc_44694_new_n4140_), .Y(_abc_44694_new_n4141_));
OR2X2 OR2X2_1314 ( .A(_abc_44694_new_n4149_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4150_));
OR2X2 OR2X2_1315 ( .A(_abc_44694_new_n4150_), .B(_abc_44694_new_n4148_), .Y(_abc_44694_new_n4151_));
OR2X2 OR2X2_1316 ( .A(_abc_44694_new_n4153_), .B(_abc_44694_new_n4154_), .Y(_abc_44694_new_n4155_));
OR2X2 OR2X2_1317 ( .A(_abc_44694_new_n4152_), .B(_abc_44694_new_n4155_), .Y(_0mem_addr_o_31_0__7_));
OR2X2 OR2X2_1318 ( .A(_abc_44694_new_n4157_), .B(_abc_44694_new_n4144_), .Y(_abc_44694_new_n4158_));
OR2X2 OR2X2_1319 ( .A(_abc_44694_new_n4126_), .B(_abc_44694_new_n4161_), .Y(_abc_44694_new_n4162_));
OR2X2 OR2X2_132 ( .A(_abc_44694_new_n952_), .B(_abc_44694_new_n817__bF_buf2), .Y(_abc_44694_new_n953_));
OR2X2 OR2X2_1320 ( .A(_abc_44694_new_n4164_), .B(_abc_44694_new_n4167_), .Y(_abc_44694_new_n4168_));
OR2X2 OR2X2_1321 ( .A(_abc_44694_new_n4174_), .B(_abc_44694_new_n4173_), .Y(_abc_44694_new_n4175_));
OR2X2 OR2X2_1322 ( .A(_abc_44694_new_n4172_), .B(_abc_44694_new_n4175_), .Y(_0mem_addr_o_31_0__8_));
OR2X2 OR2X2_1323 ( .A(_abc_44694_new_n4181_), .B(_abc_44694_new_n4179_), .Y(_abc_44694_new_n4184_));
OR2X2 OR2X2_1324 ( .A(_abc_44694_new_n4188_), .B(_abc_44694_new_n4187_), .Y(_abc_44694_new_n4189_));
OR2X2 OR2X2_1325 ( .A(_abc_44694_new_n4186_), .B(_abc_44694_new_n4189_), .Y(_0mem_addr_o_31_0__9_));
OR2X2 OR2X2_1326 ( .A(_abc_44694_new_n4163_), .B(_abc_44694_new_n4192_), .Y(_abc_44694_new_n4193_));
OR2X2 OR2X2_1327 ( .A(_abc_44694_new_n4194_), .B(_abc_44694_new_n4177_), .Y(_abc_44694_new_n4195_));
OR2X2 OR2X2_1328 ( .A(_abc_44694_new_n4198_), .B(_abc_44694_new_n4201_), .Y(_abc_44694_new_n4204_));
OR2X2 OR2X2_1329 ( .A(_abc_44694_new_n4208_), .B(_abc_44694_new_n4207_), .Y(_abc_44694_new_n4209_));
OR2X2 OR2X2_133 ( .A(state_q_1_bF_buf2_), .B(alu_p_o_29_), .Y(_abc_44694_new_n954_));
OR2X2 OR2X2_1330 ( .A(_abc_44694_new_n4206_), .B(_abc_44694_new_n4209_), .Y(_0mem_addr_o_31_0__10_));
OR2X2 OR2X2_1331 ( .A(_abc_44694_new_n4213_), .B(_abc_44694_new_n4212_), .Y(_abc_44694_new_n4214_));
OR2X2 OR2X2_1332 ( .A(_abc_44694_new_n4214_), .B(REGFILE_SIM_reg_bank_reg_ra_o_11_), .Y(_abc_44694_new_n4217_));
OR2X2 OR2X2_1333 ( .A(_abc_44694_new_n4222_), .B(_abc_44694_new_n4219_), .Y(_abc_44694_new_n4223_));
OR2X2 OR2X2_1334 ( .A(_abc_44694_new_n4226_), .B(_abc_44694_new_n4225_), .Y(_abc_44694_new_n4227_));
OR2X2 OR2X2_1335 ( .A(_abc_44694_new_n4224_), .B(_abc_44694_new_n4227_), .Y(_0mem_addr_o_31_0__11_));
OR2X2 OR2X2_1336 ( .A(_abc_44694_new_n4230_), .B(_abc_44694_new_n4229_), .Y(_abc_44694_new_n4231_));
OR2X2 OR2X2_1337 ( .A(_abc_44694_new_n4231_), .B(REGFILE_SIM_reg_bank_reg_ra_o_12_), .Y(_abc_44694_new_n4234_));
OR2X2 OR2X2_1338 ( .A(_abc_44694_new_n4215_), .B(_abc_44694_new_n4199_), .Y(_abc_44694_new_n4236_));
OR2X2 OR2X2_1339 ( .A(_abc_44694_new_n4239_), .B(_abc_44694_new_n4237_), .Y(_abc_44694_new_n4240_));
OR2X2 OR2X2_134 ( .A(_abc_44694_new_n956_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n957_));
OR2X2 OR2X2_1340 ( .A(_abc_44694_new_n4242_), .B(_abc_44694_new_n4240_), .Y(_abc_44694_new_n4243_));
OR2X2 OR2X2_1341 ( .A(_abc_44694_new_n4243_), .B(_abc_44694_new_n4235_), .Y(_abc_44694_new_n4244_));
OR2X2 OR2X2_1342 ( .A(_abc_44694_new_n4250_), .B(_abc_44694_new_n4249_), .Y(_abc_44694_new_n4251_));
OR2X2 OR2X2_1343 ( .A(_abc_44694_new_n4248_), .B(_abc_44694_new_n4251_), .Y(_0mem_addr_o_31_0__12_));
OR2X2 OR2X2_1344 ( .A(_abc_44694_new_n4254_), .B(_abc_44694_new_n4253_), .Y(_abc_44694_new_n4255_));
OR2X2 OR2X2_1345 ( .A(_abc_44694_new_n4255_), .B(REGFILE_SIM_reg_bank_reg_ra_o_13_), .Y(_abc_44694_new_n4258_));
OR2X2 OR2X2_1346 ( .A(_abc_44694_new_n4259_), .B(_abc_44694_new_n4232_), .Y(_abc_44694_new_n4260_));
OR2X2 OR2X2_1347 ( .A(_abc_44694_new_n4245_), .B(_abc_44694_new_n4260_), .Y(_abc_44694_new_n4261_));
OR2X2 OR2X2_1348 ( .A(_abc_44694_new_n4271_), .B(_abc_44694_new_n4270_), .Y(_abc_44694_new_n4272_));
OR2X2 OR2X2_1349 ( .A(_abc_44694_new_n4269_), .B(_abc_44694_new_n4272_), .Y(_0mem_addr_o_31_0__13_));
OR2X2 OR2X2_135 ( .A(_abc_44694_new_n958_), .B(_abc_44694_new_n817__bF_buf1), .Y(_abc_44694_new_n959_));
OR2X2 OR2X2_1350 ( .A(_abc_44694_new_n4278_), .B(_abc_44694_new_n4277_), .Y(_abc_44694_new_n4279_));
OR2X2 OR2X2_1351 ( .A(_abc_44694_new_n4279_), .B(REGFILE_SIM_reg_bank_reg_ra_o_14_), .Y(_abc_44694_new_n4282_));
OR2X2 OR2X2_1352 ( .A(_abc_44694_new_n4276_), .B(_abc_44694_new_n4283_), .Y(_abc_44694_new_n4284_));
OR2X2 OR2X2_1353 ( .A(_abc_44694_new_n4290_), .B(_abc_44694_new_n4289_), .Y(_abc_44694_new_n4291_));
OR2X2 OR2X2_1354 ( .A(_abc_44694_new_n4288_), .B(_abc_44694_new_n4291_), .Y(_0mem_addr_o_31_0__14_));
OR2X2 OR2X2_1355 ( .A(_abc_44694_new_n4296_), .B(_abc_44694_new_n4295_), .Y(_abc_44694_new_n4297_));
OR2X2 OR2X2_1356 ( .A(_abc_44694_new_n4306_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4307_));
OR2X2 OR2X2_1357 ( .A(_abc_44694_new_n4307_), .B(_abc_44694_new_n4305_), .Y(_abc_44694_new_n4308_));
OR2X2 OR2X2_1358 ( .A(_abc_44694_new_n667_), .B(_auto_iopadmap_cc_368_execute_48711_15_), .Y(_abc_44694_new_n4309_));
OR2X2 OR2X2_1359 ( .A(_abc_44694_new_n4312_), .B(_abc_44694_new_n4313_), .Y(_abc_44694_new_n4314_));
OR2X2 OR2X2_136 ( .A(state_q_1_bF_buf1_), .B(alu_p_o_30_), .Y(_abc_44694_new_n960_));
OR2X2 OR2X2_1360 ( .A(_abc_44694_new_n4311_), .B(_abc_44694_new_n4314_), .Y(_0mem_addr_o_31_0__15_));
OR2X2 OR2X2_1361 ( .A(_abc_44694_new_n4297__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_16_), .Y(_abc_44694_new_n4318_));
OR2X2 OR2X2_1362 ( .A(_abc_44694_new_n4320_), .B(_abc_44694_new_n4298_), .Y(_abc_44694_new_n4321_));
OR2X2 OR2X2_1363 ( .A(_abc_44694_new_n4263_), .B(_abc_44694_new_n4324_), .Y(_abc_44694_new_n4325_));
OR2X2 OR2X2_1364 ( .A(_abc_44694_new_n4321_), .B(_abc_44694_new_n4326_), .Y(_abc_44694_new_n4327_));
OR2X2 OR2X2_1365 ( .A(_abc_44694_new_n4328_), .B(_abc_44694_new_n4319_), .Y(_abc_44694_new_n4329_));
OR2X2 OR2X2_1366 ( .A(_abc_44694_new_n4335_), .B(_abc_44694_new_n4334_), .Y(_abc_44694_new_n4336_));
OR2X2 OR2X2_1367 ( .A(_abc_44694_new_n4333_), .B(_abc_44694_new_n4336_), .Y(_0mem_addr_o_31_0__16_));
OR2X2 OR2X2_1368 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_17_), .Y(_abc_44694_new_n4342_));
OR2X2 OR2X2_1369 ( .A(_abc_44694_new_n4346_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4347_));
OR2X2 OR2X2_137 ( .A(_abc_44694_new_n962_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n963_));
OR2X2 OR2X2_1370 ( .A(_abc_44694_new_n4347_), .B(_abc_44694_new_n4345_), .Y(_abc_44694_new_n4348_));
OR2X2 OR2X2_1371 ( .A(_abc_44694_new_n667_), .B(_auto_iopadmap_cc_368_execute_48711_17_), .Y(_abc_44694_new_n4349_));
OR2X2 OR2X2_1372 ( .A(_abc_44694_new_n4352_), .B(_abc_44694_new_n4353_), .Y(_abc_44694_new_n4354_));
OR2X2 OR2X2_1373 ( .A(_abc_44694_new_n4351_), .B(_abc_44694_new_n4354_), .Y(_0mem_addr_o_31_0__17_));
OR2X2 OR2X2_1374 ( .A(_abc_44694_new_n4297__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_18_), .Y(_abc_44694_new_n4358_));
OR2X2 OR2X2_1375 ( .A(_abc_44694_new_n4363_), .B(_abc_44694_new_n4361_), .Y(_abc_44694_new_n4364_));
OR2X2 OR2X2_1376 ( .A(_abc_44694_new_n4364_), .B(_abc_44694_new_n4359_), .Y(_abc_44694_new_n4365_));
OR2X2 OR2X2_1377 ( .A(_abc_44694_new_n4371_), .B(_abc_44694_new_n4370_), .Y(_abc_44694_new_n4372_));
OR2X2 OR2X2_1378 ( .A(_abc_44694_new_n4369_), .B(_abc_44694_new_n4372_), .Y(_0mem_addr_o_31_0__18_));
OR2X2 OR2X2_1379 ( .A(_abc_44694_new_n4297__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_19_), .Y(_abc_44694_new_n4378_));
OR2X2 OR2X2_138 ( .A(_abc_44694_new_n964_), .B(_abc_44694_new_n817__bF_buf0), .Y(_abc_44694_new_n965_));
OR2X2 OR2X2_1380 ( .A(_abc_44694_new_n4382_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4383_));
OR2X2 OR2X2_1381 ( .A(_abc_44694_new_n4383_), .B(_abc_44694_new_n4381_), .Y(_abc_44694_new_n4384_));
OR2X2 OR2X2_1382 ( .A(_abc_44694_new_n667_), .B(_auto_iopadmap_cc_368_execute_48711_19_), .Y(_abc_44694_new_n4385_));
OR2X2 OR2X2_1383 ( .A(_abc_44694_new_n4388_), .B(_abc_44694_new_n4389_), .Y(_abc_44694_new_n4390_));
OR2X2 OR2X2_1384 ( .A(_abc_44694_new_n4387_), .B(_abc_44694_new_n4390_), .Y(_0mem_addr_o_31_0__19_));
OR2X2 OR2X2_1385 ( .A(_abc_44694_new_n4394_), .B(_abc_44694_new_n4399_), .Y(_abc_44694_new_n4400_));
OR2X2 OR2X2_1386 ( .A(_abc_44694_new_n4297__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_20_), .Y(_abc_44694_new_n4403_));
OR2X2 OR2X2_1387 ( .A(_abc_44694_new_n4400_), .B(_abc_44694_new_n4404_), .Y(_abc_44694_new_n4405_));
OR2X2 OR2X2_1388 ( .A(_abc_44694_new_n4411_), .B(_abc_44694_new_n4410_), .Y(_abc_44694_new_n4412_));
OR2X2 OR2X2_1389 ( .A(_abc_44694_new_n4409_), .B(_abc_44694_new_n4412_), .Y(_0mem_addr_o_31_0__20_));
OR2X2 OR2X2_139 ( .A(state_q_1_bF_buf0_), .B(alu_p_o_31_), .Y(_abc_44694_new_n966_));
OR2X2 OR2X2_1390 ( .A(_abc_44694_new_n4297__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_21_), .Y(_abc_44694_new_n4417_));
OR2X2 OR2X2_1391 ( .A(_abc_44694_new_n4414_), .B(_abc_44694_new_n4419_), .Y(_abc_44694_new_n4420_));
OR2X2 OR2X2_1392 ( .A(_abc_44694_new_n4421_), .B(_abc_44694_new_n4418_), .Y(_abc_44694_new_n4422_));
OR2X2 OR2X2_1393 ( .A(_abc_44694_new_n4426_), .B(_abc_44694_new_n4425_), .Y(_abc_44694_new_n4427_));
OR2X2 OR2X2_1394 ( .A(_abc_44694_new_n4424_), .B(_abc_44694_new_n4427_), .Y(_0mem_addr_o_31_0__21_));
OR2X2 OR2X2_1395 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_22_), .Y(_abc_44694_new_n4431_));
OR2X2 OR2X2_1396 ( .A(_abc_44694_new_n4436_), .B(_abc_44694_new_n4434_), .Y(_abc_44694_new_n4437_));
OR2X2 OR2X2_1397 ( .A(_abc_44694_new_n4437_), .B(_abc_44694_new_n4432_), .Y(_abc_44694_new_n4438_));
OR2X2 OR2X2_1398 ( .A(_abc_44694_new_n4444_), .B(_abc_44694_new_n4443_), .Y(_abc_44694_new_n4445_));
OR2X2 OR2X2_1399 ( .A(_abc_44694_new_n4442_), .B(_abc_44694_new_n4445_), .Y(_0mem_addr_o_31_0__22_));
OR2X2 OR2X2_14 ( .A(_abc_44694_new_n697_), .B(_abc_44694_new_n672_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_0_));
OR2X2 OR2X2_140 ( .A(_abc_44694_new_n660_), .B(state_q_4_), .Y(REGFILE_SIM_reg_bank_wr_i));
OR2X2 OR2X2_1400 ( .A(_abc_44694_new_n4297__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_ra_o_23_), .Y(_abc_44694_new_n4451_));
OR2X2 OR2X2_1401 ( .A(_abc_44694_new_n4455_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4456_));
OR2X2 OR2X2_1402 ( .A(_abc_44694_new_n4456_), .B(_abc_44694_new_n4454_), .Y(_abc_44694_new_n4457_));
OR2X2 OR2X2_1403 ( .A(_abc_44694_new_n667_), .B(_auto_iopadmap_cc_368_execute_48711_23_), .Y(_abc_44694_new_n4458_));
OR2X2 OR2X2_1404 ( .A(_abc_44694_new_n4461_), .B(_abc_44694_new_n4462_), .Y(_abc_44694_new_n4463_));
OR2X2 OR2X2_1405 ( .A(_abc_44694_new_n4460_), .B(_abc_44694_new_n4463_), .Y(_0mem_addr_o_31_0__23_));
OR2X2 OR2X2_1406 ( .A(_abc_44694_new_n4398_), .B(_abc_44694_new_n4471_), .Y(_abc_44694_new_n4472_));
OR2X2 OR2X2_1407 ( .A(_abc_44694_new_n4474_), .B(_abc_44694_new_n4476_), .Y(_abc_44694_new_n4477_));
OR2X2 OR2X2_1408 ( .A(_abc_44694_new_n4297__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_24_), .Y(_abc_44694_new_n4482_));
OR2X2 OR2X2_1409 ( .A(_abc_44694_new_n4479_), .B(_abc_44694_new_n4483_), .Y(_abc_44694_new_n4484_));
OR2X2 OR2X2_141 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_8_), .B(alu_op_r_6_), .Y(_abc_44694_new_n972_));
OR2X2 OR2X2_1410 ( .A(_abc_44694_new_n4490_), .B(_abc_44694_new_n4489_), .Y(_abc_44694_new_n4491_));
OR2X2 OR2X2_1411 ( .A(_abc_44694_new_n4488_), .B(_abc_44694_new_n4491_), .Y(_0mem_addr_o_31_0__24_));
OR2X2 OR2X2_1412 ( .A(_abc_44694_new_n4297__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_ra_o_25_), .Y(_abc_44694_new_n4497_));
OR2X2 OR2X2_1413 ( .A(_abc_44694_new_n4501_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4502_));
OR2X2 OR2X2_1414 ( .A(_abc_44694_new_n4502_), .B(_abc_44694_new_n4500_), .Y(_abc_44694_new_n4503_));
OR2X2 OR2X2_1415 ( .A(_abc_44694_new_n667_), .B(_auto_iopadmap_cc_368_execute_48711_25_), .Y(_abc_44694_new_n4504_));
OR2X2 OR2X2_1416 ( .A(_abc_44694_new_n4507_), .B(_abc_44694_new_n4508_), .Y(_abc_44694_new_n4509_));
OR2X2 OR2X2_1417 ( .A(_abc_44694_new_n4506_), .B(_abc_44694_new_n4509_), .Y(_0mem_addr_o_31_0__25_));
OR2X2 OR2X2_1418 ( .A(_abc_44694_new_n4478_), .B(_abc_44694_new_n4512_), .Y(_abc_44694_new_n4513_));
OR2X2 OR2X2_1419 ( .A(_abc_44694_new_n4297__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_ra_o_26_), .Y(_abc_44694_new_n4519_));
OR2X2 OR2X2_142 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_9_), .B(alu_op_r_7_), .Y(_abc_44694_new_n974_));
OR2X2 OR2X2_1420 ( .A(_abc_44694_new_n4516_), .B(_abc_44694_new_n4520_), .Y(_abc_44694_new_n4521_));
OR2X2 OR2X2_1421 ( .A(_abc_44694_new_n4527_), .B(_abc_44694_new_n4526_), .Y(_abc_44694_new_n4528_));
OR2X2 OR2X2_1422 ( .A(_abc_44694_new_n4525_), .B(_abc_44694_new_n4528_), .Y(_0mem_addr_o_31_0__26_));
OR2X2 OR2X2_1423 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_27_), .Y(_abc_44694_new_n4534_));
OR2X2 OR2X2_1424 ( .A(_abc_44694_new_n4531_), .B(_abc_44694_new_n4535_), .Y(_abc_44694_new_n4536_));
OR2X2 OR2X2_1425 ( .A(_abc_44694_new_n4530_), .B(_abc_44694_new_n4537_), .Y(_abc_44694_new_n4538_));
OR2X2 OR2X2_1426 ( .A(_abc_44694_new_n4542_), .B(_abc_44694_new_n4541_), .Y(_abc_44694_new_n4543_));
OR2X2 OR2X2_1427 ( .A(_abc_44694_new_n4540_), .B(_abc_44694_new_n4543_), .Y(_0mem_addr_o_31_0__27_));
OR2X2 OR2X2_1428 ( .A(_abc_44694_new_n4549_), .B(_abc_44694_new_n4514_), .Y(_abc_44694_new_n4550_));
OR2X2 OR2X2_1429 ( .A(_abc_44694_new_n4557_), .B(_abc_44694_new_n4555_), .Y(_abc_44694_new_n4558_));
OR2X2 OR2X2_143 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_10_), .B(int32_r_10_), .Y(_abc_44694_new_n985_));
OR2X2 OR2X2_1430 ( .A(_abc_44694_new_n4554_), .B(_abc_44694_new_n4559_), .Y(_abc_44694_new_n4560_));
OR2X2 OR2X2_1431 ( .A(_abc_44694_new_n4566_), .B(_abc_44694_new_n4565_), .Y(_abc_44694_new_n4567_));
OR2X2 OR2X2_1432 ( .A(_abc_44694_new_n4564_), .B(_abc_44694_new_n4567_), .Y(_0mem_addr_o_31_0__28_));
OR2X2 OR2X2_1433 ( .A(_abc_44694_new_n4561_), .B(_abc_44694_new_n4555_), .Y(_abc_44694_new_n4569_));
OR2X2 OR2X2_1434 ( .A(_abc_44694_new_n4573_), .B(_abc_44694_new_n4571_), .Y(_abc_44694_new_n4574_));
OR2X2 OR2X2_1435 ( .A(_abc_44694_new_n4577_), .B(_abc_44694_new_n655_), .Y(_abc_44694_new_n4578_));
OR2X2 OR2X2_1436 ( .A(_abc_44694_new_n4578_), .B(_abc_44694_new_n4576_), .Y(_abc_44694_new_n4579_));
OR2X2 OR2X2_1437 ( .A(_abc_44694_new_n667_), .B(_auto_iopadmap_cc_368_execute_48711_29_), .Y(_abc_44694_new_n4580_));
OR2X2 OR2X2_1438 ( .A(_abc_44694_new_n4583_), .B(_abc_44694_new_n4584_), .Y(_abc_44694_new_n4585_));
OR2X2 OR2X2_1439 ( .A(_abc_44694_new_n4582_), .B(_abc_44694_new_n4585_), .Y(_0mem_addr_o_31_0__29_));
OR2X2 OR2X2_144 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_5_), .B(int32_r_5_), .Y(_abc_44694_new_n990_));
OR2X2 OR2X2_1440 ( .A(_abc_44694_new_n4297__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_ra_o_30_), .Y(_abc_44694_new_n4589_));
OR2X2 OR2X2_1441 ( .A(_abc_44694_new_n4300_), .B(_abc_44694_new_n4591_), .Y(_abc_44694_new_n4592_));
OR2X2 OR2X2_1442 ( .A(_abc_44694_new_n4553_), .B(_abc_44694_new_n4594_), .Y(_abc_44694_new_n4595_));
OR2X2 OR2X2_1443 ( .A(_abc_44694_new_n4597_), .B(_abc_44694_new_n4590_), .Y(_abc_44694_new_n4598_));
OR2X2 OR2X2_1444 ( .A(_abc_44694_new_n4596_), .B(_abc_44694_new_n4599_), .Y(_abc_44694_new_n4600_));
OR2X2 OR2X2_1445 ( .A(_abc_44694_new_n4604_), .B(_abc_44694_new_n4603_), .Y(_abc_44694_new_n4605_));
OR2X2 OR2X2_1446 ( .A(_abc_44694_new_n4602_), .B(_abc_44694_new_n4605_), .Y(_0mem_addr_o_31_0__30_));
OR2X2 OR2X2_1447 ( .A(_abc_44694_new_n4300_), .B(_abc_44694_new_n4609_), .Y(_abc_44694_new_n4610_));
OR2X2 OR2X2_1448 ( .A(_abc_44694_new_n4297__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_ra_o_31_), .Y(_abc_44694_new_n4611_));
OR2X2 OR2X2_1449 ( .A(_abc_44694_new_n4614_), .B(_abc_44694_new_n4615_), .Y(_abc_44694_new_n4616_));
OR2X2 OR2X2_145 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_0_), .B(alu_op_r_0_), .Y(_abc_44694_new_n992_));
OR2X2 OR2X2_1450 ( .A(_abc_44694_new_n4619_), .B(_abc_44694_new_n4618_), .Y(_abc_44694_new_n4620_));
OR2X2 OR2X2_1451 ( .A(_abc_44694_new_n4617_), .B(_abc_44694_new_n4620_), .Y(_0mem_addr_o_31_0__31_));
OR2X2 OR2X2_1452 ( .A(_abc_44694_new_n4625_), .B(_auto_iopadmap_cc_368_execute_48709), .Y(_abc_44694_new_n4626_));
OR2X2 OR2X2_1453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2104_));
OR2X2 OR2X2_1454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2109_));
OR2X2 OR2X2_1455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2114_));
OR2X2 OR2X2_1456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2119_));
OR2X2 OR2X2_1457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2124_));
OR2X2 OR2X2_1458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2129_));
OR2X2 OR2X2_1459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2134_));
OR2X2 OR2X2_146 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_4_), .B(int32_r_4_), .Y(_abc_44694_new_n994_));
OR2X2 OR2X2_1460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2139_));
OR2X2 OR2X2_1461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2144_));
OR2X2 OR2X2_1462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2149_));
OR2X2 OR2X2_1463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2154_));
OR2X2 OR2X2_1464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2159_));
OR2X2 OR2X2_1465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2164_));
OR2X2 OR2X2_1466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2169_));
OR2X2 OR2X2_1467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2174_));
OR2X2 OR2X2_1468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2179_));
OR2X2 OR2X2_1469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2184_));
OR2X2 OR2X2_147 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_1_), .B(alu_op_r_1_), .Y(_abc_44694_new_n995_));
OR2X2 OR2X2_1470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2189_));
OR2X2 OR2X2_1471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2194_));
OR2X2 OR2X2_1472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2199_));
OR2X2 OR2X2_1473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2204_));
OR2X2 OR2X2_1474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2209_));
OR2X2 OR2X2_1475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2214_));
OR2X2 OR2X2_1476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2219_));
OR2X2 OR2X2_1477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2224_));
OR2X2 OR2X2_1478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2229_));
OR2X2 OR2X2_1479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2234_));
OR2X2 OR2X2_148 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_7_), .B(alu_op_r_5_), .Y(_abc_44694_new_n999_));
OR2X2 OR2X2_1480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2239_));
OR2X2 OR2X2_1481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r31_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2244_));
OR2X2 OR2X2_1482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r31_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2249_));
OR2X2 OR2X2_1483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r31_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2254_));
OR2X2 OR2X2_1484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2103__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r31_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2259_));
OR2X2 OR2X2_1485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2268_));
OR2X2 OR2X2_1486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2270_));
OR2X2 OR2X2_1487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2272_));
OR2X2 OR2X2_1488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2273_));
OR2X2 OR2X2_1489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2275_));
OR2X2 OR2X2_149 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_6_), .B(alu_op_r_4_), .Y(_abc_44694_new_n1001_));
OR2X2 OR2X2_1490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2276_));
OR2X2 OR2X2_1491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2278_));
OR2X2 OR2X2_1492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2279_));
OR2X2 OR2X2_1493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2281_));
OR2X2 OR2X2_1494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2282_));
OR2X2 OR2X2_1495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2284_));
OR2X2 OR2X2_1496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2285_));
OR2X2 OR2X2_1497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2287_));
OR2X2 OR2X2_1498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2288_));
OR2X2 OR2X2_1499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2290_));
OR2X2 OR2X2_15 ( .A(_abc_44694_new_n701_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n702_));
OR2X2 OR2X2_150 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_3_), .B(alu_op_r_3_), .Y(_abc_44694_new_n1004_));
OR2X2 OR2X2_1500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2291_));
OR2X2 OR2X2_1501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2293_));
OR2X2 OR2X2_1502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2294_));
OR2X2 OR2X2_1503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2296_));
OR2X2 OR2X2_1504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2297_));
OR2X2 OR2X2_1505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2299_));
OR2X2 OR2X2_1506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2300_));
OR2X2 OR2X2_1507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2302_));
OR2X2 OR2X2_1508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2303_));
OR2X2 OR2X2_1509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2305_));
OR2X2 OR2X2_151 ( .A(REGFILE_SIM_reg_bank_reg_ra_o_2_), .B(alu_op_r_2_), .Y(_abc_44694_new_n1006_));
OR2X2 OR2X2_1510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2306_));
OR2X2 OR2X2_1511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2308_));
OR2X2 OR2X2_1512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2309_));
OR2X2 OR2X2_1513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2311_));
OR2X2 OR2X2_1514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2312_));
OR2X2 OR2X2_1515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2314_));
OR2X2 OR2X2_1516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2315_));
OR2X2 OR2X2_1517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2317_));
OR2X2 OR2X2_1518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2318_));
OR2X2 OR2X2_1519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2320_));
OR2X2 OR2X2_152 ( .A(_abc_44694_new_n1011_), .B(_abc_44694_new_n971_), .Y(_abc_44694_new_n1012_));
OR2X2 OR2X2_1520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2321_));
OR2X2 OR2X2_1521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2323_));
OR2X2 OR2X2_1522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2324_));
OR2X2 OR2X2_1523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2326_));
OR2X2 OR2X2_1524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2327_));
OR2X2 OR2X2_1525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2329_));
OR2X2 OR2X2_1526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2330_));
OR2X2 OR2X2_1527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2332_));
OR2X2 OR2X2_1528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2333_));
OR2X2 OR2X2_1529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2335_));
OR2X2 OR2X2_153 ( .A(_abc_44694_new_n1022_), .B(_abc_44694_new_n1020_), .Y(_abc_44694_new_n1023_));
OR2X2 OR2X2_1530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2336_));
OR2X2 OR2X2_1531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2338_));
OR2X2 OR2X2_1532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2339_));
OR2X2 OR2X2_1533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2341_));
OR2X2 OR2X2_1534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2342_));
OR2X2 OR2X2_1535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2344_));
OR2X2 OR2X2_1536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2345_));
OR2X2 OR2X2_1537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2347_));
OR2X2 OR2X2_1538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2348_));
OR2X2 OR2X2_1539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r30_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2350_));
OR2X2 OR2X2_154 ( .A(_abc_44694_new_n1016_), .B(_abc_44694_new_n1025_), .Y(_abc_44694_new_n1026_));
OR2X2 OR2X2_1540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2351_));
OR2X2 OR2X2_1541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r30_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2353_));
OR2X2 OR2X2_1542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2354_));
OR2X2 OR2X2_1543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r30_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2356_));
OR2X2 OR2X2_1544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2357_));
OR2X2 OR2X2_1545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r30_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2359_));
OR2X2 OR2X2_1546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2360_));
OR2X2 OR2X2_1547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2267__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r30_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2362_));
OR2X2 OR2X2_1548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2269__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2363_));
OR2X2 OR2X2_1549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2369_));
OR2X2 OR2X2_155 ( .A(_abc_44694_new_n1040_), .B(_abc_44694_new_n1041_), .Y(_abc_44694_new_n1042_));
OR2X2 OR2X2_1550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2371_));
OR2X2 OR2X2_1551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2373_));
OR2X2 OR2X2_1552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2374_));
OR2X2 OR2X2_1553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2376_));
OR2X2 OR2X2_1554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2377_));
OR2X2 OR2X2_1555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2379_));
OR2X2 OR2X2_1556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2380_));
OR2X2 OR2X2_1557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2382_));
OR2X2 OR2X2_1558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2383_));
OR2X2 OR2X2_1559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2385_));
OR2X2 OR2X2_156 ( .A(_abc_44694_new_n1028_), .B(_abc_44694_new_n1042_), .Y(_abc_44694_new_n1043_));
OR2X2 OR2X2_1560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2386_));
OR2X2 OR2X2_1561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2388_));
OR2X2 OR2X2_1562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2389_));
OR2X2 OR2X2_1563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2391_));
OR2X2 OR2X2_1564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2392_));
OR2X2 OR2X2_1565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2394_));
OR2X2 OR2X2_1566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2395_));
OR2X2 OR2X2_1567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2397_));
OR2X2 OR2X2_1568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2398_));
OR2X2 OR2X2_1569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2400_));
OR2X2 OR2X2_157 ( .A(nmi_q), .B(nmi_i), .Y(_abc_44694_new_n1044_));
OR2X2 OR2X2_1570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2401_));
OR2X2 OR2X2_1571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2403_));
OR2X2 OR2X2_1572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2404_));
OR2X2 OR2X2_1573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2406_));
OR2X2 OR2X2_1574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2407_));
OR2X2 OR2X2_1575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2409_));
OR2X2 OR2X2_1576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2410_));
OR2X2 OR2X2_1577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2412_));
OR2X2 OR2X2_1578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2413_));
OR2X2 OR2X2_1579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2415_));
OR2X2 OR2X2_158 ( .A(inst_trap_w), .B(_abc_44694_new_n1048_), .Y(_abc_44694_new_n1049_));
OR2X2 OR2X2_1580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2416_));
OR2X2 OR2X2_1581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2418_));
OR2X2 OR2X2_1582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2419_));
OR2X2 OR2X2_1583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2421_));
OR2X2 OR2X2_1584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2422_));
OR2X2 OR2X2_1585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2424_));
OR2X2 OR2X2_1586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2425_));
OR2X2 OR2X2_1587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2427_));
OR2X2 OR2X2_1588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2428_));
OR2X2 OR2X2_1589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2430_));
OR2X2 OR2X2_159 ( .A(_abc_44694_new_n1067_), .B(_abc_44694_new_n1070_), .Y(_abc_44694_new_n1071_));
OR2X2 OR2X2_1590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2431_));
OR2X2 OR2X2_1591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2433_));
OR2X2 OR2X2_1592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2434_));
OR2X2 OR2X2_1593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2436_));
OR2X2 OR2X2_1594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2437_));
OR2X2 OR2X2_1595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2439_));
OR2X2 OR2X2_1596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2440_));
OR2X2 OR2X2_1597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2442_));
OR2X2 OR2X2_1598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2443_));
OR2X2 OR2X2_1599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2445_));
OR2X2 OR2X2_16 ( .A(_abc_44694_new_n702_), .B(_abc_44694_new_n700_), .Y(_abc_44694_new_n703_));
OR2X2 OR2X2_160 ( .A(_abc_44694_new_n1075_), .B(_abc_44694_new_n1078_), .Y(_abc_44694_new_n1079_));
OR2X2 OR2X2_1600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2446_));
OR2X2 OR2X2_1601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2448_));
OR2X2 OR2X2_1602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2449_));
OR2X2 OR2X2_1603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r29_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2451_));
OR2X2 OR2X2_1604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2452_));
OR2X2 OR2X2_1605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r29_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2454_));
OR2X2 OR2X2_1606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2455_));
OR2X2 OR2X2_1607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r29_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2457_));
OR2X2 OR2X2_1608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2458_));
OR2X2 OR2X2_1609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r29_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2460_));
OR2X2 OR2X2_161 ( .A(_abc_44694_new_n1072_), .B(_abc_44694_new_n1079_), .Y(_abc_44694_new_n1080_));
OR2X2 OR2X2_1610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2461_));
OR2X2 OR2X2_1611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2368__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r29_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2463_));
OR2X2 OR2X2_1612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2370__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2464_));
OR2X2 OR2X2_1613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2469_));
OR2X2 OR2X2_1614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2473_));
OR2X2 OR2X2_1615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2477_));
OR2X2 OR2X2_1616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2481_));
OR2X2 OR2X2_1617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2485_));
OR2X2 OR2X2_1618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2489_));
OR2X2 OR2X2_1619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2493_));
OR2X2 OR2X2_162 ( .A(_abc_44694_new_n1110_), .B(_abc_44694_new_n1104_), .Y(_abc_44694_new_n1111_));
OR2X2 OR2X2_1620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2497_));
OR2X2 OR2X2_1621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2501_));
OR2X2 OR2X2_1622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2505_));
OR2X2 OR2X2_1623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2509_));
OR2X2 OR2X2_1624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2513_));
OR2X2 OR2X2_1625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2517_));
OR2X2 OR2X2_1626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2521_));
OR2X2 OR2X2_1627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2525_));
OR2X2 OR2X2_1628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2529_));
OR2X2 OR2X2_1629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2533_));
OR2X2 OR2X2_163 ( .A(_abc_44694_new_n1111_), .B(_abc_44694_new_n1099_), .Y(_abc_44694_new_n1112_));
OR2X2 OR2X2_1630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2537_));
OR2X2 OR2X2_1631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2541_));
OR2X2 OR2X2_1632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2545_));
OR2X2 OR2X2_1633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2549_));
OR2X2 OR2X2_1634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2553_));
OR2X2 OR2X2_1635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2557_));
OR2X2 OR2X2_1636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2561_));
OR2X2 OR2X2_1637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2565_));
OR2X2 OR2X2_1638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2569_));
OR2X2 OR2X2_1639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2573_));
OR2X2 OR2X2_164 ( .A(_abc_44694_new_n1121_), .B(_abc_44694_new_n1123_), .Y(_abc_44694_new_n1124_));
OR2X2 OR2X2_1640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2577_));
OR2X2 OR2X2_1641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r28_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2581_));
OR2X2 OR2X2_1642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r28_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2585_));
OR2X2 OR2X2_1643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r28_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2589_));
OR2X2 OR2X2_1644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2468__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r28_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2593_));
OR2X2 OR2X2_1645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2601_));
OR2X2 OR2X2_1646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2603_));
OR2X2 OR2X2_1647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2605_));
OR2X2 OR2X2_1648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2606_));
OR2X2 OR2X2_1649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2608_));
OR2X2 OR2X2_165 ( .A(_abc_44694_new_n1124_), .B(_abc_44694_new_n1118_), .Y(_abc_44694_new_n1125_));
OR2X2 OR2X2_1650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2609_));
OR2X2 OR2X2_1651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2611_));
OR2X2 OR2X2_1652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2612_));
OR2X2 OR2X2_1653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2614_));
OR2X2 OR2X2_1654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2615_));
OR2X2 OR2X2_1655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2617_));
OR2X2 OR2X2_1656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2618_));
OR2X2 OR2X2_1657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2620_));
OR2X2 OR2X2_1658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2621_));
OR2X2 OR2X2_1659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2623_));
OR2X2 OR2X2_166 ( .A(_abc_44694_new_n1095_), .B(opcode_q_22_), .Y(_abc_44694_new_n1128_));
OR2X2 OR2X2_1660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2624_));
OR2X2 OR2X2_1661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2626_));
OR2X2 OR2X2_1662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2627_));
OR2X2 OR2X2_1663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2629_));
OR2X2 OR2X2_1664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2630_));
OR2X2 OR2X2_1665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2632_));
OR2X2 OR2X2_1666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2633_));
OR2X2 OR2X2_1667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2635_));
OR2X2 OR2X2_1668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2636_));
OR2X2 OR2X2_1669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2638_));
OR2X2 OR2X2_167 ( .A(_abc_44694_new_n1147_), .B(_abc_44694_new_n1146_), .Y(_abc_44694_new_n1148_));
OR2X2 OR2X2_1670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2639_));
OR2X2 OR2X2_1671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2641_));
OR2X2 OR2X2_1672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2642_));
OR2X2 OR2X2_1673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2644_));
OR2X2 OR2X2_1674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2645_));
OR2X2 OR2X2_1675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2647_));
OR2X2 OR2X2_1676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2648_));
OR2X2 OR2X2_1677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2650_));
OR2X2 OR2X2_1678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2651_));
OR2X2 OR2X2_1679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2653_));
OR2X2 OR2X2_168 ( .A(_abc_44694_new_n1148_), .B(_abc_44694_new_n1144_), .Y(_abc_44694_new_n1149_));
OR2X2 OR2X2_1680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2654_));
OR2X2 OR2X2_1681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2656_));
OR2X2 OR2X2_1682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2657_));
OR2X2 OR2X2_1683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2659_));
OR2X2 OR2X2_1684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2660_));
OR2X2 OR2X2_1685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2662_));
OR2X2 OR2X2_1686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2663_));
OR2X2 OR2X2_1687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2665_));
OR2X2 OR2X2_1688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2666_));
OR2X2 OR2X2_1689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2668_));
OR2X2 OR2X2_169 ( .A(_abc_44694_new_n1155_), .B(_abc_44694_new_n1159_), .Y(_abc_44694_new_n1160_));
OR2X2 OR2X2_1690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2669_));
OR2X2 OR2X2_1691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2671_));
OR2X2 OR2X2_1692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2672_));
OR2X2 OR2X2_1693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2674_));
OR2X2 OR2X2_1694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2675_));
OR2X2 OR2X2_1695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2677_));
OR2X2 OR2X2_1696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2678_));
OR2X2 OR2X2_1697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2680_));
OR2X2 OR2X2_1698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2681_));
OR2X2 OR2X2_1699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r27_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2683_));
OR2X2 OR2X2_17 ( .A(_abc_44694_new_n704_), .B(_abc_44694_new_n705_), .Y(_abc_44694_new_n706_));
OR2X2 OR2X2_170 ( .A(_abc_44694_new_n1160_), .B(_abc_44694_new_n1152_), .Y(_abc_44694_new_n1161_));
OR2X2 OR2X2_1700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2684_));
OR2X2 OR2X2_1701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r27_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2686_));
OR2X2 OR2X2_1702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2687_));
OR2X2 OR2X2_1703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r27_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2689_));
OR2X2 OR2X2_1704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2690_));
OR2X2 OR2X2_1705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r27_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2692_));
OR2X2 OR2X2_1706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2693_));
OR2X2 OR2X2_1707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2600__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r27_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2695_));
OR2X2 OR2X2_1708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2602__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2696_));
OR2X2 OR2X2_1709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2700_));
OR2X2 OR2X2_171 ( .A(_abc_44694_new_n1161_), .B(_abc_44694_new_n1149_), .Y(_abc_44694_new_n1162_));
OR2X2 OR2X2_1710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2704_));
OR2X2 OR2X2_1711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2708_));
OR2X2 OR2X2_1712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2712_));
OR2X2 OR2X2_1713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2716_));
OR2X2 OR2X2_1714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2720_));
OR2X2 OR2X2_1715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2724_));
OR2X2 OR2X2_1716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2728_));
OR2X2 OR2X2_1717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2732_));
OR2X2 OR2X2_1718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2736_));
OR2X2 OR2X2_1719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2740_));
OR2X2 OR2X2_172 ( .A(_abc_44694_new_n1166_), .B(_abc_44694_new_n1170_), .Y(_abc_44694_new_n1171_));
OR2X2 OR2X2_1720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2744_));
OR2X2 OR2X2_1721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2748_));
OR2X2 OR2X2_1722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2752_));
OR2X2 OR2X2_1723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2756_));
OR2X2 OR2X2_1724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2760_));
OR2X2 OR2X2_1725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2764_));
OR2X2 OR2X2_1726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2768_));
OR2X2 OR2X2_1727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2772_));
OR2X2 OR2X2_1728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2776_));
OR2X2 OR2X2_1729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2780_));
OR2X2 OR2X2_173 ( .A(_abc_44694_new_n1176_), .B(_abc_44694_new_n1177_), .Y(_abc_44694_new_n1178_));
OR2X2 OR2X2_1730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2784_));
OR2X2 OR2X2_1731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2788_));
OR2X2 OR2X2_1732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2792_));
OR2X2 OR2X2_1733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2796_));
OR2X2 OR2X2_1734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2800_));
OR2X2 OR2X2_1735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2804_));
OR2X2 OR2X2_1736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2808_));
OR2X2 OR2X2_1737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r26_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2812_));
OR2X2 OR2X2_1738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r26_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2816_));
OR2X2 OR2X2_1739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r26_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2820_));
OR2X2 OR2X2_174 ( .A(_abc_44694_new_n1182_), .B(_abc_44694_new_n1181__bF_buf3), .Y(_abc_44694_new_n1183_));
OR2X2 OR2X2_1740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2699__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r26_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2824_));
OR2X2 OR2X2_1741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2830_));
OR2X2 OR2X2_1742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2834_));
OR2X2 OR2X2_1743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2838_));
OR2X2 OR2X2_1744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2842_));
OR2X2 OR2X2_1745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2846_));
OR2X2 OR2X2_1746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2850_));
OR2X2 OR2X2_1747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2854_));
OR2X2 OR2X2_1748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2858_));
OR2X2 OR2X2_1749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2862_));
OR2X2 OR2X2_175 ( .A(_abc_44694_new_n1196_), .B(_abc_44694_new_n1197_), .Y(_abc_44694_new_n1198_));
OR2X2 OR2X2_1750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2866_));
OR2X2 OR2X2_1751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2870_));
OR2X2 OR2X2_1752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2874_));
OR2X2 OR2X2_1753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2878_));
OR2X2 OR2X2_1754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2882_));
OR2X2 OR2X2_1755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2886_));
OR2X2 OR2X2_1756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2890_));
OR2X2 OR2X2_1757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2894_));
OR2X2 OR2X2_1758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2898_));
OR2X2 OR2X2_1759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2902_));
OR2X2 OR2X2_176 ( .A(next_pc_r_1_), .B(next_pc_r_0_), .Y(_abc_44694_new_n1204_));
OR2X2 OR2X2_1760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2906_));
OR2X2 OR2X2_1761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2910_));
OR2X2 OR2X2_1762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2914_));
OR2X2 OR2X2_1763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2918_));
OR2X2 OR2X2_1764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2922_));
OR2X2 OR2X2_1765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2926_));
OR2X2 OR2X2_1766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2930_));
OR2X2 OR2X2_1767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2934_));
OR2X2 OR2X2_1768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2938_));
OR2X2 OR2X2_1769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r25_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2942_));
OR2X2 OR2X2_177 ( .A(_abc_44694_new_n1203_), .B(_abc_44694_new_n1204_), .Y(_abc_44694_new_n1205_));
OR2X2 OR2X2_1770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r25_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2946_));
OR2X2 OR2X2_1771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r25_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2950_));
OR2X2 OR2X2_1772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2829__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r25_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2954_));
OR2X2 OR2X2_1773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2959_));
OR2X2 OR2X2_1774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2961_));
OR2X2 OR2X2_1775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2963_));
OR2X2 OR2X2_1776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2964_));
OR2X2 OR2X2_1777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2966_));
OR2X2 OR2X2_1778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2967_));
OR2X2 OR2X2_1779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2969_));
OR2X2 OR2X2_178 ( .A(_abc_44694_new_n1212_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n1213_));
OR2X2 OR2X2_1780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2970_));
OR2X2 OR2X2_1781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2972_));
OR2X2 OR2X2_1782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2973_));
OR2X2 OR2X2_1783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2975_));
OR2X2 OR2X2_1784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2976_));
OR2X2 OR2X2_1785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2978_));
OR2X2 OR2X2_1786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2979_));
OR2X2 OR2X2_1787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2981_));
OR2X2 OR2X2_1788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2982_));
OR2X2 OR2X2_1789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2984_));
OR2X2 OR2X2_179 ( .A(_abc_44694_new_n1213_), .B(_abc_44694_new_n1209_), .Y(_abc_44694_new_n1214_));
OR2X2 OR2X2_1790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2985_));
OR2X2 OR2X2_1791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2987_));
OR2X2 OR2X2_1792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2988_));
OR2X2 OR2X2_1793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2990_));
OR2X2 OR2X2_1794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2991_));
OR2X2 OR2X2_1795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2993_));
OR2X2 OR2X2_1796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2994_));
OR2X2 OR2X2_1797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2996_));
OR2X2 OR2X2_1798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2997_));
OR2X2 OR2X2_1799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n2999_));
OR2X2 OR2X2_18 ( .A(_abc_44694_new_n707_), .B(_abc_44694_new_n708_), .Y(_abc_44694_new_n709_));
OR2X2 OR2X2_180 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(esr_q_2_), .Y(_abc_44694_new_n1215_));
OR2X2 OR2X2_1800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3000_));
OR2X2 OR2X2_1801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3002_));
OR2X2 OR2X2_1802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3003_));
OR2X2 OR2X2_1803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3005_));
OR2X2 OR2X2_1804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3006_));
OR2X2 OR2X2_1805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3008_));
OR2X2 OR2X2_1806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3009_));
OR2X2 OR2X2_1807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3011_));
OR2X2 OR2X2_1808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3012_));
OR2X2 OR2X2_1809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3014_));
OR2X2 OR2X2_181 ( .A(_abc_44694_new_n1196_), .B(alu_equal_o), .Y(_abc_44694_new_n1221_));
OR2X2 OR2X2_1810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3015_));
OR2X2 OR2X2_1811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3017_));
OR2X2 OR2X2_1812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3018_));
OR2X2 OR2X2_1813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3020_));
OR2X2 OR2X2_1814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3021_));
OR2X2 OR2X2_1815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3023_));
OR2X2 OR2X2_1816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3024_));
OR2X2 OR2X2_1817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3026_));
OR2X2 OR2X2_1818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3027_));
OR2X2 OR2X2_1819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3029_));
OR2X2 OR2X2_182 ( .A(_abc_44694_new_n1224_), .B(_abc_44694_new_n1099_), .Y(_abc_44694_new_n1225_));
OR2X2 OR2X2_1820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3030_));
OR2X2 OR2X2_1821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3032_));
OR2X2 OR2X2_1822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3033_));
OR2X2 OR2X2_1823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3035_));
OR2X2 OR2X2_1824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3036_));
OR2X2 OR2X2_1825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3038_));
OR2X2 OR2X2_1826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3039_));
OR2X2 OR2X2_1827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r24_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3041_));
OR2X2 OR2X2_1828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3042_));
OR2X2 OR2X2_1829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r24_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3044_));
OR2X2 OR2X2_183 ( .A(_abc_44694_new_n1226_), .B(alu_less_than_o), .Y(_abc_44694_new_n1227_));
OR2X2 OR2X2_1830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3045_));
OR2X2 OR2X2_1831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r24_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3047_));
OR2X2 OR2X2_1832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3048_));
OR2X2 OR2X2_1833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r24_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3050_));
OR2X2 OR2X2_1834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3051_));
OR2X2 OR2X2_1835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2958__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r24_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3053_));
OR2X2 OR2X2_1836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n2960__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3054_));
OR2X2 OR2X2_1837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3060_));
OR2X2 OR2X2_1838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3062_));
OR2X2 OR2X2_1839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3064_));
OR2X2 OR2X2_184 ( .A(_abc_44694_new_n1228_), .B(_abc_44694_new_n1197_), .Y(_abc_44694_new_n1229_));
OR2X2 OR2X2_1840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3065_));
OR2X2 OR2X2_1841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3067_));
OR2X2 OR2X2_1842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3068_));
OR2X2 OR2X2_1843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3070_));
OR2X2 OR2X2_1844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3071_));
OR2X2 OR2X2_1845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3073_));
OR2X2 OR2X2_1846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3074_));
OR2X2 OR2X2_1847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3076_));
OR2X2 OR2X2_1848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3077_));
OR2X2 OR2X2_1849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3079_));
OR2X2 OR2X2_185 ( .A(alu_equal_o), .B(alu_less_than_o), .Y(_abc_44694_new_n1235_));
OR2X2 OR2X2_1850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3080_));
OR2X2 OR2X2_1851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3082_));
OR2X2 OR2X2_1852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3083_));
OR2X2 OR2X2_1853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3085_));
OR2X2 OR2X2_1854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3086_));
OR2X2 OR2X2_1855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3088_));
OR2X2 OR2X2_1856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3089_));
OR2X2 OR2X2_1857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3091_));
OR2X2 OR2X2_1858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3092_));
OR2X2 OR2X2_1859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3094_));
OR2X2 OR2X2_186 ( .A(_abc_44694_new_n1166_), .B(_abc_44694_new_n1236_), .Y(_abc_44694_new_n1237_));
OR2X2 OR2X2_1860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3095_));
OR2X2 OR2X2_1861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3097_));
OR2X2 OR2X2_1862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3098_));
OR2X2 OR2X2_1863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3100_));
OR2X2 OR2X2_1864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3101_));
OR2X2 OR2X2_1865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3103_));
OR2X2 OR2X2_1866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3104_));
OR2X2 OR2X2_1867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3106_));
OR2X2 OR2X2_1868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3107_));
OR2X2 OR2X2_1869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3109_));
OR2X2 OR2X2_187 ( .A(_abc_44694_new_n1234_), .B(_abc_44694_new_n1237_), .Y(_abc_44694_new_n1238_));
OR2X2 OR2X2_1870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3110_));
OR2X2 OR2X2_1871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3112_));
OR2X2 OR2X2_1872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3113_));
OR2X2 OR2X2_1873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3115_));
OR2X2 OR2X2_1874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3116_));
OR2X2 OR2X2_1875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3118_));
OR2X2 OR2X2_1876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3119_));
OR2X2 OR2X2_1877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3121_));
OR2X2 OR2X2_1878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3122_));
OR2X2 OR2X2_1879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3124_));
OR2X2 OR2X2_188 ( .A(_abc_44694_new_n1243_), .B(_abc_44694_new_n1220_), .Y(_abc_44694_new_n1244_));
OR2X2 OR2X2_1880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3125_));
OR2X2 OR2X2_1881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3127_));
OR2X2 OR2X2_1882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3128_));
OR2X2 OR2X2_1883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3130_));
OR2X2 OR2X2_1884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3131_));
OR2X2 OR2X2_1885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3133_));
OR2X2 OR2X2_1886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3134_));
OR2X2 OR2X2_1887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3136_));
OR2X2 OR2X2_1888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3137_));
OR2X2 OR2X2_1889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3139_));
OR2X2 OR2X2_189 ( .A(_abc_44694_new_n1173_), .B(_abc_44694_new_n1251_), .Y(_abc_44694_new_n1252_));
OR2X2 OR2X2_1890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3140_));
OR2X2 OR2X2_1891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r23_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3142_));
OR2X2 OR2X2_1892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3143_));
OR2X2 OR2X2_1893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r23_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3145_));
OR2X2 OR2X2_1894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3146_));
OR2X2 OR2X2_1895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r23_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3148_));
OR2X2 OR2X2_1896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3149_));
OR2X2 OR2X2_1897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r23_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3151_));
OR2X2 OR2X2_1898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3152_));
OR2X2 OR2X2_1899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3059__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r23_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3154_));
OR2X2 OR2X2_19 ( .A(_abc_44694_new_n706_), .B(_abc_44694_new_n709_), .Y(_abc_44694_new_n710_));
OR2X2 OR2X2_190 ( .A(_abc_44694_new_n1250_), .B(_abc_44694_new_n1252_), .Y(_abc_44694_new_n1253_));
OR2X2 OR2X2_1900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3061__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3155_));
OR2X2 OR2X2_1901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3159_));
OR2X2 OR2X2_1902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3163_));
OR2X2 OR2X2_1903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3167_));
OR2X2 OR2X2_1904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3171_));
OR2X2 OR2X2_1905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3175_));
OR2X2 OR2X2_1906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3179_));
OR2X2 OR2X2_1907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3183_));
OR2X2 OR2X2_1908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3187_));
OR2X2 OR2X2_1909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3191_));
OR2X2 OR2X2_191 ( .A(alu_equal_o), .B(alu_greater_than_o), .Y(_abc_44694_new_n1254_));
OR2X2 OR2X2_1910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3195_));
OR2X2 OR2X2_1911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3199_));
OR2X2 OR2X2_1912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3203_));
OR2X2 OR2X2_1913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3207_));
OR2X2 OR2X2_1914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3211_));
OR2X2 OR2X2_1915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3215_));
OR2X2 OR2X2_1916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3219_));
OR2X2 OR2X2_1917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3223_));
OR2X2 OR2X2_1918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3227_));
OR2X2 OR2X2_1919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3231_));
OR2X2 OR2X2_192 ( .A(_abc_44694_new_n1174_), .B(_abc_44694_new_n1254_), .Y(_abc_44694_new_n1255_));
OR2X2 OR2X2_1920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3235_));
OR2X2 OR2X2_1921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3239_));
OR2X2 OR2X2_1922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3243_));
OR2X2 OR2X2_1923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3247_));
OR2X2 OR2X2_1924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3251_));
OR2X2 OR2X2_1925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3255_));
OR2X2 OR2X2_1926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3259_));
OR2X2 OR2X2_1927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3263_));
OR2X2 OR2X2_1928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3267_));
OR2X2 OR2X2_1929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r22_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3271_));
OR2X2 OR2X2_193 ( .A(alu_equal_o), .B(alu_greater_than_signed_o), .Y(_abc_44694_new_n1258_));
OR2X2 OR2X2_1930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r22_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3275_));
OR2X2 OR2X2_1931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r22_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3279_));
OR2X2 OR2X2_1932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3158__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r22_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3283_));
OR2X2 OR2X2_1933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3289_));
OR2X2 OR2X2_1934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3293_));
OR2X2 OR2X2_1935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3297_));
OR2X2 OR2X2_1936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3301_));
OR2X2 OR2X2_1937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3305_));
OR2X2 OR2X2_1938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3309_));
OR2X2 OR2X2_1939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3313_));
OR2X2 OR2X2_194 ( .A(_abc_44694_new_n1257_), .B(_abc_44694_new_n1259_), .Y(_abc_44694_new_n1260_));
OR2X2 OR2X2_1940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3317_));
OR2X2 OR2X2_1941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3321_));
OR2X2 OR2X2_1942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3325_));
OR2X2 OR2X2_1943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3329_));
OR2X2 OR2X2_1944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3333_));
OR2X2 OR2X2_1945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3337_));
OR2X2 OR2X2_1946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3341_));
OR2X2 OR2X2_1947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3345_));
OR2X2 OR2X2_1948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3349_));
OR2X2 OR2X2_1949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3353_));
OR2X2 OR2X2_195 ( .A(_abc_44694_new_n1261_), .B(_abc_44694_new_n1219_), .Y(_abc_44694_new_n1262_));
OR2X2 OR2X2_1950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3357_));
OR2X2 OR2X2_1951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3361_));
OR2X2 OR2X2_1952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3365_));
OR2X2 OR2X2_1953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3369_));
OR2X2 OR2X2_1954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3373_));
OR2X2 OR2X2_1955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3377_));
OR2X2 OR2X2_1956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3381_));
OR2X2 OR2X2_1957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3385_));
OR2X2 OR2X2_1958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3389_));
OR2X2 OR2X2_1959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3393_));
OR2X2 OR2X2_196 ( .A(_abc_44694_new_n1264_), .B(_abc_44694_new_n1019__bF_buf2), .Y(_abc_44694_new_n1265_));
OR2X2 OR2X2_1960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3397_));
OR2X2 OR2X2_1961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r21_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3401_));
OR2X2 OR2X2_1962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r21_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3405_));
OR2X2 OR2X2_1963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r21_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3409_));
OR2X2 OR2X2_1964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3288__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r21_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3413_));
OR2X2 OR2X2_1965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3418_));
OR2X2 OR2X2_1966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3420_));
OR2X2 OR2X2_1967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3422_));
OR2X2 OR2X2_1968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3423_));
OR2X2 OR2X2_1969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3425_));
OR2X2 OR2X2_197 ( .A(_abc_44694_new_n1263_), .B(_abc_44694_new_n1265_), .Y(_abc_44694_new_n1266_));
OR2X2 OR2X2_1970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3426_));
OR2X2 OR2X2_1971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3428_));
OR2X2 OR2X2_1972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3429_));
OR2X2 OR2X2_1973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3431_));
OR2X2 OR2X2_1974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3432_));
OR2X2 OR2X2_1975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3434_));
OR2X2 OR2X2_1976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3435_));
OR2X2 OR2X2_1977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3437_));
OR2X2 OR2X2_1978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3438_));
OR2X2 OR2X2_1979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3440_));
OR2X2 OR2X2_198 ( .A(_abc_44694_new_n1021_), .B(esr_q_9_), .Y(_abc_44694_new_n1267_));
OR2X2 OR2X2_1980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3441_));
OR2X2 OR2X2_1981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3443_));
OR2X2 OR2X2_1982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3444_));
OR2X2 OR2X2_1983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3446_));
OR2X2 OR2X2_1984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3447_));
OR2X2 OR2X2_1985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3449_));
OR2X2 OR2X2_1986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3450_));
OR2X2 OR2X2_1987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3452_));
OR2X2 OR2X2_1988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3453_));
OR2X2 OR2X2_1989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3455_));
OR2X2 OR2X2_199 ( .A(_abc_44694_new_n1262_), .B(_abc_44694_new_n1011_), .Y(_abc_44694_new_n1270_));
OR2X2 OR2X2_1990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3456_));
OR2X2 OR2X2_1991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3458_));
OR2X2 OR2X2_1992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3459_));
OR2X2 OR2X2_1993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3461_));
OR2X2 OR2X2_1994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3462_));
OR2X2 OR2X2_1995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3464_));
OR2X2 OR2X2_1996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3465_));
OR2X2 OR2X2_1997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3467_));
OR2X2 OR2X2_1998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3468_));
OR2X2 OR2X2_1999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3470_));
OR2X2 OR2X2_2 ( .A(_abc_44694_new_n644_), .B(_abc_44694_new_n652_), .Y(_abc_44694_new_n653_));
OR2X2 OR2X2_20 ( .A(_abc_44694_new_n673__bF_buf3), .B(_abc_44694_new_n710_), .Y(_abc_44694_new_n711_));
OR2X2 OR2X2_200 ( .A(_abc_44694_new_n1269_), .B(_abc_44694_new_n1275_), .Y(_abc_44694_new_n1276_));
OR2X2 OR2X2_2000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3471_));
OR2X2 OR2X2_2001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3473_));
OR2X2 OR2X2_2002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3474_));
OR2X2 OR2X2_2003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3476_));
OR2X2 OR2X2_2004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3477_));
OR2X2 OR2X2_2005 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3479_));
OR2X2 OR2X2_2006 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3480_));
OR2X2 OR2X2_2007 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3482_));
OR2X2 OR2X2_2008 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3483_));
OR2X2 OR2X2_2009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3485_));
OR2X2 OR2X2_201 ( .A(_abc_44694_new_n1282_), .B(_abc_44694_new_n1283_), .Y(_abc_44694_new_n1284_));
OR2X2 OR2X2_2010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3486_));
OR2X2 OR2X2_2011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3488_));
OR2X2 OR2X2_2012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3489_));
OR2X2 OR2X2_2013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3491_));
OR2X2 OR2X2_2014 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3492_));
OR2X2 OR2X2_2015 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3494_));
OR2X2 OR2X2_2016 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3495_));
OR2X2 OR2X2_2017 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3497_));
OR2X2 OR2X2_2018 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3498_));
OR2X2 OR2X2_2019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r20_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3500_));
OR2X2 OR2X2_202 ( .A(_abc_44694_new_n1285_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n1286_));
OR2X2 OR2X2_2020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3501_));
OR2X2 OR2X2_2021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r20_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3503_));
OR2X2 OR2X2_2022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3504_));
OR2X2 OR2X2_2023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r20_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3506_));
OR2X2 OR2X2_2024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3507_));
OR2X2 OR2X2_2025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r20_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3509_));
OR2X2 OR2X2_2026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3510_));
OR2X2 OR2X2_2027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3417__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r20_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3512_));
OR2X2 OR2X2_2028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3419__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3513_));
OR2X2 OR2X2_2029 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3518_));
OR2X2 OR2X2_203 ( .A(_abc_44694_new_n1281_), .B(_abc_44694_new_n1286_), .Y(_abc_44694_new_n1287_));
OR2X2 OR2X2_2030 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3520_));
OR2X2 OR2X2_2031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3522_));
OR2X2 OR2X2_2032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3523_));
OR2X2 OR2X2_2033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3525_));
OR2X2 OR2X2_2034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3526_));
OR2X2 OR2X2_2035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3528_));
OR2X2 OR2X2_2036 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3529_));
OR2X2 OR2X2_2037 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3531_));
OR2X2 OR2X2_2038 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3532_));
OR2X2 OR2X2_2039 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3534_));
OR2X2 OR2X2_204 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(esr_q_9_), .Y(_abc_44694_new_n1288_));
OR2X2 OR2X2_2040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3535_));
OR2X2 OR2X2_2041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3537_));
OR2X2 OR2X2_2042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3538_));
OR2X2 OR2X2_2043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3540_));
OR2X2 OR2X2_2044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3541_));
OR2X2 OR2X2_2045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3543_));
OR2X2 OR2X2_2046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3544_));
OR2X2 OR2X2_2047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3546_));
OR2X2 OR2X2_2048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3547_));
OR2X2 OR2X2_2049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3549_));
OR2X2 OR2X2_205 ( .A(_abc_44694_new_n1291_), .B(_abc_44694_new_n1292_), .Y(_abc_44694_new_n1293_));
OR2X2 OR2X2_2050 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3550_));
OR2X2 OR2X2_2051 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3552_));
OR2X2 OR2X2_2052 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3553_));
OR2X2 OR2X2_2053 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3555_));
OR2X2 OR2X2_2054 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3556_));
OR2X2 OR2X2_2055 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3558_));
OR2X2 OR2X2_2056 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3559_));
OR2X2 OR2X2_2057 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3561_));
OR2X2 OR2X2_2058 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3562_));
OR2X2 OR2X2_2059 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3564_));
OR2X2 OR2X2_206 ( .A(alu_c_i), .B(alu_c_update_o), .Y(_abc_44694_new_n1295_));
OR2X2 OR2X2_2060 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3565_));
OR2X2 OR2X2_2061 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3567_));
OR2X2 OR2X2_2062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3568_));
OR2X2 OR2X2_2063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3570_));
OR2X2 OR2X2_2064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3571_));
OR2X2 OR2X2_2065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3573_));
OR2X2 OR2X2_2066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3574_));
OR2X2 OR2X2_2067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3576_));
OR2X2 OR2X2_2068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3577_));
OR2X2 OR2X2_2069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3579_));
OR2X2 OR2X2_207 ( .A(_abc_44694_new_n1296_), .B(alu_c_o), .Y(_abc_44694_new_n1297_));
OR2X2 OR2X2_2070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3580_));
OR2X2 OR2X2_2071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3582_));
OR2X2 OR2X2_2072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3583_));
OR2X2 OR2X2_2073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3585_));
OR2X2 OR2X2_2074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3586_));
OR2X2 OR2X2_2075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3588_));
OR2X2 OR2X2_2076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3589_));
OR2X2 OR2X2_2077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3591_));
OR2X2 OR2X2_2078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3592_));
OR2X2 OR2X2_2079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3594_));
OR2X2 OR2X2_208 ( .A(_abc_44694_new_n1019__bF_buf1), .B(_abc_44694_new_n1298_), .Y(_abc_44694_new_n1299_));
OR2X2 OR2X2_2080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3595_));
OR2X2 OR2X2_2081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3597_));
OR2X2 OR2X2_2082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3598_));
OR2X2 OR2X2_2083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r19_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3600_));
OR2X2 OR2X2_2084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3601_));
OR2X2 OR2X2_2085 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r19_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3603_));
OR2X2 OR2X2_2086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3604_));
OR2X2 OR2X2_2087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r19_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3606_));
OR2X2 OR2X2_2088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3607_));
OR2X2 OR2X2_2089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r19_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3609_));
OR2X2 OR2X2_209 ( .A(_abc_44694_new_n1021_), .B(esr_q_10_), .Y(_abc_44694_new_n1300_));
OR2X2 OR2X2_2090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3610_));
OR2X2 OR2X2_2091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3517__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r19_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3612_));
OR2X2 OR2X2_2092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3519__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3613_));
OR2X2 OR2X2_2093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3617_));
OR2X2 OR2X2_2094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3619_));
OR2X2 OR2X2_2095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3621_));
OR2X2 OR2X2_2096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3622_));
OR2X2 OR2X2_2097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3624_));
OR2X2 OR2X2_2098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3625_));
OR2X2 OR2X2_2099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3627_));
OR2X2 OR2X2_21 ( .A(_abc_44694_new_n713_), .B(_abc_44694_new_n699_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_1_));
OR2X2 OR2X2_210 ( .A(_abc_44694_new_n1301_), .B(_abc_44694_new_n970_), .Y(_abc_44694_new_n1302_));
OR2X2 OR2X2_2100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3628_));
OR2X2 OR2X2_2101 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3630_));
OR2X2 OR2X2_2102 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3631_));
OR2X2 OR2X2_2103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3633_));
OR2X2 OR2X2_2104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3634_));
OR2X2 OR2X2_2105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3636_));
OR2X2 OR2X2_2106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3637_));
OR2X2 OR2X2_2107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3639_));
OR2X2 OR2X2_2108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3640_));
OR2X2 OR2X2_2109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3642_));
OR2X2 OR2X2_211 ( .A(_abc_44694_new_n1011_), .B(_abc_44694_new_n1298_), .Y(_abc_44694_new_n1303_));
OR2X2 OR2X2_2110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3643_));
OR2X2 OR2X2_2111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3645_));
OR2X2 OR2X2_2112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3646_));
OR2X2 OR2X2_2113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3648_));
OR2X2 OR2X2_2114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3649_));
OR2X2 OR2X2_2115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3651_));
OR2X2 OR2X2_2116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3652_));
OR2X2 OR2X2_2117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3654_));
OR2X2 OR2X2_2118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3655_));
OR2X2 OR2X2_2119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3657_));
OR2X2 OR2X2_212 ( .A(_abc_44694_new_n1307_), .B(_abc_44694_new_n1017_), .Y(_abc_44694_new_n1308_));
OR2X2 OR2X2_2120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3658_));
OR2X2 OR2X2_2121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3660_));
OR2X2 OR2X2_2122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3661_));
OR2X2 OR2X2_2123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3663_));
OR2X2 OR2X2_2124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3664_));
OR2X2 OR2X2_2125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3666_));
OR2X2 OR2X2_2126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3667_));
OR2X2 OR2X2_2127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3669_));
OR2X2 OR2X2_2128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3670_));
OR2X2 OR2X2_2129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3672_));
OR2X2 OR2X2_213 ( .A(_abc_44694_new_n1310_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n1311_));
OR2X2 OR2X2_2130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3673_));
OR2X2 OR2X2_2131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3675_));
OR2X2 OR2X2_2132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3676_));
OR2X2 OR2X2_2133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3678_));
OR2X2 OR2X2_2134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3679_));
OR2X2 OR2X2_2135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3681_));
OR2X2 OR2X2_2136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3682_));
OR2X2 OR2X2_2137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3684_));
OR2X2 OR2X2_2138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3685_));
OR2X2 OR2X2_2139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3687_));
OR2X2 OR2X2_214 ( .A(_abc_44694_new_n1311_), .B(_abc_44694_new_n1294_), .Y(_abc_44694_new_n1312_));
OR2X2 OR2X2_2140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3688_));
OR2X2 OR2X2_2141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3690_));
OR2X2 OR2X2_2142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3691_));
OR2X2 OR2X2_2143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3693_));
OR2X2 OR2X2_2144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3694_));
OR2X2 OR2X2_2145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3696_));
OR2X2 OR2X2_2146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3697_));
OR2X2 OR2X2_2147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r18_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3699_));
OR2X2 OR2X2_2148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3700_));
OR2X2 OR2X2_2149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r18_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3702_));
OR2X2 OR2X2_215 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(esr_q_10_), .Y(_abc_44694_new_n1313_));
OR2X2 OR2X2_2150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3703_));
OR2X2 OR2X2_2151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r18_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3705_));
OR2X2 OR2X2_2152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3706_));
OR2X2 OR2X2_2153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r18_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3708_));
OR2X2 OR2X2_2154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3709_));
OR2X2 OR2X2_2155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3616__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r18_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3711_));
OR2X2 OR2X2_2156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3618__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3712_));
OR2X2 OR2X2_2157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3716_));
OR2X2 OR2X2_2158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3718_));
OR2X2 OR2X2_2159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3720_));
OR2X2 OR2X2_216 ( .A(_abc_44694_new_n1318_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n1319_));
OR2X2 OR2X2_2160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3721_));
OR2X2 OR2X2_2161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3723_));
OR2X2 OR2X2_2162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3724_));
OR2X2 OR2X2_2163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3726_));
OR2X2 OR2X2_2164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3727_));
OR2X2 OR2X2_2165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3729_));
OR2X2 OR2X2_2166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3730_));
OR2X2 OR2X2_2167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3732_));
OR2X2 OR2X2_2168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3733_));
OR2X2 OR2X2_2169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3735_));
OR2X2 OR2X2_217 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(sr_q_2_), .Y(_abc_44694_new_n1320_));
OR2X2 OR2X2_2170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3736_));
OR2X2 OR2X2_2171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3738_));
OR2X2 OR2X2_2172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3739_));
OR2X2 OR2X2_2173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3741_));
OR2X2 OR2X2_2174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3742_));
OR2X2 OR2X2_2175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3744_));
OR2X2 OR2X2_2176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3745_));
OR2X2 OR2X2_2177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3747_));
OR2X2 OR2X2_2178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3748_));
OR2X2 OR2X2_2179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3750_));
OR2X2 OR2X2_218 ( .A(_abc_44694_new_n1323_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n1324_));
OR2X2 OR2X2_2180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3751_));
OR2X2 OR2X2_2181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3753_));
OR2X2 OR2X2_2182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3754_));
OR2X2 OR2X2_2183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3756_));
OR2X2 OR2X2_2184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3757_));
OR2X2 OR2X2_2185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3759_));
OR2X2 OR2X2_2186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3760_));
OR2X2 OR2X2_2187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3762_));
OR2X2 OR2X2_2188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3763_));
OR2X2 OR2X2_2189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3765_));
OR2X2 OR2X2_219 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(sr_q_9_), .Y(_abc_44694_new_n1325_));
OR2X2 OR2X2_2190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3766_));
OR2X2 OR2X2_2191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3768_));
OR2X2 OR2X2_2192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3769_));
OR2X2 OR2X2_2193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3771_));
OR2X2 OR2X2_2194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3772_));
OR2X2 OR2X2_2195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3774_));
OR2X2 OR2X2_2196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3775_));
OR2X2 OR2X2_2197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3777_));
OR2X2 OR2X2_2198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3778_));
OR2X2 OR2X2_2199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3780_));
OR2X2 OR2X2_22 ( .A(_abc_44694_new_n717_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n718_));
OR2X2 OR2X2_220 ( .A(_abc_44694_new_n1331_), .B(_abc_44694_new_n1328_), .Y(_abc_44694_new_n1332_));
OR2X2 OR2X2_2200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3781_));
OR2X2 OR2X2_2201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3783_));
OR2X2 OR2X2_2202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3784_));
OR2X2 OR2X2_2203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3786_));
OR2X2 OR2X2_2204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3787_));
OR2X2 OR2X2_2205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3789_));
OR2X2 OR2X2_2206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3790_));
OR2X2 OR2X2_2207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3792_));
OR2X2 OR2X2_2208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3793_));
OR2X2 OR2X2_2209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3795_));
OR2X2 OR2X2_221 ( .A(_abc_44694_new_n1121_), .B(_abc_44694_new_n1176_), .Y(_abc_44694_new_n1337_));
OR2X2 OR2X2_2210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3796_));
OR2X2 OR2X2_2211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r17_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3798_));
OR2X2 OR2X2_2212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3799_));
OR2X2 OR2X2_2213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r17_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3801_));
OR2X2 OR2X2_2214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3802_));
OR2X2 OR2X2_2215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r17_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3804_));
OR2X2 OR2X2_2216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3805_));
OR2X2 OR2X2_2217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r17_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3807_));
OR2X2 OR2X2_2218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3808_));
OR2X2 OR2X2_2219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3715__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r17_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3810_));
OR2X2 OR2X2_222 ( .A(_abc_44694_new_n1337__bF_buf4), .B(_abc_44694_new_n1336_), .Y(_abc_44694_new_n1338_));
OR2X2 OR2X2_2220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3717__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3811_));
OR2X2 OR2X2_2221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3814_));
OR2X2 OR2X2_2222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3816_));
OR2X2 OR2X2_2223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3818_));
OR2X2 OR2X2_2224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3819_));
OR2X2 OR2X2_2225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3821_));
OR2X2 OR2X2_2226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3822_));
OR2X2 OR2X2_2227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3824_));
OR2X2 OR2X2_2228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3825_));
OR2X2 OR2X2_2229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3827_));
OR2X2 OR2X2_223 ( .A(_abc_44694_new_n1335_), .B(_abc_44694_new_n1338_), .Y(_abc_44694_new_n1339_));
OR2X2 OR2X2_2230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3828_));
OR2X2 OR2X2_2231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3830_));
OR2X2 OR2X2_2232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3831_));
OR2X2 OR2X2_2233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3833_));
OR2X2 OR2X2_2234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3834_));
OR2X2 OR2X2_2235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3836_));
OR2X2 OR2X2_2236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3837_));
OR2X2 OR2X2_2237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3839_));
OR2X2 OR2X2_2238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3840_));
OR2X2 OR2X2_2239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3842_));
OR2X2 OR2X2_224 ( .A(_abc_44694_new_n1340__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rb_o_0_), .Y(_abc_44694_new_n1341_));
OR2X2 OR2X2_2240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3843_));
OR2X2 OR2X2_2241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3845_));
OR2X2 OR2X2_2242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3846_));
OR2X2 OR2X2_2243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3848_));
OR2X2 OR2X2_2244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3849_));
OR2X2 OR2X2_2245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3851_));
OR2X2 OR2X2_2246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3852_));
OR2X2 OR2X2_2247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3854_));
OR2X2 OR2X2_2248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3855_));
OR2X2 OR2X2_2249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3857_));
OR2X2 OR2X2_225 ( .A(_abc_44694_new_n1348__bF_buf5), .B(epc_q_0_), .Y(_abc_44694_new_n1349_));
OR2X2 OR2X2_2250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3858_));
OR2X2 OR2X2_2251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3860_));
OR2X2 OR2X2_2252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3861_));
OR2X2 OR2X2_2253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3863_));
OR2X2 OR2X2_2254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3864_));
OR2X2 OR2X2_2255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3866_));
OR2X2 OR2X2_2256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3867_));
OR2X2 OR2X2_2257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3869_));
OR2X2 OR2X2_2258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3870_));
OR2X2 OR2X2_2259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3872_));
OR2X2 OR2X2_226 ( .A(_abc_44694_new_n1343_), .B(_abc_44694_new_n1354_), .Y(_abc_44694_new_n1355_));
OR2X2 OR2X2_2260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3873_));
OR2X2 OR2X2_2261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3875_));
OR2X2 OR2X2_2262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3876_));
OR2X2 OR2X2_2263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3878_));
OR2X2 OR2X2_2264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3879_));
OR2X2 OR2X2_2265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3881_));
OR2X2 OR2X2_2266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3882_));
OR2X2 OR2X2_2267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3884_));
OR2X2 OR2X2_2268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3885_));
OR2X2 OR2X2_2269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3887_));
OR2X2 OR2X2_227 ( .A(_abc_44694_new_n1210__bF_buf1), .B(next_pc_r_0_), .Y(_abc_44694_new_n1357_));
OR2X2 OR2X2_2270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3888_));
OR2X2 OR2X2_2271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3890_));
OR2X2 OR2X2_2272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3891_));
OR2X2 OR2X2_2273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3893_));
OR2X2 OR2X2_2274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3894_));
OR2X2 OR2X2_2275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r16_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3896_));
OR2X2 OR2X2_2276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3897_));
OR2X2 OR2X2_2277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r16_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3899_));
OR2X2 OR2X2_2278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3900_));
OR2X2 OR2X2_2279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r16_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3902_));
OR2X2 OR2X2_228 ( .A(_abc_44694_new_n1356_), .B(_abc_44694_new_n1357_), .Y(_abc_44694_new_n1358_));
OR2X2 OR2X2_2280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3903_));
OR2X2 OR2X2_2281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r16_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3905_));
OR2X2 OR2X2_2282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3906_));
OR2X2 OR2X2_2283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3813__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r16_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3908_));
OR2X2 OR2X2_2284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3815__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3909_));
OR2X2 OR2X2_2285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3914_));
OR2X2 OR2X2_2286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3918_));
OR2X2 OR2X2_2287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3922_));
OR2X2 OR2X2_2288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3926_));
OR2X2 OR2X2_2289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3930_));
OR2X2 OR2X2_229 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_0_), .Y(_abc_44694_new_n1359_));
OR2X2 OR2X2_2290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3934_));
OR2X2 OR2X2_2291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3938_));
OR2X2 OR2X2_2292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3942_));
OR2X2 OR2X2_2293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3946_));
OR2X2 OR2X2_2294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3950_));
OR2X2 OR2X2_2295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3954_));
OR2X2 OR2X2_2296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3958_));
OR2X2 OR2X2_2297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3962_));
OR2X2 OR2X2_2298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3966_));
OR2X2 OR2X2_2299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3970_));
OR2X2 OR2X2_23 ( .A(_abc_44694_new_n718_), .B(_abc_44694_new_n716_), .Y(_abc_44694_new_n719_));
OR2X2 OR2X2_230 ( .A(_abc_44694_new_n1337__bF_buf2), .B(_abc_44694_new_n1363_), .Y(_abc_44694_new_n1364_));
OR2X2 OR2X2_2300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3974_));
OR2X2 OR2X2_2301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3978_));
OR2X2 OR2X2_2302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3982_));
OR2X2 OR2X2_2303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3986_));
OR2X2 OR2X2_2304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3990_));
OR2X2 OR2X2_2305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3994_));
OR2X2 OR2X2_2306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n3998_));
OR2X2 OR2X2_2307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4002_));
OR2X2 OR2X2_2308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4006_));
OR2X2 OR2X2_2309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4010_));
OR2X2 OR2X2_231 ( .A(_abc_44694_new_n1362_), .B(_abc_44694_new_n1364_), .Y(_abc_44694_new_n1365_));
OR2X2 OR2X2_2310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4014_));
OR2X2 OR2X2_2311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4018_));
OR2X2 OR2X2_2312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4022_));
OR2X2 OR2X2_2313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r15_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4026_));
OR2X2 OR2X2_2314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r15_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4030_));
OR2X2 OR2X2_2315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r15_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4034_));
OR2X2 OR2X2_2316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n3913__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r15_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4038_));
OR2X2 OR2X2_2317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4043_));
OR2X2 OR2X2_2318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4045_));
OR2X2 OR2X2_2319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4047_));
OR2X2 OR2X2_232 ( .A(_abc_44694_new_n1340__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_1_), .Y(_abc_44694_new_n1366_));
OR2X2 OR2X2_2320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4048_));
OR2X2 OR2X2_2321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4050_));
OR2X2 OR2X2_2322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4051_));
OR2X2 OR2X2_2323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4053_));
OR2X2 OR2X2_2324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4054_));
OR2X2 OR2X2_2325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4056_));
OR2X2 OR2X2_2326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4057_));
OR2X2 OR2X2_2327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4059_));
OR2X2 OR2X2_2328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4060_));
OR2X2 OR2X2_2329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4062_));
OR2X2 OR2X2_233 ( .A(_abc_44694_new_n1348__bF_buf3), .B(epc_q_1_), .Y(_abc_44694_new_n1369_));
OR2X2 OR2X2_2330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4063_));
OR2X2 OR2X2_2331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4065_));
OR2X2 OR2X2_2332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4066_));
OR2X2 OR2X2_2333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4068_));
OR2X2 OR2X2_2334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4069_));
OR2X2 OR2X2_2335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4071_));
OR2X2 OR2X2_2336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4072_));
OR2X2 OR2X2_2337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4074_));
OR2X2 OR2X2_2338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4075_));
OR2X2 OR2X2_2339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4077_));
OR2X2 OR2X2_234 ( .A(_abc_44694_new_n1368_), .B(_abc_44694_new_n1374_), .Y(_abc_44694_new_n1375_));
OR2X2 OR2X2_2340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4078_));
OR2X2 OR2X2_2341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4080_));
OR2X2 OR2X2_2342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4081_));
OR2X2 OR2X2_2343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4083_));
OR2X2 OR2X2_2344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4084_));
OR2X2 OR2X2_2345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4086_));
OR2X2 OR2X2_2346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4087_));
OR2X2 OR2X2_2347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4089_));
OR2X2 OR2X2_2348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4090_));
OR2X2 OR2X2_2349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4092_));
OR2X2 OR2X2_235 ( .A(_abc_44694_new_n1210__bF_buf0), .B(next_pc_r_1_), .Y(_abc_44694_new_n1377_));
OR2X2 OR2X2_2350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4093_));
OR2X2 OR2X2_2351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4095_));
OR2X2 OR2X2_2352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4096_));
OR2X2 OR2X2_2353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4098_));
OR2X2 OR2X2_2354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4099_));
OR2X2 OR2X2_2355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4101_));
OR2X2 OR2X2_2356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4102_));
OR2X2 OR2X2_2357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4104_));
OR2X2 OR2X2_2358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4105_));
OR2X2 OR2X2_2359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4107_));
OR2X2 OR2X2_236 ( .A(_abc_44694_new_n1376_), .B(_abc_44694_new_n1377_), .Y(_abc_44694_new_n1378_));
OR2X2 OR2X2_2360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4108_));
OR2X2 OR2X2_2361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4110_));
OR2X2 OR2X2_2362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4111_));
OR2X2 OR2X2_2363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4113_));
OR2X2 OR2X2_2364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4114_));
OR2X2 OR2X2_2365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4116_));
OR2X2 OR2X2_2366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4117_));
OR2X2 OR2X2_2367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4119_));
OR2X2 OR2X2_2368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4120_));
OR2X2 OR2X2_2369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4122_));
OR2X2 OR2X2_237 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(epc_q_1_), .Y(_abc_44694_new_n1379_));
OR2X2 OR2X2_2370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4123_));
OR2X2 OR2X2_2371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r14_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4125_));
OR2X2 OR2X2_2372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4126_));
OR2X2 OR2X2_2373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r14_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4128_));
OR2X2 OR2X2_2374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4129_));
OR2X2 OR2X2_2375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r14_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4131_));
OR2X2 OR2X2_2376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4132_));
OR2X2 OR2X2_2377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r14_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4134_));
OR2X2 OR2X2_2378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4135_));
OR2X2 OR2X2_2379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4042__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r14_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4137_));
OR2X2 OR2X2_238 ( .A(_abc_44694_new_n1348__bF_buf0), .B(epc_q_2_), .Y(_abc_44694_new_n1386_));
OR2X2 OR2X2_2380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4044__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4138_));
OR2X2 OR2X2_2381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4141_));
OR2X2 OR2X2_2382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4143_));
OR2X2 OR2X2_2383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4145_));
OR2X2 OR2X2_2384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4146_));
OR2X2 OR2X2_2385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4148_));
OR2X2 OR2X2_2386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4149_));
OR2X2 OR2X2_2387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4151_));
OR2X2 OR2X2_2388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4152_));
OR2X2 OR2X2_2389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4154_));
OR2X2 OR2X2_239 ( .A(_abc_44694_new_n1334__bF_buf2), .B(_abc_44694_new_n1387_), .Y(_abc_44694_new_n1388_));
OR2X2 OR2X2_2390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4155_));
OR2X2 OR2X2_2391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4157_));
OR2X2 OR2X2_2392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4158_));
OR2X2 OR2X2_2393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4160_));
OR2X2 OR2X2_2394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4161_));
OR2X2 OR2X2_2395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4163_));
OR2X2 OR2X2_2396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4164_));
OR2X2 OR2X2_2397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4166_));
OR2X2 OR2X2_2398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4167_));
OR2X2 OR2X2_2399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4169_));
OR2X2 OR2X2_24 ( .A(_abc_44694_new_n720_), .B(_abc_44694_new_n721_), .Y(_abc_44694_new_n722_));
OR2X2 OR2X2_240 ( .A(_abc_44694_new_n1337__bF_buf1), .B(_abc_44694_new_n1390_), .Y(_abc_44694_new_n1391_));
OR2X2 OR2X2_2400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4170_));
OR2X2 OR2X2_2401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4172_));
OR2X2 OR2X2_2402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4173_));
OR2X2 OR2X2_2403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4175_));
OR2X2 OR2X2_2404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4176_));
OR2X2 OR2X2_2405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4178_));
OR2X2 OR2X2_2406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4179_));
OR2X2 OR2X2_2407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4181_));
OR2X2 OR2X2_2408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4182_));
OR2X2 OR2X2_2409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4184_));
OR2X2 OR2X2_241 ( .A(_abc_44694_new_n1389_), .B(_abc_44694_new_n1391_), .Y(_abc_44694_new_n1392_));
OR2X2 OR2X2_2410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4185_));
OR2X2 OR2X2_2411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4187_));
OR2X2 OR2X2_2412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4188_));
OR2X2 OR2X2_2413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4190_));
OR2X2 OR2X2_2414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4191_));
OR2X2 OR2X2_2415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4193_));
OR2X2 OR2X2_2416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4194_));
OR2X2 OR2X2_2417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4196_));
OR2X2 OR2X2_2418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4197_));
OR2X2 OR2X2_2419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4199_));
OR2X2 OR2X2_242 ( .A(_abc_44694_new_n1396_), .B(_abc_44694_new_n1398_), .Y(_abc_44694_new_n1399_));
OR2X2 OR2X2_2420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4200_));
OR2X2 OR2X2_2421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4202_));
OR2X2 OR2X2_2422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4203_));
OR2X2 OR2X2_2423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4205_));
OR2X2 OR2X2_2424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4206_));
OR2X2 OR2X2_2425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4208_));
OR2X2 OR2X2_2426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4209_));
OR2X2 OR2X2_2427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4211_));
OR2X2 OR2X2_2428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4212_));
OR2X2 OR2X2_2429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4214_));
OR2X2 OR2X2_243 ( .A(_abc_44694_new_n1340__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_2_), .Y(_abc_44694_new_n1401_));
OR2X2 OR2X2_2430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4215_));
OR2X2 OR2X2_2431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4217_));
OR2X2 OR2X2_2432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4218_));
OR2X2 OR2X2_2433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4220_));
OR2X2 OR2X2_2434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4221_));
OR2X2 OR2X2_2435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r13_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4223_));
OR2X2 OR2X2_2436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4224_));
OR2X2 OR2X2_2437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r13_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4226_));
OR2X2 OR2X2_2438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4227_));
OR2X2 OR2X2_2439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r13_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4229_));
OR2X2 OR2X2_244 ( .A(alu_op_r_0_), .B(pc_q_2_), .Y(_abc_44694_new_n1402_));
OR2X2 OR2X2_2440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4230_));
OR2X2 OR2X2_2441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r13_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4232_));
OR2X2 OR2X2_2442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4233_));
OR2X2 OR2X2_2443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4140__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r13_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4235_));
OR2X2 OR2X2_2444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4142__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4236_));
OR2X2 OR2X2_2445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4240_));
OR2X2 OR2X2_2446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4242_));
OR2X2 OR2X2_2447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4244_));
OR2X2 OR2X2_2448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4245_));
OR2X2 OR2X2_2449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4247_));
OR2X2 OR2X2_245 ( .A(_abc_44694_new_n1337__bF_buf0), .B(_abc_44694_new_n1407_), .Y(_abc_44694_new_n1408_));
OR2X2 OR2X2_2450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4248_));
OR2X2 OR2X2_2451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4250_));
OR2X2 OR2X2_2452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4251_));
OR2X2 OR2X2_2453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4253_));
OR2X2 OR2X2_2454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4254_));
OR2X2 OR2X2_2455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4256_));
OR2X2 OR2X2_2456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4257_));
OR2X2 OR2X2_2457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4259_));
OR2X2 OR2X2_2458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4260_));
OR2X2 OR2X2_2459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4262_));
OR2X2 OR2X2_246 ( .A(_abc_44694_new_n1406_), .B(_abc_44694_new_n1408_), .Y(_abc_44694_new_n1409_));
OR2X2 OR2X2_2460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4263_));
OR2X2 OR2X2_2461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4265_));
OR2X2 OR2X2_2462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4266_));
OR2X2 OR2X2_2463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4268_));
OR2X2 OR2X2_2464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4269_));
OR2X2 OR2X2_2465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4271_));
OR2X2 OR2X2_2466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4272_));
OR2X2 OR2X2_2467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4274_));
OR2X2 OR2X2_2468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4275_));
OR2X2 OR2X2_2469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4277_));
OR2X2 OR2X2_247 ( .A(_abc_44694_new_n1400__bF_buf4), .B(_abc_44694_new_n1410_), .Y(_abc_44694_new_n1411_));
OR2X2 OR2X2_2470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4278_));
OR2X2 OR2X2_2471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4280_));
OR2X2 OR2X2_2472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4281_));
OR2X2 OR2X2_2473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4283_));
OR2X2 OR2X2_2474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4284_));
OR2X2 OR2X2_2475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4286_));
OR2X2 OR2X2_2476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4287_));
OR2X2 OR2X2_2477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4289_));
OR2X2 OR2X2_2478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4290_));
OR2X2 OR2X2_2479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4292_));
OR2X2 OR2X2_248 ( .A(_abc_44694_new_n1399__bF_buf3), .B(_abc_44694_new_n1412_), .Y(_abc_44694_new_n1413_));
OR2X2 OR2X2_2480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4293_));
OR2X2 OR2X2_2481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4295_));
OR2X2 OR2X2_2482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4296_));
OR2X2 OR2X2_2483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4298_));
OR2X2 OR2X2_2484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4299_));
OR2X2 OR2X2_2485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4301_));
OR2X2 OR2X2_2486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4302_));
OR2X2 OR2X2_2487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4304_));
OR2X2 OR2X2_2488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4305_));
OR2X2 OR2X2_2489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4307_));
OR2X2 OR2X2_249 ( .A(_abc_44694_new_n1414_), .B(_abc_44694_new_n1278__bF_buf0), .Y(_abc_44694_new_n1415_));
OR2X2 OR2X2_2490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4308_));
OR2X2 OR2X2_2491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4310_));
OR2X2 OR2X2_2492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4311_));
OR2X2 OR2X2_2493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4313_));
OR2X2 OR2X2_2494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4314_));
OR2X2 OR2X2_2495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4316_));
OR2X2 OR2X2_2496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4317_));
OR2X2 OR2X2_2497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4319_));
OR2X2 OR2X2_2498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4320_));
OR2X2 OR2X2_2499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r12_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4322_));
OR2X2 OR2X2_25 ( .A(_abc_44694_new_n723_), .B(_abc_44694_new_n724_), .Y(_abc_44694_new_n725_));
OR2X2 OR2X2_250 ( .A(_abc_44694_new_n1382__bF_buf3), .B(_abc_44694_new_n1416_), .Y(_abc_44694_new_n1417_));
OR2X2 OR2X2_2500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4323_));
OR2X2 OR2X2_2501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r12_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4325_));
OR2X2 OR2X2_2502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4326_));
OR2X2 OR2X2_2503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r12_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4328_));
OR2X2 OR2X2_2504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4329_));
OR2X2 OR2X2_2505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r12_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4331_));
OR2X2 OR2X2_2506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4332_));
OR2X2 OR2X2_2507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4239__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r12_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4334_));
OR2X2 OR2X2_2508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4241__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4335_));
OR2X2 OR2X2_2509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4338_));
OR2X2 OR2X2_251 ( .A(_abc_44694_new_n1207__bF_buf5), .B(_abc_44694_new_n1412_), .Y(_abc_44694_new_n1418_));
OR2X2 OR2X2_2510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4340_));
OR2X2 OR2X2_2511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4342_));
OR2X2 OR2X2_2512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4343_));
OR2X2 OR2X2_2513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4345_));
OR2X2 OR2X2_2514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4346_));
OR2X2 OR2X2_2515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4348_));
OR2X2 OR2X2_2516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4349_));
OR2X2 OR2X2_2517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4351_));
OR2X2 OR2X2_2518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4352_));
OR2X2 OR2X2_2519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4354_));
OR2X2 OR2X2_252 ( .A(_abc_44694_new_n1419_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n1420_));
OR2X2 OR2X2_2520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4355_));
OR2X2 OR2X2_2521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4357_));
OR2X2 OR2X2_2522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4358_));
OR2X2 OR2X2_2523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4360_));
OR2X2 OR2X2_2524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4361_));
OR2X2 OR2X2_2525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4363_));
OR2X2 OR2X2_2526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4364_));
OR2X2 OR2X2_2527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4366_));
OR2X2 OR2X2_2528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4367_));
OR2X2 OR2X2_2529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4369_));
OR2X2 OR2X2_253 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(epc_q_2_), .Y(_abc_44694_new_n1421_));
OR2X2 OR2X2_2530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4370_));
OR2X2 OR2X2_2531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4372_));
OR2X2 OR2X2_2532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4373_));
OR2X2 OR2X2_2533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4375_));
OR2X2 OR2X2_2534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4376_));
OR2X2 OR2X2_2535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4378_));
OR2X2 OR2X2_2536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4379_));
OR2X2 OR2X2_2537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4381_));
OR2X2 OR2X2_2538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4382_));
OR2X2 OR2X2_2539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4384_));
OR2X2 OR2X2_254 ( .A(_abc_44694_new_n1348__bF_buf4), .B(epc_q_3_), .Y(_abc_44694_new_n1427_));
OR2X2 OR2X2_2540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4385_));
OR2X2 OR2X2_2541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4387_));
OR2X2 OR2X2_2542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4388_));
OR2X2 OR2X2_2543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4390_));
OR2X2 OR2X2_2544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4391_));
OR2X2 OR2X2_2545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4393_));
OR2X2 OR2X2_2546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4394_));
OR2X2 OR2X2_2547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4396_));
OR2X2 OR2X2_2548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4397_));
OR2X2 OR2X2_2549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4399_));
OR2X2 OR2X2_255 ( .A(_abc_44694_new_n1334__bF_buf1), .B(_abc_44694_new_n1428_), .Y(_abc_44694_new_n1429_));
OR2X2 OR2X2_2550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4400_));
OR2X2 OR2X2_2551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4402_));
OR2X2 OR2X2_2552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4403_));
OR2X2 OR2X2_2553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4405_));
OR2X2 OR2X2_2554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4406_));
OR2X2 OR2X2_2555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4408_));
OR2X2 OR2X2_2556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4409_));
OR2X2 OR2X2_2557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4411_));
OR2X2 OR2X2_2558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4412_));
OR2X2 OR2X2_2559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4414_));
OR2X2 OR2X2_256 ( .A(alu_op_r_1_), .B(pc_q_3_), .Y(_abc_44694_new_n1430_));
OR2X2 OR2X2_2560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4415_));
OR2X2 OR2X2_2561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4417_));
OR2X2 OR2X2_2562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4418_));
OR2X2 OR2X2_2563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r11_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4420_));
OR2X2 OR2X2_2564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4421_));
OR2X2 OR2X2_2565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r11_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4423_));
OR2X2 OR2X2_2566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4424_));
OR2X2 OR2X2_2567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r11_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4426_));
OR2X2 OR2X2_2568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4427_));
OR2X2 OR2X2_2569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r11_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4429_));
OR2X2 OR2X2_257 ( .A(_abc_44694_new_n1433_), .B(_abc_44694_new_n1403_), .Y(_abc_44694_new_n1434_));
OR2X2 OR2X2_2570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4430_));
OR2X2 OR2X2_2571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4337__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r11_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4432_));
OR2X2 OR2X2_2572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4339__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4433_));
OR2X2 OR2X2_2573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4436_));
OR2X2 OR2X2_2574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4440_));
OR2X2 OR2X2_2575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4444_));
OR2X2 OR2X2_2576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4448_));
OR2X2 OR2X2_2577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4452_));
OR2X2 OR2X2_2578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4456_));
OR2X2 OR2X2_2579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4460_));
OR2X2 OR2X2_258 ( .A(_abc_44694_new_n1337__bF_buf4), .B(_abc_44694_new_n1439_), .Y(_abc_44694_new_n1440_));
OR2X2 OR2X2_2580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4464_));
OR2X2 OR2X2_2581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4468_));
OR2X2 OR2X2_2582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4472_));
OR2X2 OR2X2_2583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4476_));
OR2X2 OR2X2_2584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4480_));
OR2X2 OR2X2_2585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4484_));
OR2X2 OR2X2_2586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4488_));
OR2X2 OR2X2_2587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4492_));
OR2X2 OR2X2_2588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4496_));
OR2X2 OR2X2_2589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4500_));
OR2X2 OR2X2_259 ( .A(_abc_44694_new_n1438_), .B(_abc_44694_new_n1440_), .Y(_abc_44694_new_n1441_));
OR2X2 OR2X2_2590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4504_));
OR2X2 OR2X2_2591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4508_));
OR2X2 OR2X2_2592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4512_));
OR2X2 OR2X2_2593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4516_));
OR2X2 OR2X2_2594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4520_));
OR2X2 OR2X2_2595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4524_));
OR2X2 OR2X2_2596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4528_));
OR2X2 OR2X2_2597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4532_));
OR2X2 OR2X2_2598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4536_));
OR2X2 OR2X2_2599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4540_));
OR2X2 OR2X2_26 ( .A(_abc_44694_new_n722_), .B(_abc_44694_new_n725_), .Y(_abc_44694_new_n726_));
OR2X2 OR2X2_260 ( .A(_abc_44694_new_n1340__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_3_), .Y(_abc_44694_new_n1442_));
OR2X2 OR2X2_2600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4544_));
OR2X2 OR2X2_2601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r10_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4548_));
OR2X2 OR2X2_2602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r10_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4552_));
OR2X2 OR2X2_2603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r10_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4556_));
OR2X2 OR2X2_2604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4435__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r10_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4560_));
OR2X2 OR2X2_2605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4565_));
OR2X2 OR2X2_2606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4567_));
OR2X2 OR2X2_2607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4569_));
OR2X2 OR2X2_2608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4570_));
OR2X2 OR2X2_2609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4572_));
OR2X2 OR2X2_261 ( .A(pc_q_2_), .B(pc_q_3_), .Y(_abc_44694_new_n1445_));
OR2X2 OR2X2_2610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4573_));
OR2X2 OR2X2_2611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4575_));
OR2X2 OR2X2_2612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4576_));
OR2X2 OR2X2_2613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4578_));
OR2X2 OR2X2_2614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4579_));
OR2X2 OR2X2_2615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4581_));
OR2X2 OR2X2_2616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4582_));
OR2X2 OR2X2_2617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4584_));
OR2X2 OR2X2_2618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4585_));
OR2X2 OR2X2_2619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4587_));
OR2X2 OR2X2_262 ( .A(_abc_44694_new_n1449_), .B(_abc_44694_new_n1444_), .Y(_abc_44694_new_n1450_));
OR2X2 OR2X2_2620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4588_));
OR2X2 OR2X2_2621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4590_));
OR2X2 OR2X2_2622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4591_));
OR2X2 OR2X2_2623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4593_));
OR2X2 OR2X2_2624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4594_));
OR2X2 OR2X2_2625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4596_));
OR2X2 OR2X2_2626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4597_));
OR2X2 OR2X2_2627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4599_));
OR2X2 OR2X2_2628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4600_));
OR2X2 OR2X2_2629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4602_));
OR2X2 OR2X2_263 ( .A(_abc_44694_new_n1450_), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n1451_));
OR2X2 OR2X2_2630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4603_));
OR2X2 OR2X2_2631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4605_));
OR2X2 OR2X2_2632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4606_));
OR2X2 OR2X2_2633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4608_));
OR2X2 OR2X2_2634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4609_));
OR2X2 OR2X2_2635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4611_));
OR2X2 OR2X2_2636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4612_));
OR2X2 OR2X2_2637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4614_));
OR2X2 OR2X2_2638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4615_));
OR2X2 OR2X2_2639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4617_));
OR2X2 OR2X2_264 ( .A(_abc_44694_new_n1382__bF_buf2), .B(_abc_44694_new_n1452_), .Y(_abc_44694_new_n1453_));
OR2X2 OR2X2_2640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4618_));
OR2X2 OR2X2_2641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4620_));
OR2X2 OR2X2_2642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4621_));
OR2X2 OR2X2_2643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4623_));
OR2X2 OR2X2_2644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4624_));
OR2X2 OR2X2_2645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4626_));
OR2X2 OR2X2_2646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4627_));
OR2X2 OR2X2_2647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4629_));
OR2X2 OR2X2_2648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4630_));
OR2X2 OR2X2_2649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4632_));
OR2X2 OR2X2_265 ( .A(_abc_44694_new_n1207__bF_buf4), .B(_abc_44694_new_n1448_), .Y(_abc_44694_new_n1454_));
OR2X2 OR2X2_2650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4633_));
OR2X2 OR2X2_2651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4635_));
OR2X2 OR2X2_2652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4636_));
OR2X2 OR2X2_2653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4638_));
OR2X2 OR2X2_2654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4639_));
OR2X2 OR2X2_2655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4641_));
OR2X2 OR2X2_2656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4642_));
OR2X2 OR2X2_2657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4644_));
OR2X2 OR2X2_2658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4645_));
OR2X2 OR2X2_2659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r1_sp_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4647_));
OR2X2 OR2X2_266 ( .A(_abc_44694_new_n1455_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n1456_));
OR2X2 OR2X2_2660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4648_));
OR2X2 OR2X2_2661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r1_sp_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4650_));
OR2X2 OR2X2_2662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4651_));
OR2X2 OR2X2_2663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r1_sp_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4653_));
OR2X2 OR2X2_2664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4654_));
OR2X2 OR2X2_2665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r1_sp_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4656_));
OR2X2 OR2X2_2666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4657_));
OR2X2 OR2X2_2667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4564__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r1_sp_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4659_));
OR2X2 OR2X2_2668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4566__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4660_));
OR2X2 OR2X2_2669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4663_));
OR2X2 OR2X2_267 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_3_), .Y(_abc_44694_new_n1457_));
OR2X2 OR2X2_2670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4667_));
OR2X2 OR2X2_2671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4671_));
OR2X2 OR2X2_2672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4675_));
OR2X2 OR2X2_2673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4679_));
OR2X2 OR2X2_2674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4683_));
OR2X2 OR2X2_2675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4687_));
OR2X2 OR2X2_2676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4691_));
OR2X2 OR2X2_2677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4695_));
OR2X2 OR2X2_2678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4699_));
OR2X2 OR2X2_2679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4703_));
OR2X2 OR2X2_268 ( .A(_abc_44694_new_n1348__bF_buf2), .B(epc_q_4_), .Y(_abc_44694_new_n1463_));
OR2X2 OR2X2_2680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4707_));
OR2X2 OR2X2_2681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4711_));
OR2X2 OR2X2_2682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4715_));
OR2X2 OR2X2_2683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4719_));
OR2X2 OR2X2_2684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4723_));
OR2X2 OR2X2_2685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4727_));
OR2X2 OR2X2_2686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4731_));
OR2X2 OR2X2_2687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4735_));
OR2X2 OR2X2_2688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4739_));
OR2X2 OR2X2_2689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4743_));
OR2X2 OR2X2_269 ( .A(_abc_44694_new_n1334__bF_buf0), .B(_abc_44694_new_n1464_), .Y(_abc_44694_new_n1465_));
OR2X2 OR2X2_2690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4747_));
OR2X2 OR2X2_2691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4751_));
OR2X2 OR2X2_2692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4755_));
OR2X2 OR2X2_2693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4759_));
OR2X2 OR2X2_2694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4763_));
OR2X2 OR2X2_2695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4767_));
OR2X2 OR2X2_2696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4771_));
OR2X2 OR2X2_2697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r9_lr_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4775_));
OR2X2 OR2X2_2698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r9_lr_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4779_));
OR2X2 OR2X2_2699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r9_lr_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4783_));
OR2X2 OR2X2_27 ( .A(_abc_44694_new_n673__bF_buf2), .B(_abc_44694_new_n726_), .Y(_abc_44694_new_n727_));
OR2X2 OR2X2_270 ( .A(alu_op_r_2_), .B(pc_q_4_), .Y(_abc_44694_new_n1467_));
OR2X2 OR2X2_2700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4662__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r9_lr_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4787_));
OR2X2 OR2X2_2701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4792_));
OR2X2 OR2X2_2702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4794_));
OR2X2 OR2X2_2703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4796_));
OR2X2 OR2X2_2704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4797_));
OR2X2 OR2X2_2705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4799_));
OR2X2 OR2X2_2706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4800_));
OR2X2 OR2X2_2707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4802_));
OR2X2 OR2X2_2708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4803_));
OR2X2 OR2X2_2709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4805_));
OR2X2 OR2X2_271 ( .A(_abc_44694_new_n1466_), .B(_abc_44694_new_n1471_), .Y(_abc_44694_new_n1472_));
OR2X2 OR2X2_2710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4806_));
OR2X2 OR2X2_2711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4808_));
OR2X2 OR2X2_2712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4809_));
OR2X2 OR2X2_2713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4811_));
OR2X2 OR2X2_2714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4812_));
OR2X2 OR2X2_2715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4814_));
OR2X2 OR2X2_2716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4815_));
OR2X2 OR2X2_2717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4817_));
OR2X2 OR2X2_2718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4818_));
OR2X2 OR2X2_2719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4820_));
OR2X2 OR2X2_272 ( .A(_abc_44694_new_n1473_), .B(_abc_44694_new_n1470_), .Y(_abc_44694_new_n1474_));
OR2X2 OR2X2_2720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4821_));
OR2X2 OR2X2_2721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4823_));
OR2X2 OR2X2_2722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4824_));
OR2X2 OR2X2_2723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4826_));
OR2X2 OR2X2_2724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4827_));
OR2X2 OR2X2_2725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4829_));
OR2X2 OR2X2_2726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4830_));
OR2X2 OR2X2_2727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4832_));
OR2X2 OR2X2_2728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4833_));
OR2X2 OR2X2_2729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4835_));
OR2X2 OR2X2_273 ( .A(_abc_44694_new_n1337__bF_buf3), .B(_abc_44694_new_n1477_), .Y(_abc_44694_new_n1478_));
OR2X2 OR2X2_2730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4836_));
OR2X2 OR2X2_2731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4838_));
OR2X2 OR2X2_2732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4839_));
OR2X2 OR2X2_2733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4841_));
OR2X2 OR2X2_2734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4842_));
OR2X2 OR2X2_2735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4844_));
OR2X2 OR2X2_2736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4845_));
OR2X2 OR2X2_2737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4847_));
OR2X2 OR2X2_2738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4848_));
OR2X2 OR2X2_2739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4850_));
OR2X2 OR2X2_274 ( .A(_abc_44694_new_n1476_), .B(_abc_44694_new_n1478_), .Y(_abc_44694_new_n1479_));
OR2X2 OR2X2_2740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4851_));
OR2X2 OR2X2_2741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4853_));
OR2X2 OR2X2_2742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4854_));
OR2X2 OR2X2_2743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4856_));
OR2X2 OR2X2_2744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4857_));
OR2X2 OR2X2_2745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4859_));
OR2X2 OR2X2_2746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4860_));
OR2X2 OR2X2_2747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4862_));
OR2X2 OR2X2_2748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4863_));
OR2X2 OR2X2_2749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4865_));
OR2X2 OR2X2_275 ( .A(_abc_44694_new_n1340__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_4_), .Y(_abc_44694_new_n1480_));
OR2X2 OR2X2_2750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4866_));
OR2X2 OR2X2_2751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4868_));
OR2X2 OR2X2_2752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4869_));
OR2X2 OR2X2_2753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4871_));
OR2X2 OR2X2_2754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4872_));
OR2X2 OR2X2_2755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r8_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4874_));
OR2X2 OR2X2_2756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4875_));
OR2X2 OR2X2_2757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r8_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4877_));
OR2X2 OR2X2_2758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4878_));
OR2X2 OR2X2_2759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r8_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4880_));
OR2X2 OR2X2_276 ( .A(_abc_44694_new_n1446_), .B(pc_q_4_), .Y(_abc_44694_new_n1483_));
OR2X2 OR2X2_2760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4881_));
OR2X2 OR2X2_2761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r8_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4883_));
OR2X2 OR2X2_2762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4884_));
OR2X2 OR2X2_2763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4791__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r8_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4886_));
OR2X2 OR2X2_2764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4793__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4887_));
OR2X2 OR2X2_2765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4890_));
OR2X2 OR2X2_2766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4892_));
OR2X2 OR2X2_2767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4894_));
OR2X2 OR2X2_2768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4895_));
OR2X2 OR2X2_2769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4897_));
OR2X2 OR2X2_277 ( .A(_abc_44694_new_n1487_), .B(_abc_44694_new_n1482_), .Y(_abc_44694_new_n1488_));
OR2X2 OR2X2_2770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4898_));
OR2X2 OR2X2_2771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4900_));
OR2X2 OR2X2_2772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4901_));
OR2X2 OR2X2_2773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4903_));
OR2X2 OR2X2_2774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4904_));
OR2X2 OR2X2_2775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4906_));
OR2X2 OR2X2_2776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4907_));
OR2X2 OR2X2_2777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4909_));
OR2X2 OR2X2_2778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4910_));
OR2X2 OR2X2_2779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4912_));
OR2X2 OR2X2_278 ( .A(_abc_44694_new_n1488_), .B(_abc_44694_new_n1278__bF_buf4), .Y(_abc_44694_new_n1489_));
OR2X2 OR2X2_2780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4913_));
OR2X2 OR2X2_2781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4915_));
OR2X2 OR2X2_2782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4916_));
OR2X2 OR2X2_2783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4918_));
OR2X2 OR2X2_2784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4919_));
OR2X2 OR2X2_2785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4921_));
OR2X2 OR2X2_2786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4922_));
OR2X2 OR2X2_2787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4924_));
OR2X2 OR2X2_2788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4925_));
OR2X2 OR2X2_2789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4927_));
OR2X2 OR2X2_279 ( .A(_abc_44694_new_n1382__bF_buf1), .B(_abc_44694_new_n1490_), .Y(_abc_44694_new_n1491_));
OR2X2 OR2X2_2790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4928_));
OR2X2 OR2X2_2791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4930_));
OR2X2 OR2X2_2792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4931_));
OR2X2 OR2X2_2793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4933_));
OR2X2 OR2X2_2794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4934_));
OR2X2 OR2X2_2795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4936_));
OR2X2 OR2X2_2796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4937_));
OR2X2 OR2X2_2797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4939_));
OR2X2 OR2X2_2798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4940_));
OR2X2 OR2X2_2799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4942_));
OR2X2 OR2X2_28 ( .A(_abc_44694_new_n729_), .B(_abc_44694_new_n715_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_2_));
OR2X2 OR2X2_280 ( .A(_abc_44694_new_n1207__bF_buf3), .B(_abc_44694_new_n1486_), .Y(_abc_44694_new_n1492_));
OR2X2 OR2X2_2800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4943_));
OR2X2 OR2X2_2801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4945_));
OR2X2 OR2X2_2802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4946_));
OR2X2 OR2X2_2803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4948_));
OR2X2 OR2X2_2804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4949_));
OR2X2 OR2X2_2805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4951_));
OR2X2 OR2X2_2806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4952_));
OR2X2 OR2X2_2807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4954_));
OR2X2 OR2X2_2808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4955_));
OR2X2 OR2X2_2809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4957_));
OR2X2 OR2X2_281 ( .A(_abc_44694_new_n1493_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n1494_));
OR2X2 OR2X2_2810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4958_));
OR2X2 OR2X2_2811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4960_));
OR2X2 OR2X2_2812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4961_));
OR2X2 OR2X2_2813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4963_));
OR2X2 OR2X2_2814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4964_));
OR2X2 OR2X2_2815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4966_));
OR2X2 OR2X2_2816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4967_));
OR2X2 OR2X2_2817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4969_));
OR2X2 OR2X2_2818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4970_));
OR2X2 OR2X2_2819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r7_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4972_));
OR2X2 OR2X2_282 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_4_), .Y(_abc_44694_new_n1495_));
OR2X2 OR2X2_2820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4973_));
OR2X2 OR2X2_2821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r7_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4975_));
OR2X2 OR2X2_2822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4976_));
OR2X2 OR2X2_2823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r7_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4978_));
OR2X2 OR2X2_2824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4979_));
OR2X2 OR2X2_2825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r7_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4981_));
OR2X2 OR2X2_2826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4982_));
OR2X2 OR2X2_2827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4889__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r7_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4984_));
OR2X2 OR2X2_2828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4891__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4985_));
OR2X2 OR2X2_2829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4988_));
OR2X2 OR2X2_283 ( .A(_abc_44694_new_n1484_), .B(pc_q_5_), .Y(_abc_44694_new_n1498_));
OR2X2 OR2X2_2830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4992_));
OR2X2 OR2X2_2831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n4996_));
OR2X2 OR2X2_2832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5000_));
OR2X2 OR2X2_2833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5004_));
OR2X2 OR2X2_2834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5008_));
OR2X2 OR2X2_2835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5012_));
OR2X2 OR2X2_2836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5016_));
OR2X2 OR2X2_2837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5020_));
OR2X2 OR2X2_2838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5024_));
OR2X2 OR2X2_2839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5028_));
OR2X2 OR2X2_284 ( .A(_abc_44694_new_n1399__bF_buf0), .B(_abc_44694_new_n1501_), .Y(_abc_44694_new_n1502_));
OR2X2 OR2X2_2840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5032_));
OR2X2 OR2X2_2841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5036_));
OR2X2 OR2X2_2842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5040_));
OR2X2 OR2X2_2843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5044_));
OR2X2 OR2X2_2844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5048_));
OR2X2 OR2X2_2845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5052_));
OR2X2 OR2X2_2846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5056_));
OR2X2 OR2X2_2847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5060_));
OR2X2 OR2X2_2848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5064_));
OR2X2 OR2X2_2849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5068_));
OR2X2 OR2X2_285 ( .A(alu_op_r_3_), .B(pc_q_5_), .Y(_abc_44694_new_n1504_));
OR2X2 OR2X2_2850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5072_));
OR2X2 OR2X2_2851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5076_));
OR2X2 OR2X2_2852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5080_));
OR2X2 OR2X2_2853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5084_));
OR2X2 OR2X2_2854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5088_));
OR2X2 OR2X2_2855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5092_));
OR2X2 OR2X2_2856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5096_));
OR2X2 OR2X2_2857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r6_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5100_));
OR2X2 OR2X2_2858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r6_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5104_));
OR2X2 OR2X2_2859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r6_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5108_));
OR2X2 OR2X2_286 ( .A(_abc_44694_new_n1511_), .B(_abc_44694_new_n1512_), .Y(_abc_44694_new_n1513_));
OR2X2 OR2X2_2860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n4987__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r6_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5112_));
OR2X2 OR2X2_2861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5117_));
OR2X2 OR2X2_2862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5121_));
OR2X2 OR2X2_2863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5125_));
OR2X2 OR2X2_2864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5129_));
OR2X2 OR2X2_2865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5133_));
OR2X2 OR2X2_2866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5137_));
OR2X2 OR2X2_2867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5141_));
OR2X2 OR2X2_2868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5145_));
OR2X2 OR2X2_2869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5149_));
OR2X2 OR2X2_287 ( .A(_abc_44694_new_n1514_), .B(_abc_44694_new_n1503_), .Y(_abc_44694_new_n1515_));
OR2X2 OR2X2_2870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5153_));
OR2X2 OR2X2_2871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5157_));
OR2X2 OR2X2_2872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5161_));
OR2X2 OR2X2_2873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5165_));
OR2X2 OR2X2_2874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5169_));
OR2X2 OR2X2_2875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5173_));
OR2X2 OR2X2_2876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5177_));
OR2X2 OR2X2_2877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5181_));
OR2X2 OR2X2_2878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5185_));
OR2X2 OR2X2_2879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5189_));
OR2X2 OR2X2_288 ( .A(_abc_44694_new_n1400__bF_buf1), .B(_abc_44694_new_n1517_), .Y(_abc_44694_new_n1518_));
OR2X2 OR2X2_2880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5193_));
OR2X2 OR2X2_2881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5197_));
OR2X2 OR2X2_2882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5201_));
OR2X2 OR2X2_2883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5205_));
OR2X2 OR2X2_2884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5209_));
OR2X2 OR2X2_2885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5213_));
OR2X2 OR2X2_2886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5217_));
OR2X2 OR2X2_2887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5221_));
OR2X2 OR2X2_2888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5225_));
OR2X2 OR2X2_2889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf7), .B(REGFILE_SIM_reg_bank_reg_r5_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5229_));
OR2X2 OR2X2_289 ( .A(_abc_44694_new_n1516_), .B(_abc_44694_new_n1518_), .Y(_abc_44694_new_n1519_));
OR2X2 OR2X2_2890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf5), .B(REGFILE_SIM_reg_bank_reg_r5_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5233_));
OR2X2 OR2X2_2891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r5_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5237_));
OR2X2 OR2X2_2892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5116__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r5_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5241_));
OR2X2 OR2X2_2893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5246_));
OR2X2 OR2X2_2894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5248_));
OR2X2 OR2X2_2895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5250_));
OR2X2 OR2X2_2896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5251_));
OR2X2 OR2X2_2897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5253_));
OR2X2 OR2X2_2898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5254_));
OR2X2 OR2X2_2899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5256_));
OR2X2 OR2X2_29 ( .A(_abc_44694_new_n733_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n734_));
OR2X2 OR2X2_290 ( .A(_abc_44694_new_n1520_), .B(_abc_44694_new_n1278__bF_buf3), .Y(_abc_44694_new_n1521_));
OR2X2 OR2X2_2900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5257_));
OR2X2 OR2X2_2901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5259_));
OR2X2 OR2X2_2902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5260_));
OR2X2 OR2X2_2903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5262_));
OR2X2 OR2X2_2904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5263_));
OR2X2 OR2X2_2905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5265_));
OR2X2 OR2X2_2906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5266_));
OR2X2 OR2X2_2907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5268_));
OR2X2 OR2X2_2908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5269_));
OR2X2 OR2X2_2909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5271_));
OR2X2 OR2X2_291 ( .A(_abc_44694_new_n1523_), .B(_abc_44694_new_n1524_), .Y(_abc_44694_new_n1525_));
OR2X2 OR2X2_2910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5272_));
OR2X2 OR2X2_2911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5274_));
OR2X2 OR2X2_2912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5275_));
OR2X2 OR2X2_2913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5277_));
OR2X2 OR2X2_2914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5278_));
OR2X2 OR2X2_2915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5280_));
OR2X2 OR2X2_2916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5281_));
OR2X2 OR2X2_2917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5283_));
OR2X2 OR2X2_2918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5284_));
OR2X2 OR2X2_2919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5286_));
OR2X2 OR2X2_292 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n1525_), .Y(_abc_44694_new_n1526_));
OR2X2 OR2X2_2920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5287_));
OR2X2 OR2X2_2921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5289_));
OR2X2 OR2X2_2922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5290_));
OR2X2 OR2X2_2923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5292_));
OR2X2 OR2X2_2924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5293_));
OR2X2 OR2X2_2925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5295_));
OR2X2 OR2X2_2926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5296_));
OR2X2 OR2X2_2927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5298_));
OR2X2 OR2X2_2928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5299_));
OR2X2 OR2X2_2929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5301_));
OR2X2 OR2X2_293 ( .A(_abc_44694_new_n1527_), .B(_abc_44694_new_n1382__bF_buf0), .Y(_abc_44694_new_n1528_));
OR2X2 OR2X2_2930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5302_));
OR2X2 OR2X2_2931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5304_));
OR2X2 OR2X2_2932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5305_));
OR2X2 OR2X2_2933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5307_));
OR2X2 OR2X2_2934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5308_));
OR2X2 OR2X2_2935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5310_));
OR2X2 OR2X2_2936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5311_));
OR2X2 OR2X2_2937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5313_));
OR2X2 OR2X2_2938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5314_));
OR2X2 OR2X2_2939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5316_));
OR2X2 OR2X2_294 ( .A(_abc_44694_new_n1207__bF_buf2), .B(_abc_44694_new_n1501_), .Y(_abc_44694_new_n1529_));
OR2X2 OR2X2_2940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5317_));
OR2X2 OR2X2_2941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5319_));
OR2X2 OR2X2_2942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5320_));
OR2X2 OR2X2_2943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5322_));
OR2X2 OR2X2_2944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5323_));
OR2X2 OR2X2_2945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5325_));
OR2X2 OR2X2_2946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5326_));
OR2X2 OR2X2_2947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r4_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5328_));
OR2X2 OR2X2_2948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5329_));
OR2X2 OR2X2_2949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r4_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5331_));
OR2X2 OR2X2_295 ( .A(_abc_44694_new_n1530_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n1531_));
OR2X2 OR2X2_2950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5332_));
OR2X2 OR2X2_2951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r4_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5334_));
OR2X2 OR2X2_2952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5335_));
OR2X2 OR2X2_2953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r4_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5337_));
OR2X2 OR2X2_2954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5338_));
OR2X2 OR2X2_2955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5245__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r4_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5340_));
OR2X2 OR2X2_2956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5247__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5341_));
OR2X2 OR2X2_2957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5344_));
OR2X2 OR2X2_2958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5346_));
OR2X2 OR2X2_2959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5348_));
OR2X2 OR2X2_296 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_5_), .Y(_abc_44694_new_n1532_));
OR2X2 OR2X2_2960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5349_));
OR2X2 OR2X2_2961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5351_));
OR2X2 OR2X2_2962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5352_));
OR2X2 OR2X2_2963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5354_));
OR2X2 OR2X2_2964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5355_));
OR2X2 OR2X2_2965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5357_));
OR2X2 OR2X2_2966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5358_));
OR2X2 OR2X2_2967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5360_));
OR2X2 OR2X2_2968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5361_));
OR2X2 OR2X2_2969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5363_));
OR2X2 OR2X2_297 ( .A(_abc_44694_new_n1499_), .B(pc_q_6_), .Y(_abc_44694_new_n1536_));
OR2X2 OR2X2_2970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5364_));
OR2X2 OR2X2_2971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5366_));
OR2X2 OR2X2_2972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5367_));
OR2X2 OR2X2_2973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5369_));
OR2X2 OR2X2_2974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5370_));
OR2X2 OR2X2_2975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5372_));
OR2X2 OR2X2_2976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5373_));
OR2X2 OR2X2_2977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5375_));
OR2X2 OR2X2_2978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5376_));
OR2X2 OR2X2_2979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5378_));
OR2X2 OR2X2_298 ( .A(_abc_44694_new_n1539_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n1540_));
OR2X2 OR2X2_2980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5379_));
OR2X2 OR2X2_2981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5381_));
OR2X2 OR2X2_2982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5382_));
OR2X2 OR2X2_2983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5384_));
OR2X2 OR2X2_2984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5385_));
OR2X2 OR2X2_2985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5387_));
OR2X2 OR2X2_2986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5388_));
OR2X2 OR2X2_2987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5390_));
OR2X2 OR2X2_2988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5391_));
OR2X2 OR2X2_2989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5393_));
OR2X2 OR2X2_299 ( .A(_abc_44694_new_n1399__bF_buf4), .B(_abc_44694_new_n1539_), .Y(_abc_44694_new_n1542_));
OR2X2 OR2X2_2990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5394_));
OR2X2 OR2X2_2991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5396_));
OR2X2 OR2X2_2992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5397_));
OR2X2 OR2X2_2993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5399_));
OR2X2 OR2X2_2994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5400_));
OR2X2 OR2X2_2995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5402_));
OR2X2 OR2X2_2996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5403_));
OR2X2 OR2X2_2997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5405_));
OR2X2 OR2X2_2998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5406_));
OR2X2 OR2X2_2999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5408_));
OR2X2 OR2X2_3 ( .A(_abc_44694_new_n656_), .B(_abc_44694_new_n658_), .Y(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_4_));
OR2X2 OR2X2_30 ( .A(_abc_44694_new_n734_), .B(_abc_44694_new_n732_), .Y(_abc_44694_new_n735_));
OR2X2 OR2X2_300 ( .A(_abc_44694_new_n1546_), .B(_abc_44694_new_n1505_), .Y(_abc_44694_new_n1547_));
OR2X2 OR2X2_3000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5409_));
OR2X2 OR2X2_3001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5411_));
OR2X2 OR2X2_3002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5412_));
OR2X2 OR2X2_3003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5414_));
OR2X2 OR2X2_3004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5415_));
OR2X2 OR2X2_3005 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5417_));
OR2X2 OR2X2_3006 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5418_));
OR2X2 OR2X2_3007 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5420_));
OR2X2 OR2X2_3008 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5421_));
OR2X2 OR2X2_3009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5423_));
OR2X2 OR2X2_301 ( .A(_abc_44694_new_n1545_), .B(_abc_44694_new_n1547_), .Y(_abc_44694_new_n1548_));
OR2X2 OR2X2_3010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5424_));
OR2X2 OR2X2_3011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r3_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5426_));
OR2X2 OR2X2_3012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5427_));
OR2X2 OR2X2_3013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r3_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5429_));
OR2X2 OR2X2_3014 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5430_));
OR2X2 OR2X2_3015 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r3_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5432_));
OR2X2 OR2X2_3016 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5433_));
OR2X2 OR2X2_3017 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r3_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5435_));
OR2X2 OR2X2_3018 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5436_));
OR2X2 OR2X2_3019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5343__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r3_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5438_));
OR2X2 OR2X2_302 ( .A(int32_r_4_), .B(pc_q_6_), .Y(_abc_44694_new_n1549_));
OR2X2 OR2X2_3020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5345__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5439_));
OR2X2 OR2X2_3021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_0_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5442_));
OR2X2 OR2X2_3022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_0_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5444_));
OR2X2 OR2X2_3023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_1_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5446_));
OR2X2 OR2X2_3024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_1_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5447_));
OR2X2 OR2X2_3025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_2_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5449_));
OR2X2 OR2X2_3026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_2_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5450_));
OR2X2 OR2X2_3027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5452_));
OR2X2 OR2X2_3028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_3_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5453_));
OR2X2 OR2X2_3029 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_4_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5455_));
OR2X2 OR2X2_303 ( .A(_abc_44694_new_n1548_), .B(_abc_44694_new_n1552_), .Y(_abc_44694_new_n1553_));
OR2X2 OR2X2_3030 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_4_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5456_));
OR2X2 OR2X2_3031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_5_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5458_));
OR2X2 OR2X2_3032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_5_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5459_));
OR2X2 OR2X2_3033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_6_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5461_));
OR2X2 OR2X2_3034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_6_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5462_));
OR2X2 OR2X2_3035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_7_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5464_));
OR2X2 OR2X2_3036 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_7_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5465_));
OR2X2 OR2X2_3037 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_8_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5467_));
OR2X2 OR2X2_3038 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_8_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5468_));
OR2X2 OR2X2_3039 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_9_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5470_));
OR2X2 OR2X2_304 ( .A(_abc_44694_new_n1557_), .B(_abc_44694_new_n1543_), .Y(_abc_44694_new_n1558_));
OR2X2 OR2X2_3040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_9_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5471_));
OR2X2 OR2X2_3041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_10_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5473_));
OR2X2 OR2X2_3042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_10_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5474_));
OR2X2 OR2X2_3043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_11_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5476_));
OR2X2 OR2X2_3044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_11_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5477_));
OR2X2 OR2X2_3045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_12_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5479_));
OR2X2 OR2X2_3046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_12_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5480_));
OR2X2 OR2X2_3047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_13_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5482_));
OR2X2 OR2X2_3048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_13_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5483_));
OR2X2 OR2X2_3049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_14_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5485_));
OR2X2 OR2X2_305 ( .A(_abc_44694_new_n1400__bF_buf0), .B(_abc_44694_new_n1560_), .Y(_abc_44694_new_n1561_));
OR2X2 OR2X2_3050 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_14_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5486_));
OR2X2 OR2X2_3051 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_15_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5488_));
OR2X2 OR2X2_3052 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_15_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5489_));
OR2X2 OR2X2_3053 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_16_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5491_));
OR2X2 OR2X2_3054 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_16_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5492_));
OR2X2 OR2X2_3055 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_17_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5494_));
OR2X2 OR2X2_3056 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_17_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5495_));
OR2X2 OR2X2_3057 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_18_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5497_));
OR2X2 OR2X2_3058 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_18_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5498_));
OR2X2 OR2X2_3059 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_19_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5500_));
OR2X2 OR2X2_306 ( .A(_abc_44694_new_n1559_), .B(_abc_44694_new_n1561_), .Y(_abc_44694_new_n1562_));
OR2X2 OR2X2_3060 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_19_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5501_));
OR2X2 OR2X2_3061 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_20_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5503_));
OR2X2 OR2X2_3062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_20_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5504_));
OR2X2 OR2X2_3063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_21_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5506_));
OR2X2 OR2X2_3064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_21_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5507_));
OR2X2 OR2X2_3065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_22_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5509_));
OR2X2 OR2X2_3066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_22_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5510_));
OR2X2 OR2X2_3067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_23_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5512_));
OR2X2 OR2X2_3068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_23_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5513_));
OR2X2 OR2X2_3069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_24_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5515_));
OR2X2 OR2X2_307 ( .A(_abc_44694_new_n1563_), .B(_abc_44694_new_n1278__bF_buf2), .Y(_abc_44694_new_n1564_));
OR2X2 OR2X2_3070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_24_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5516_));
OR2X2 OR2X2_3071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_25_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5518_));
OR2X2 OR2X2_3072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_25_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5519_));
OR2X2 OR2X2_3073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_26_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5521_));
OR2X2 OR2X2_3074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_26_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5522_));
OR2X2 OR2X2_3075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_r2_fp_27_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5524_));
OR2X2 OR2X2_3076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rd_i_27_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5525_));
OR2X2 OR2X2_3077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_r2_fp_28_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5527_));
OR2X2 OR2X2_3078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rd_i_28_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5528_));
OR2X2 OR2X2_3079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_r2_fp_29_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5530_));
OR2X2 OR2X2_308 ( .A(_abc_44694_new_n1565_), .B(_abc_44694_new_n1566_), .Y(_abc_44694_new_n1567_));
OR2X2 OR2X2_3080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rd_i_29_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5531_));
OR2X2 OR2X2_3081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_r2_fp_30_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5533_));
OR2X2 OR2X2_3082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf4), .B(REGFILE_SIM_reg_bank_reg_rd_i_30_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5534_));
OR2X2 OR2X2_3083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5441__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_r2_fp_31_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5536_));
OR2X2 OR2X2_3084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5443__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rd_i_31_bF_buf3_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5537_));
OR2X2 OR2X2_3085 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5549_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5544_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5550_));
OR2X2 OR2X2_3086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5555_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5559_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5560_));
OR2X2 OR2X2_3087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5560_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5550_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5561_));
OR2X2 OR2X2_3088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5566_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5569_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5570_));
OR2X2 OR2X2_3089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5573_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5576_));
OR2X2 OR2X2_309 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n1567_), .Y(_abc_44694_new_n1568_));
OR2X2 OR2X2_3090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5576_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5570_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5577_));
OR2X2 OR2X2_3091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5577_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5561_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5578_));
OR2X2 OR2X2_3092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5586_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5589_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5590_));
OR2X2 OR2X2_3093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5590_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5583_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5591_));
OR2X2 OR2X2_3094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5595_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5597_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5598_));
OR2X2 OR2X2_3095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5604_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5601_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5605_));
OR2X2 OR2X2_3096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5598_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5605_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5606_));
OR2X2 OR2X2_3097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5606_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5591_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5607_));
OR2X2 OR2X2_3098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5607_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5608_));
OR2X2 OR2X2_3099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5612_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5613_));
OR2X2 OR2X2_31 ( .A(_abc_44694_new_n736_), .B(_abc_44694_new_n737_), .Y(_abc_44694_new_n738_));
OR2X2 OR2X2_310 ( .A(_abc_44694_new_n1541_), .B(_abc_44694_new_n1570_), .Y(_abc_44694_new_n1571_));
OR2X2 OR2X2_3100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5616_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5619_));
OR2X2 OR2X2_3101 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5619_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5620_));
OR2X2 OR2X2_3102 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5622_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5624_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5625_));
OR2X2 OR2X2_3103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5627_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5629_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5630_));
OR2X2 OR2X2_3104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5625_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5630_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5631_));
OR2X2 OR2X2_3105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5631_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5620_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5632_));
OR2X2 OR2X2_3106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5634_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5637_));
OR2X2 OR2X2_3107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5639_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5641_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5642_));
OR2X2 OR2X2_3108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5637_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5642_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5643_));
OR2X2 OR2X2_3109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5645_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5647_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5648_));
OR2X2 OR2X2_311 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_6_), .Y(_abc_44694_new_n1572_));
OR2X2 OR2X2_3110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5650_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5652_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5653_));
OR2X2 OR2X2_3111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5648_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5653_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5654_));
OR2X2 OR2X2_3112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5643_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5654_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5655_));
OR2X2 OR2X2_3113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5655_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5632_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5656_));
OR2X2 OR2X2_3114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5608_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5656_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_0_));
OR2X2 OR2X2_3115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5659_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5658_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5660_));
OR2X2 OR2X2_3116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5661_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5663_));
OR2X2 OR2X2_3117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5663_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5660_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5664_));
OR2X2 OR2X2_3118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5665_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5666_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5667_));
OR2X2 OR2X2_3119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5668_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5669_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5670_));
OR2X2 OR2X2_312 ( .A(_abc_44694_new_n1537_), .B(pc_q_7_), .Y(_abc_44694_new_n1575_));
OR2X2 OR2X2_3120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5670_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5667_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5671_));
OR2X2 OR2X2_3121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5671_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5664_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5672_));
OR2X2 OR2X2_3122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5674_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5675_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5676_));
OR2X2 OR2X2_3123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5676_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5673_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5677_));
OR2X2 OR2X2_3124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5678_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5679_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5680_));
OR2X2 OR2X2_3125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5682_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5681_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5683_));
OR2X2 OR2X2_3126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5680_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5683_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5684_));
OR2X2 OR2X2_3127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5684_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5677_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5685_));
OR2X2 OR2X2_3128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5685_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5672_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5686_));
OR2X2 OR2X2_3129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5688_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5687_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5689_));
OR2X2 OR2X2_313 ( .A(_abc_44694_new_n1578_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n1579_));
OR2X2 OR2X2_3130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5690_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5691_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5692_));
OR2X2 OR2X2_3131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5692_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5689_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5693_));
OR2X2 OR2X2_3132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5694_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5695_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5696_));
OR2X2 OR2X2_3133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5697_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5698_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5699_));
OR2X2 OR2X2_3134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5696_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5700_));
OR2X2 OR2X2_3135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5700_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5693_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5701_));
OR2X2 OR2X2_3136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5702_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5703_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5704_));
OR2X2 OR2X2_3137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5705_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5706_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5707_));
OR2X2 OR2X2_3138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5704_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5707_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5708_));
OR2X2 OR2X2_3139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5709_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5710_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5711_));
OR2X2 OR2X2_314 ( .A(_abc_44694_new_n1399__bF_buf3), .B(_abc_44694_new_n1578_), .Y(_abc_44694_new_n1581_));
OR2X2 OR2X2_3140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5712_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5713_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5714_));
OR2X2 OR2X2_3141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5711_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5714_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5715_));
OR2X2 OR2X2_3142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5708_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5715_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5716_));
OR2X2 OR2X2_3143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5716_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5701_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5717_));
OR2X2 OR2X2_3144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5686_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5717_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_1_));
OR2X2 OR2X2_3145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5720_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5719_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5721_));
OR2X2 OR2X2_3146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5722_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5723_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5724_));
OR2X2 OR2X2_3147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5724_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5721_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5725_));
OR2X2 OR2X2_3148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5726_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5727_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5728_));
OR2X2 OR2X2_3149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5729_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5730_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5731_));
OR2X2 OR2X2_315 ( .A(int32_r_5_), .B(pc_q_7_), .Y(_abc_44694_new_n1583_));
OR2X2 OR2X2_3150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5731_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5728_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5732_));
OR2X2 OR2X2_3151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5732_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5725_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5733_));
OR2X2 OR2X2_3152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5735_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5736_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5737_));
OR2X2 OR2X2_3153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5737_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5734_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5738_));
OR2X2 OR2X2_3154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5739_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5740_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5741_));
OR2X2 OR2X2_3155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5743_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5742_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5744_));
OR2X2 OR2X2_3156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5741_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5744_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5745_));
OR2X2 OR2X2_3157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5745_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5738_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5746_));
OR2X2 OR2X2_3158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5746_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5733_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5747_));
OR2X2 OR2X2_3159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5749_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5748_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5750_));
OR2X2 OR2X2_316 ( .A(_abc_44694_new_n1586_), .B(_abc_44694_new_n1550_), .Y(_abc_44694_new_n1587_));
OR2X2 OR2X2_3160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5751_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5752_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5753_));
OR2X2 OR2X2_3161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5753_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5750_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5754_));
OR2X2 OR2X2_3162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5755_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5756_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5757_));
OR2X2 OR2X2_3163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5758_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5759_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5760_));
OR2X2 OR2X2_3164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5757_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5760_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5761_));
OR2X2 OR2X2_3165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5761_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5754_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5762_));
OR2X2 OR2X2_3166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5763_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5764_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5765_));
OR2X2 OR2X2_3167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5766_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5767_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5768_));
OR2X2 OR2X2_3168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5765_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5768_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5769_));
OR2X2 OR2X2_3169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5770_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5771_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5772_));
OR2X2 OR2X2_317 ( .A(_abc_44694_new_n1554_), .B(_abc_44694_new_n1587_), .Y(_abc_44694_new_n1588_));
OR2X2 OR2X2_3170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5773_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5774_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5775_));
OR2X2 OR2X2_3171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5772_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5775_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5776_));
OR2X2 OR2X2_3172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5769_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5776_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5777_));
OR2X2 OR2X2_3173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5777_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5762_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5778_));
OR2X2 OR2X2_3174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5747_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5778_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_2_));
OR2X2 OR2X2_3175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5781_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5780_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5782_));
OR2X2 OR2X2_3176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5783_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5784_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5785_));
OR2X2 OR2X2_3177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5785_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5782_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5786_));
OR2X2 OR2X2_3178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5787_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5788_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5789_));
OR2X2 OR2X2_3179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5790_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5792_));
OR2X2 OR2X2_318 ( .A(_abc_44694_new_n1596_), .B(_abc_44694_new_n1582_), .Y(_abc_44694_new_n1597_));
OR2X2 OR2X2_3180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5792_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5789_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5793_));
OR2X2 OR2X2_3181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5793_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5786_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5794_));
OR2X2 OR2X2_3182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5796_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5797_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5798_));
OR2X2 OR2X2_3183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5798_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5795_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5799_));
OR2X2 OR2X2_3184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5800_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5801_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5802_));
OR2X2 OR2X2_3185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5804_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5803_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5805_));
OR2X2 OR2X2_3186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5802_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5805_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5806_));
OR2X2 OR2X2_3187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5806_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5799_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5807_));
OR2X2 OR2X2_3188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5807_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5794_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5808_));
OR2X2 OR2X2_3189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5810_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5809_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5811_));
OR2X2 OR2X2_319 ( .A(_abc_44694_new_n1400__bF_buf4), .B(_abc_44694_new_n1599_), .Y(_abc_44694_new_n1600_));
OR2X2 OR2X2_3190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5812_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5814_));
OR2X2 OR2X2_3191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5814_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5811_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5815_));
OR2X2 OR2X2_3192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5816_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5817_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5818_));
OR2X2 OR2X2_3193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5819_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5820_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5821_));
OR2X2 OR2X2_3194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5818_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5821_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5822_));
OR2X2 OR2X2_3195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5822_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5823_));
OR2X2 OR2X2_3196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5824_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5825_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5826_));
OR2X2 OR2X2_3197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5827_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5828_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5829_));
OR2X2 OR2X2_3198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5826_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5830_));
OR2X2 OR2X2_3199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5831_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5832_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5833_));
OR2X2 OR2X2_32 ( .A(_abc_44694_new_n739_), .B(_abc_44694_new_n740_), .Y(_abc_44694_new_n741_));
OR2X2 OR2X2_320 ( .A(_abc_44694_new_n1598_), .B(_abc_44694_new_n1600_), .Y(_abc_44694_new_n1601_));
OR2X2 OR2X2_3200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5834_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5835_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5836_));
OR2X2 OR2X2_3201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5833_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5836_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5837_));
OR2X2 OR2X2_3202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5830_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5837_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5838_));
OR2X2 OR2X2_3203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5838_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5823_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5839_));
OR2X2 OR2X2_3204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5808_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5839_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_3_));
OR2X2 OR2X2_3205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5842_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5841_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5843_));
OR2X2 OR2X2_3206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5844_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5845_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5846_));
OR2X2 OR2X2_3207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5846_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5843_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5847_));
OR2X2 OR2X2_3208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5848_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5849_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5850_));
OR2X2 OR2X2_3209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5851_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5852_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5853_));
OR2X2 OR2X2_321 ( .A(_abc_44694_new_n1602_), .B(_abc_44694_new_n1278__bF_buf1), .Y(_abc_44694_new_n1603_));
OR2X2 OR2X2_3210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5853_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5850_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5854_));
OR2X2 OR2X2_3211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5854_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5847_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5855_));
OR2X2 OR2X2_3212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5857_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5858_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5859_));
OR2X2 OR2X2_3213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5859_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5856_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5860_));
OR2X2 OR2X2_3214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5861_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5862_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5863_));
OR2X2 OR2X2_3215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5865_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5864_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5866_));
OR2X2 OR2X2_3216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5863_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5866_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5867_));
OR2X2 OR2X2_3217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5867_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5860_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5868_));
OR2X2 OR2X2_3218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5868_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5855_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5869_));
OR2X2 OR2X2_3219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5871_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5870_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5872_));
OR2X2 OR2X2_322 ( .A(_abc_44694_new_n1604_), .B(_abc_44694_new_n1605_), .Y(_abc_44694_new_n1606_));
OR2X2 OR2X2_3220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5873_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5874_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5875_));
OR2X2 OR2X2_3221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5875_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5872_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5876_));
OR2X2 OR2X2_3222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5877_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5878_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5879_));
OR2X2 OR2X2_3223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5880_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5881_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5882_));
OR2X2 OR2X2_3224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5879_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5882_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5883_));
OR2X2 OR2X2_3225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5883_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5876_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5884_));
OR2X2 OR2X2_3226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5885_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5886_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5887_));
OR2X2 OR2X2_3227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5888_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5890_));
OR2X2 OR2X2_3228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5887_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5890_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5891_));
OR2X2 OR2X2_3229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5892_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5893_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5894_));
OR2X2 OR2X2_323 ( .A(_abc_44694_new_n1334__bF_buf2), .B(_abc_44694_new_n1606_), .Y(_abc_44694_new_n1607_));
OR2X2 OR2X2_3230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5895_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5896_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5897_));
OR2X2 OR2X2_3231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5894_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5897_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5898_));
OR2X2 OR2X2_3232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5891_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5898_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5899_));
OR2X2 OR2X2_3233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5899_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5884_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5900_));
OR2X2 OR2X2_3234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5869_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5900_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_4_));
OR2X2 OR2X2_3235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5903_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5902_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5904_));
OR2X2 OR2X2_3236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5905_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5906_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5907_));
OR2X2 OR2X2_3237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5907_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5904_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5908_));
OR2X2 OR2X2_3238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5909_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5910_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5911_));
OR2X2 OR2X2_3239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5912_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5914_));
OR2X2 OR2X2_324 ( .A(_abc_44694_new_n1580_), .B(_abc_44694_new_n1609_), .Y(_abc_44694_new_n1610_));
OR2X2 OR2X2_3240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5914_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5911_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5915_));
OR2X2 OR2X2_3241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5915_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5908_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5916_));
OR2X2 OR2X2_3242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5918_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5919_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5920_));
OR2X2 OR2X2_3243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5920_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5917_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5921_));
OR2X2 OR2X2_3244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5922_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5923_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5924_));
OR2X2 OR2X2_3245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5926_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5925_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5927_));
OR2X2 OR2X2_3246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5924_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5927_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5928_));
OR2X2 OR2X2_3247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5928_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5921_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5929_));
OR2X2 OR2X2_3248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5929_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5916_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5930_));
OR2X2 OR2X2_3249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5932_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5931_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5933_));
OR2X2 OR2X2_325 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_7_), .Y(_abc_44694_new_n1611_));
OR2X2 OR2X2_3250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5934_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5935_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5936_));
OR2X2 OR2X2_3251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5936_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5933_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5937_));
OR2X2 OR2X2_3252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5938_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5939_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5940_));
OR2X2 OR2X2_3253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5941_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5942_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5943_));
OR2X2 OR2X2_3254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5940_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5943_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5944_));
OR2X2 OR2X2_3255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5944_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5937_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5945_));
OR2X2 OR2X2_3256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5946_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5947_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5948_));
OR2X2 OR2X2_3257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5949_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5950_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5951_));
OR2X2 OR2X2_3258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5948_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5951_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5952_));
OR2X2 OR2X2_3259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5953_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5954_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5955_));
OR2X2 OR2X2_326 ( .A(_abc_44694_new_n1576_), .B(pc_q_8_), .Y(_abc_44694_new_n1614_));
OR2X2 OR2X2_3260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5956_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5957_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5958_));
OR2X2 OR2X2_3261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5955_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5959_));
OR2X2 OR2X2_3262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5952_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5959_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5960_));
OR2X2 OR2X2_3263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5960_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5945_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5961_));
OR2X2 OR2X2_3264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5930_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5961_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_5_));
OR2X2 OR2X2_3265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5964_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5963_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5965_));
OR2X2 OR2X2_3266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5966_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5967_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5968_));
OR2X2 OR2X2_3267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5968_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5965_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5969_));
OR2X2 OR2X2_3268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5970_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5971_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5972_));
OR2X2 OR2X2_3269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5973_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5974_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5975_));
OR2X2 OR2X2_327 ( .A(_abc_44694_new_n1617_), .B(_abc_44694_new_n1210__bF_buf1), .Y(_abc_44694_new_n1618_));
OR2X2 OR2X2_3270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5975_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5972_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5976_));
OR2X2 OR2X2_3271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5976_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5969_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5977_));
OR2X2 OR2X2_3272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5979_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5980_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5981_));
OR2X2 OR2X2_3273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5981_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5978_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5982_));
OR2X2 OR2X2_3274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5983_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5984_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5985_));
OR2X2 OR2X2_3275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5987_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5986_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5988_));
OR2X2 OR2X2_3276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5985_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5988_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5989_));
OR2X2 OR2X2_3277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5989_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5982_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5990_));
OR2X2 OR2X2_3278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5990_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5977_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5991_));
OR2X2 OR2X2_3279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5993_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5992_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5994_));
OR2X2 OR2X2_328 ( .A(_abc_44694_new_n1399__bF_buf2), .B(_abc_44694_new_n1617_), .Y(_abc_44694_new_n1620_));
OR2X2 OR2X2_3280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5995_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5996_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5997_));
OR2X2 OR2X2_3281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5997_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5994_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n5998_));
OR2X2 OR2X2_3282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5999_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6000_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6001_));
OR2X2 OR2X2_3283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6002_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6003_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6004_));
OR2X2 OR2X2_3284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6001_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6004_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6005_));
OR2X2 OR2X2_3285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6005_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n5998_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6006_));
OR2X2 OR2X2_3286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6007_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6008_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6009_));
OR2X2 OR2X2_3287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6010_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6011_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6012_));
OR2X2 OR2X2_3288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6009_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6012_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6013_));
OR2X2 OR2X2_3289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6014_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6015_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6016_));
OR2X2 OR2X2_329 ( .A(_abc_44694_new_n1590_), .B(_abc_44694_new_n1623_), .Y(_abc_44694_new_n1624_));
OR2X2 OR2X2_3290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6017_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6018_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6019_));
OR2X2 OR2X2_3291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6016_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6019_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6020_));
OR2X2 OR2X2_3292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6013_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6020_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6021_));
OR2X2 OR2X2_3293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6021_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6006_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6022_));
OR2X2 OR2X2_3294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n5991_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6022_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_6_));
OR2X2 OR2X2_3295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6025_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6024_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6026_));
OR2X2 OR2X2_3296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6027_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6028_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6029_));
OR2X2 OR2X2_3297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6029_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6026_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6030_));
OR2X2 OR2X2_3298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6031_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6032_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6033_));
OR2X2 OR2X2_3299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6034_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6035_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6036_));
OR2X2 OR2X2_33 ( .A(_abc_44694_new_n738_), .B(_abc_44694_new_n741_), .Y(_abc_44694_new_n742_));
OR2X2 OR2X2_330 ( .A(alu_op_r_4_), .B(pc_q_8_), .Y(_abc_44694_new_n1625_));
OR2X2 OR2X2_3300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6036_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6033_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6037_));
OR2X2 OR2X2_3301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6037_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6030_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6038_));
OR2X2 OR2X2_3302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6040_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6041_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6042_));
OR2X2 OR2X2_3303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6042_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6039_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6043_));
OR2X2 OR2X2_3304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6044_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6045_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6046_));
OR2X2 OR2X2_3305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6048_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6047_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6049_));
OR2X2 OR2X2_3306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6046_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6049_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6050_));
OR2X2 OR2X2_3307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6050_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6043_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6051_));
OR2X2 OR2X2_3308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6051_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6038_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6052_));
OR2X2 OR2X2_3309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6053_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6055_));
OR2X2 OR2X2_331 ( .A(_abc_44694_new_n1624_), .B(_abc_44694_new_n1628_), .Y(_abc_44694_new_n1629_));
OR2X2 OR2X2_3310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6056_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6058_));
OR2X2 OR2X2_3311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6058_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6055_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6059_));
OR2X2 OR2X2_3312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6060_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6062_));
OR2X2 OR2X2_3313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6063_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6064_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6065_));
OR2X2 OR2X2_3314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6062_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6065_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6066_));
OR2X2 OR2X2_3315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6066_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6067_));
OR2X2 OR2X2_3316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6068_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6069_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6070_));
OR2X2 OR2X2_3317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6071_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6072_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6073_));
OR2X2 OR2X2_3318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6070_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6073_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6074_));
OR2X2 OR2X2_3319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6075_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6076_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6077_));
OR2X2 OR2X2_332 ( .A(_abc_44694_new_n1633_), .B(_abc_44694_new_n1621_), .Y(_abc_44694_new_n1634_));
OR2X2 OR2X2_3320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6078_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6079_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6080_));
OR2X2 OR2X2_3321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6077_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6080_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6081_));
OR2X2 OR2X2_3322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6074_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6081_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6082_));
OR2X2 OR2X2_3323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6082_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6067_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6083_));
OR2X2 OR2X2_3324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6052_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6083_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_7_));
OR2X2 OR2X2_3325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6086_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6085_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6087_));
OR2X2 OR2X2_3326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6088_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6089_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6090_));
OR2X2 OR2X2_3327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6090_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6087_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6091_));
OR2X2 OR2X2_3328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6092_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6093_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6094_));
OR2X2 OR2X2_3329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6095_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6096_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6097_));
OR2X2 OR2X2_333 ( .A(_abc_44694_new_n1400__bF_buf3), .B(_abc_44694_new_n1636_), .Y(_abc_44694_new_n1637_));
OR2X2 OR2X2_3330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6097_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6094_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6098_));
OR2X2 OR2X2_3331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6098_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6091_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6099_));
OR2X2 OR2X2_3332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6101_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6103_));
OR2X2 OR2X2_3333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6103_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6100_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6104_));
OR2X2 OR2X2_3334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6105_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6106_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6107_));
OR2X2 OR2X2_3335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6109_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6108_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6110_));
OR2X2 OR2X2_3336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6107_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6111_));
OR2X2 OR2X2_3337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6111_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6104_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6112_));
OR2X2 OR2X2_3338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6112_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6099_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6113_));
OR2X2 OR2X2_3339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6115_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6114_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6116_));
OR2X2 OR2X2_334 ( .A(_abc_44694_new_n1635_), .B(_abc_44694_new_n1637_), .Y(_abc_44694_new_n1638_));
OR2X2 OR2X2_3340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6117_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6118_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6119_));
OR2X2 OR2X2_3341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6119_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6120_));
OR2X2 OR2X2_3342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6121_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6122_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6123_));
OR2X2 OR2X2_3343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6124_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6125_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6126_));
OR2X2 OR2X2_3344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6123_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6126_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6127_));
OR2X2 OR2X2_3345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6127_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6128_));
OR2X2 OR2X2_3346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6129_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6131_));
OR2X2 OR2X2_3347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6132_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6133_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6134_));
OR2X2 OR2X2_3348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6131_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6134_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6135_));
OR2X2 OR2X2_3349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6136_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6137_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6138_));
OR2X2 OR2X2_335 ( .A(_abc_44694_new_n1639_), .B(_abc_44694_new_n1278__bF_buf0), .Y(_abc_44694_new_n1640_));
OR2X2 OR2X2_3350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6139_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6141_));
OR2X2 OR2X2_3351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6138_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6141_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6142_));
OR2X2 OR2X2_3352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6135_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6142_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6143_));
OR2X2 OR2X2_3353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6143_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6128_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6144_));
OR2X2 OR2X2_3354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6113_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6144_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_8_));
OR2X2 OR2X2_3355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6147_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6146_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6148_));
OR2X2 OR2X2_3356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6149_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6151_));
OR2X2 OR2X2_3357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6151_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6148_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6152_));
OR2X2 OR2X2_3358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6153_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6154_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6155_));
OR2X2 OR2X2_3359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6156_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6157_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6158_));
OR2X2 OR2X2_336 ( .A(_abc_44694_new_n1641_), .B(_abc_44694_new_n1642_), .Y(_abc_44694_new_n1643_));
OR2X2 OR2X2_3360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6158_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6159_));
OR2X2 OR2X2_3361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6159_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6152_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6160_));
OR2X2 OR2X2_3362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6162_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6163_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6164_));
OR2X2 OR2X2_3363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6164_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6161_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6165_));
OR2X2 OR2X2_3364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6166_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6167_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6168_));
OR2X2 OR2X2_3365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6170_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6169_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6171_));
OR2X2 OR2X2_3366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6168_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6171_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6172_));
OR2X2 OR2X2_3367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6172_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6173_));
OR2X2 OR2X2_3368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6173_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6174_));
OR2X2 OR2X2_3369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6176_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6177_));
OR2X2 OR2X2_337 ( .A(_abc_44694_new_n1334__bF_buf1), .B(_abc_44694_new_n1643_), .Y(_abc_44694_new_n1644_));
OR2X2 OR2X2_3370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6178_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6179_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6180_));
OR2X2 OR2X2_3371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6180_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6177_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6181_));
OR2X2 OR2X2_3372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6182_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6183_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6184_));
OR2X2 OR2X2_3373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6185_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6186_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6187_));
OR2X2 OR2X2_3374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6184_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6187_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6188_));
OR2X2 OR2X2_3375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6188_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6181_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6189_));
OR2X2 OR2X2_3376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6190_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6191_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6192_));
OR2X2 OR2X2_3377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6193_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6194_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6195_));
OR2X2 OR2X2_3378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6192_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6196_));
OR2X2 OR2X2_3379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6197_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6198_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6199_));
OR2X2 OR2X2_338 ( .A(_abc_44694_new_n1646_), .B(_abc_44694_new_n1619_), .Y(_abc_44694_new_n1647_));
OR2X2 OR2X2_3380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6200_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6201_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6202_));
OR2X2 OR2X2_3381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6199_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6202_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6203_));
OR2X2 OR2X2_3382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6196_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6203_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6204_));
OR2X2 OR2X2_3383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6204_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6189_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6205_));
OR2X2 OR2X2_3384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6174_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6205_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_9_));
OR2X2 OR2X2_3385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6208_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6207_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6209_));
OR2X2 OR2X2_3386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6210_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6211_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6212_));
OR2X2 OR2X2_3387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6212_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6209_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6213_));
OR2X2 OR2X2_3388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6214_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6215_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6216_));
OR2X2 OR2X2_3389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6217_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6218_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6219_));
OR2X2 OR2X2_339 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_8_), .Y(_abc_44694_new_n1648_));
OR2X2 OR2X2_3390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6219_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6216_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6220_));
OR2X2 OR2X2_3391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6220_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6213_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6221_));
OR2X2 OR2X2_3392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6223_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6224_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6225_));
OR2X2 OR2X2_3393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6225_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6222_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6226_));
OR2X2 OR2X2_3394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6228_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6229_));
OR2X2 OR2X2_3395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6231_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6232_));
OR2X2 OR2X2_3396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6229_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6232_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6233_));
OR2X2 OR2X2_3397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6233_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6226_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6234_));
OR2X2 OR2X2_3398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6234_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6221_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6235_));
OR2X2 OR2X2_3399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6237_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6236_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6238_));
OR2X2 OR2X2_34 ( .A(_abc_44694_new_n673__bF_buf1), .B(_abc_44694_new_n742_), .Y(_abc_44694_new_n743_));
OR2X2 OR2X2_340 ( .A(_abc_44694_new_n1615_), .B(pc_q_9_), .Y(_abc_44694_new_n1651_));
OR2X2 OR2X2_3400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6239_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6241_));
OR2X2 OR2X2_3401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6241_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6238_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6242_));
OR2X2 OR2X2_3402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6243_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6244_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6245_));
OR2X2 OR2X2_3403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6246_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6247_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6248_));
OR2X2 OR2X2_3404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6245_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6248_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6249_));
OR2X2 OR2X2_3405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6249_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6242_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6250_));
OR2X2 OR2X2_3406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6251_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6252_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6253_));
OR2X2 OR2X2_3407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6254_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6256_));
OR2X2 OR2X2_3408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6253_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6256_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6257_));
OR2X2 OR2X2_3409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6258_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6259_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6260_));
OR2X2 OR2X2_341 ( .A(_abc_44694_new_n1654_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n1655_));
OR2X2 OR2X2_3410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6261_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6262_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6263_));
OR2X2 OR2X2_3411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6260_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6263_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6264_));
OR2X2 OR2X2_3412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6264_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6265_));
OR2X2 OR2X2_3413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6265_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6266_));
OR2X2 OR2X2_3414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6235_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6266_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_10_));
OR2X2 OR2X2_3415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6269_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6268_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6270_));
OR2X2 OR2X2_3416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6271_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6272_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6273_));
OR2X2 OR2X2_3417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6273_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6270_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6274_));
OR2X2 OR2X2_3418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6275_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6276_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6277_));
OR2X2 OR2X2_3419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6278_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6279_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6280_));
OR2X2 OR2X2_342 ( .A(_abc_44694_new_n1399__bF_buf1), .B(_abc_44694_new_n1654_), .Y(_abc_44694_new_n1657_));
OR2X2 OR2X2_3420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6280_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6277_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6281_));
OR2X2 OR2X2_3421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6281_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6274_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6282_));
OR2X2 OR2X2_3422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6284_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6285_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6286_));
OR2X2 OR2X2_3423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6286_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6283_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6287_));
OR2X2 OR2X2_3424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6288_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6289_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6290_));
OR2X2 OR2X2_3425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6292_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6291_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6293_));
OR2X2 OR2X2_3426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6290_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6293_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6294_));
OR2X2 OR2X2_3427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6294_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6287_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6295_));
OR2X2 OR2X2_3428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6295_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6282_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6296_));
OR2X2 OR2X2_3429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6298_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6297_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6299_));
OR2X2 OR2X2_343 ( .A(alu_op_r_5_), .B(pc_q_9_), .Y(_abc_44694_new_n1661_));
OR2X2 OR2X2_3430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6300_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6301_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6302_));
OR2X2 OR2X2_3431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6302_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6299_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6303_));
OR2X2 OR2X2_3432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6304_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6305_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6306_));
OR2X2 OR2X2_3433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6307_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6308_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6309_));
OR2X2 OR2X2_3434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6306_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6309_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6310_));
OR2X2 OR2X2_3435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6310_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6303_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6311_));
OR2X2 OR2X2_3436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6312_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6313_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6314_));
OR2X2 OR2X2_3437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6315_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6316_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6317_));
OR2X2 OR2X2_3438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6314_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6317_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6318_));
OR2X2 OR2X2_3439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6319_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6320_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6321_));
OR2X2 OR2X2_344 ( .A(_abc_44694_new_n1664_), .B(_abc_44694_new_n1626_), .Y(_abc_44694_new_n1665_));
OR2X2 OR2X2_3440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6322_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6323_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6324_));
OR2X2 OR2X2_3441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6321_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6324_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6325_));
OR2X2 OR2X2_3442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6318_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6325_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6326_));
OR2X2 OR2X2_3443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6326_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6311_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6327_));
OR2X2 OR2X2_3444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6296_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6327_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_11_));
OR2X2 OR2X2_3445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6330_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6329_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6331_));
OR2X2 OR2X2_3446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6332_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6333_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6334_));
OR2X2 OR2X2_3447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6334_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6331_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6335_));
OR2X2 OR2X2_3448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6336_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6337_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6338_));
OR2X2 OR2X2_3449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6339_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6340_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6341_));
OR2X2 OR2X2_345 ( .A(_abc_44694_new_n1630_), .B(_abc_44694_new_n1665_), .Y(_abc_44694_new_n1666_));
OR2X2 OR2X2_3450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6341_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6338_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6342_));
OR2X2 OR2X2_3451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6342_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6335_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6343_));
OR2X2 OR2X2_3452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6345_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6346_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6347_));
OR2X2 OR2X2_3453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6347_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6344_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6348_));
OR2X2 OR2X2_3454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6349_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6350_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6351_));
OR2X2 OR2X2_3455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6353_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6352_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6354_));
OR2X2 OR2X2_3456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6351_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6354_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6355_));
OR2X2 OR2X2_3457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6355_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6348_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6356_));
OR2X2 OR2X2_3458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6356_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6357_));
OR2X2 OR2X2_3459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6359_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6358_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6360_));
OR2X2 OR2X2_346 ( .A(_abc_44694_new_n1673_), .B(inst_trap_w), .Y(_abc_44694_new_n1674_));
OR2X2 OR2X2_3460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6361_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6362_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6363_));
OR2X2 OR2X2_3461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6363_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6360_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6364_));
OR2X2 OR2X2_3462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6365_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6366_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6367_));
OR2X2 OR2X2_3463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6368_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6369_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6370_));
OR2X2 OR2X2_3464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6371_));
OR2X2 OR2X2_3465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6371_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6364_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6372_));
OR2X2 OR2X2_3466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6373_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6374_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6375_));
OR2X2 OR2X2_3467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6376_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6377_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6378_));
OR2X2 OR2X2_3468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6375_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6378_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6379_));
OR2X2 OR2X2_3469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6380_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6381_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6382_));
OR2X2 OR2X2_347 ( .A(_abc_44694_new_n1675_), .B(_abc_44694_new_n1658_), .Y(_abc_44694_new_n1676_));
OR2X2 OR2X2_3470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6383_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6384_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6385_));
OR2X2 OR2X2_3471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6382_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6385_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6386_));
OR2X2 OR2X2_3472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6379_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6386_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6387_));
OR2X2 OR2X2_3473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6387_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6372_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6388_));
OR2X2 OR2X2_3474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6357_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6388_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_12_));
OR2X2 OR2X2_3475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6391_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6390_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6392_));
OR2X2 OR2X2_3476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6393_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6394_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6395_));
OR2X2 OR2X2_3477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6395_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6392_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6396_));
OR2X2 OR2X2_3478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6397_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6398_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6399_));
OR2X2 OR2X2_3479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6400_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6401_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6402_));
OR2X2 OR2X2_348 ( .A(_abc_44694_new_n1400__bF_buf2), .B(_abc_44694_new_n1678_), .Y(_abc_44694_new_n1679_));
OR2X2 OR2X2_3480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6402_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6399_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6403_));
OR2X2 OR2X2_3481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6403_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6396_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6404_));
OR2X2 OR2X2_3482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6406_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6407_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6408_));
OR2X2 OR2X2_3483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6408_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6405_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6409_));
OR2X2 OR2X2_3484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6410_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6411_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6412_));
OR2X2 OR2X2_3485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6414_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6413_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6415_));
OR2X2 OR2X2_3486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6412_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6415_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6416_));
OR2X2 OR2X2_3487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6416_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6409_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6417_));
OR2X2 OR2X2_3488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6417_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6404_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6418_));
OR2X2 OR2X2_3489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6420_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6421_));
OR2X2 OR2X2_349 ( .A(_abc_44694_new_n1677_), .B(_abc_44694_new_n1679_), .Y(_abc_44694_new_n1680_));
OR2X2 OR2X2_3490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6422_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6423_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6424_));
OR2X2 OR2X2_3491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6424_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6421_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6425_));
OR2X2 OR2X2_3492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6426_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6427_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6428_));
OR2X2 OR2X2_3493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6429_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6430_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6431_));
OR2X2 OR2X2_3494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6428_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6431_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6432_));
OR2X2 OR2X2_3495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6432_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6425_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6433_));
OR2X2 OR2X2_3496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6434_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6436_));
OR2X2 OR2X2_3497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6437_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6438_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6439_));
OR2X2 OR2X2_3498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6436_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6439_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6440_));
OR2X2 OR2X2_3499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6441_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6442_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6443_));
OR2X2 OR2X2_35 ( .A(_abc_44694_new_n745_), .B(_abc_44694_new_n731_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_3_));
OR2X2 OR2X2_350 ( .A(_abc_44694_new_n1681_), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n1682_));
OR2X2 OR2X2_3500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6444_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6445_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6446_));
OR2X2 OR2X2_3501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6443_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6446_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6447_));
OR2X2 OR2X2_3502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6440_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6447_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6448_));
OR2X2 OR2X2_3503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6448_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6433_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6449_));
OR2X2 OR2X2_3504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6418_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6449_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_13_));
OR2X2 OR2X2_3505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6452_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6451_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6453_));
OR2X2 OR2X2_3506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6454_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6455_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6456_));
OR2X2 OR2X2_3507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6456_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6453_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6457_));
OR2X2 OR2X2_3508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6458_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6459_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6460_));
OR2X2 OR2X2_3509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6461_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6462_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6463_));
OR2X2 OR2X2_351 ( .A(_abc_44694_new_n1683_), .B(_abc_44694_new_n1684_), .Y(_abc_44694_new_n1685_));
OR2X2 OR2X2_3510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6463_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6460_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6464_));
OR2X2 OR2X2_3511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6464_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6457_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6465_));
OR2X2 OR2X2_3512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6467_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6469_));
OR2X2 OR2X2_3513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6469_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6466_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6470_));
OR2X2 OR2X2_3514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6472_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6473_));
OR2X2 OR2X2_3515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6475_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6474_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6476_));
OR2X2 OR2X2_3516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6473_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6476_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6477_));
OR2X2 OR2X2_3517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6477_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6470_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6478_));
OR2X2 OR2X2_3518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6478_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6465_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6479_));
OR2X2 OR2X2_3519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6481_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6480_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6482_));
OR2X2 OR2X2_352 ( .A(_abc_44694_new_n1334__bF_buf0), .B(_abc_44694_new_n1685_), .Y(_abc_44694_new_n1686_));
OR2X2 OR2X2_3520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6483_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6484_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6485_));
OR2X2 OR2X2_3521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6485_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6482_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6486_));
OR2X2 OR2X2_3522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6487_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6488_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6489_));
OR2X2 OR2X2_3523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6490_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6491_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6492_));
OR2X2 OR2X2_3524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6489_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6492_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6493_));
OR2X2 OR2X2_3525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6493_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6486_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6494_));
OR2X2 OR2X2_3526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6496_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6497_));
OR2X2 OR2X2_3527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6498_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6499_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6500_));
OR2X2 OR2X2_3528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6497_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6500_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6501_));
OR2X2 OR2X2_3529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6502_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6503_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6504_));
OR2X2 OR2X2_353 ( .A(_abc_44694_new_n1688_), .B(_abc_44694_new_n1656_), .Y(_abc_44694_new_n1689_));
OR2X2 OR2X2_3530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6505_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6506_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6507_));
OR2X2 OR2X2_3531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6504_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6507_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6508_));
OR2X2 OR2X2_3532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6501_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6508_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6509_));
OR2X2 OR2X2_3533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6509_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6494_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6510_));
OR2X2 OR2X2_3534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6479_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6510_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_14_));
OR2X2 OR2X2_3535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6513_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6512_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6514_));
OR2X2 OR2X2_3536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6516_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6517_));
OR2X2 OR2X2_3537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6517_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6514_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6518_));
OR2X2 OR2X2_3538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6519_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6520_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6521_));
OR2X2 OR2X2_3539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6522_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6523_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6524_));
OR2X2 OR2X2_354 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(epc_q_9_), .Y(_abc_44694_new_n1690_));
OR2X2 OR2X2_3540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6524_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6521_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6525_));
OR2X2 OR2X2_3541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6525_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6518_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6526_));
OR2X2 OR2X2_3542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6528_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6529_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6530_));
OR2X2 OR2X2_3543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6530_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6527_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6531_));
OR2X2 OR2X2_3544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6532_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6533_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6534_));
OR2X2 OR2X2_3545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6536_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6535_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6537_));
OR2X2 OR2X2_3546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6534_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6537_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6538_));
OR2X2 OR2X2_3547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6538_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6531_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6539_));
OR2X2 OR2X2_3548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6539_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6526_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6540_));
OR2X2 OR2X2_3549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6542_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6543_));
OR2X2 OR2X2_355 ( .A(_abc_44694_new_n1652_), .B(pc_q_10_), .Y(_abc_44694_new_n1693_));
OR2X2 OR2X2_3550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6544_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6545_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6546_));
OR2X2 OR2X2_3551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6546_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6547_));
OR2X2 OR2X2_3552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6548_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6549_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6550_));
OR2X2 OR2X2_3553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6551_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6552_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6553_));
OR2X2 OR2X2_3554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6550_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6554_));
OR2X2 OR2X2_3555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6554_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6547_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6555_));
OR2X2 OR2X2_3556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6557_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6558_));
OR2X2 OR2X2_3557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6559_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6560_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6561_));
OR2X2 OR2X2_3558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6558_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6561_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6562_));
OR2X2 OR2X2_3559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6563_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6564_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6565_));
OR2X2 OR2X2_356 ( .A(_abc_44694_new_n1696_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n1697_));
OR2X2 OR2X2_3560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6566_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6567_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6568_));
OR2X2 OR2X2_3561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6565_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6568_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6569_));
OR2X2 OR2X2_3562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6562_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6569_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6570_));
OR2X2 OR2X2_3563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6570_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6555_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6571_));
OR2X2 OR2X2_3564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6540_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6571_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_15_));
OR2X2 OR2X2_3565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6574_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6573_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6575_));
OR2X2 OR2X2_3566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6576_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6577_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6578_));
OR2X2 OR2X2_3567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6578_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6575_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6579_));
OR2X2 OR2X2_3568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6580_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6581_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6582_));
OR2X2 OR2X2_3569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6583_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6584_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6585_));
OR2X2 OR2X2_357 ( .A(_abc_44694_new_n1667_), .B(_abc_44694_new_n1662_), .Y(_abc_44694_new_n1699_));
OR2X2 OR2X2_3570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6585_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6582_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6586_));
OR2X2 OR2X2_3571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6586_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6579_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6587_));
OR2X2 OR2X2_3572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6589_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6590_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6591_));
OR2X2 OR2X2_3573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6591_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6592_));
OR2X2 OR2X2_3574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6593_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6595_));
OR2X2 OR2X2_3575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6597_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6596_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6598_));
OR2X2 OR2X2_3576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6595_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6599_));
OR2X2 OR2X2_3577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6599_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6600_));
OR2X2 OR2X2_3578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6600_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6587_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6601_));
OR2X2 OR2X2_3579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6603_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6604_));
OR2X2 OR2X2_358 ( .A(alu_op_r_6_), .B(pc_q_10_), .Y(_abc_44694_new_n1703_));
OR2X2 OR2X2_3580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6605_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6607_));
OR2X2 OR2X2_3581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6607_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6608_));
OR2X2 OR2X2_3582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6609_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6610_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6611_));
OR2X2 OR2X2_3583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6612_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6613_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6614_));
OR2X2 OR2X2_3584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6611_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6614_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6615_));
OR2X2 OR2X2_3585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6615_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6608_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6616_));
OR2X2 OR2X2_3586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6617_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6619_));
OR2X2 OR2X2_3587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6620_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6621_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6622_));
OR2X2 OR2X2_3588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6619_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6622_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6623_));
OR2X2 OR2X2_3589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6624_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6625_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6626_));
OR2X2 OR2X2_359 ( .A(_abc_44694_new_n1702_), .B(_abc_44694_new_n1706_), .Y(_abc_44694_new_n1709_));
OR2X2 OR2X2_3590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6627_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6629_));
OR2X2 OR2X2_3591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6626_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6629_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6630_));
OR2X2 OR2X2_3592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6623_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6630_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6631_));
OR2X2 OR2X2_3593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6631_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6632_));
OR2X2 OR2X2_3594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6601_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6632_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_16_));
OR2X2 OR2X2_3595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6635_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6634_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6636_));
OR2X2 OR2X2_3596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6637_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6639_));
OR2X2 OR2X2_3597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6639_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6636_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6640_));
OR2X2 OR2X2_3598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6641_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6642_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6643_));
OR2X2 OR2X2_3599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6644_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6645_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6646_));
OR2X2 OR2X2_36 ( .A(_abc_44694_new_n748_), .B(_abc_44694_new_n749_), .Y(_abc_44694_new_n750_));
OR2X2 OR2X2_360 ( .A(_abc_44694_new_n1710_), .B(_abc_44694_new_n1389_), .Y(_abc_44694_new_n1711_));
OR2X2 OR2X2_3600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6646_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6643_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6647_));
OR2X2 OR2X2_3601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6647_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6648_));
OR2X2 OR2X2_3602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6650_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6652_));
OR2X2 OR2X2_3603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6652_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6649_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6653_));
OR2X2 OR2X2_3604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6654_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6655_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6656_));
OR2X2 OR2X2_3605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6658_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6657_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6659_));
OR2X2 OR2X2_3606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6656_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6660_));
OR2X2 OR2X2_3607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6660_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6653_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6661_));
OR2X2 OR2X2_3608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6661_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6662_));
OR2X2 OR2X2_3609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6664_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6663_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6665_));
OR2X2 OR2X2_361 ( .A(_abc_44694_new_n1021_), .B(epc_q_10_), .Y(_abc_44694_new_n1712_));
OR2X2 OR2X2_3610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6666_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6667_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6668_));
OR2X2 OR2X2_3611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6668_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6665_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6669_));
OR2X2 OR2X2_3612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6670_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6671_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6672_));
OR2X2 OR2X2_3613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6673_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6674_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6675_));
OR2X2 OR2X2_3614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6672_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6675_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6676_));
OR2X2 OR2X2_3615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6676_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6669_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6677_));
OR2X2 OR2X2_3616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6678_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6679_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6680_));
OR2X2 OR2X2_3617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6681_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6682_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6683_));
OR2X2 OR2X2_3618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6680_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6683_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6684_));
OR2X2 OR2X2_3619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6685_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6686_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6687_));
OR2X2 OR2X2_362 ( .A(_abc_44694_new_n1714_), .B(_abc_44694_new_n1715_), .Y(_abc_44694_new_n1716_));
OR2X2 OR2X2_3620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6688_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6689_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6690_));
OR2X2 OR2X2_3621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6687_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6690_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6691_));
OR2X2 OR2X2_3622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6684_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6691_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6692_));
OR2X2 OR2X2_3623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6692_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6677_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6693_));
OR2X2 OR2X2_3624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6662_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6693_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_17_));
OR2X2 OR2X2_3625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6696_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6695_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6697_));
OR2X2 OR2X2_3626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6698_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6700_));
OR2X2 OR2X2_3627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6700_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6697_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6701_));
OR2X2 OR2X2_3628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6702_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6703_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6704_));
OR2X2 OR2X2_3629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6705_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6706_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6707_));
OR2X2 OR2X2_363 ( .A(_abc_44694_new_n1717_), .B(_abc_44694_new_n1718_), .Y(_abc_44694_new_n1719_));
OR2X2 OR2X2_3630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6707_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6704_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6708_));
OR2X2 OR2X2_3631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6708_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6701_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6709_));
OR2X2 OR2X2_3632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6711_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6712_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6713_));
OR2X2 OR2X2_3633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6713_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6710_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6714_));
OR2X2 OR2X2_3634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6715_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6716_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6717_));
OR2X2 OR2X2_3635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6719_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6718_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6720_));
OR2X2 OR2X2_3636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6717_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6720_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6721_));
OR2X2 OR2X2_3637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6721_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6714_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6722_));
OR2X2 OR2X2_3638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6722_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6709_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6723_));
OR2X2 OR2X2_3639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6725_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6724_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6726_));
OR2X2 OR2X2_364 ( .A(_abc_44694_new_n1719_), .B(_abc_44694_new_n1278__bF_buf4), .Y(_abc_44694_new_n1720_));
OR2X2 OR2X2_3640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6727_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6728_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6729_));
OR2X2 OR2X2_3641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6729_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6726_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6730_));
OR2X2 OR2X2_3642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6731_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6732_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6733_));
OR2X2 OR2X2_3643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6734_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6735_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6736_));
OR2X2 OR2X2_3644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6733_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6736_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6737_));
OR2X2 OR2X2_3645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6737_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6730_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6738_));
OR2X2 OR2X2_3646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6739_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6740_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6741_));
OR2X2 OR2X2_3647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6742_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6743_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6744_));
OR2X2 OR2X2_3648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6741_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6744_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6745_));
OR2X2 OR2X2_3649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6746_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6747_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6748_));
OR2X2 OR2X2_365 ( .A(_abc_44694_new_n1721_), .B(_abc_44694_new_n1722_), .Y(_abc_44694_new_n1723_));
OR2X2 OR2X2_3650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6749_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6750_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6751_));
OR2X2 OR2X2_3651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6748_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6751_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6752_));
OR2X2 OR2X2_3652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6745_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6752_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6753_));
OR2X2 OR2X2_3653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6753_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6738_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6754_));
OR2X2 OR2X2_3654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6723_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6754_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_18_));
OR2X2 OR2X2_3655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6757_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6756_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6758_));
OR2X2 OR2X2_3656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6759_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6760_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6761_));
OR2X2 OR2X2_3657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6761_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6758_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6762_));
OR2X2 OR2X2_3658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6763_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6764_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6765_));
OR2X2 OR2X2_3659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6766_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6767_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6768_));
OR2X2 OR2X2_366 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n1723_), .Y(_abc_44694_new_n1724_));
OR2X2 OR2X2_3660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6768_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6765_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6769_));
OR2X2 OR2X2_3661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6769_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6762_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6770_));
OR2X2 OR2X2_3662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6772_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6773_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6774_));
OR2X2 OR2X2_3663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6774_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6771_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6775_));
OR2X2 OR2X2_3664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6776_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6777_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6778_));
OR2X2 OR2X2_3665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6780_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6779_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6781_));
OR2X2 OR2X2_3666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6778_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6781_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6782_));
OR2X2 OR2X2_3667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6782_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6775_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6783_));
OR2X2 OR2X2_3668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6783_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6770_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6784_));
OR2X2 OR2X2_3669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6786_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6785_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6787_));
OR2X2 OR2X2_367 ( .A(_abc_44694_new_n1726_), .B(_abc_44694_new_n1698_), .Y(_abc_44694_new_n1727_));
OR2X2 OR2X2_3670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6788_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6789_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6790_));
OR2X2 OR2X2_3671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6790_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6787_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6791_));
OR2X2 OR2X2_3672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6792_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6793_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6794_));
OR2X2 OR2X2_3673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6795_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6796_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6797_));
OR2X2 OR2X2_3674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6794_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6797_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6798_));
OR2X2 OR2X2_3675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6798_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6799_));
OR2X2 OR2X2_3676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6800_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6801_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6802_));
OR2X2 OR2X2_3677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6803_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6804_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6805_));
OR2X2 OR2X2_3678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6802_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6805_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6806_));
OR2X2 OR2X2_3679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6807_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6808_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6809_));
OR2X2 OR2X2_368 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(epc_q_10_), .Y(_abc_44694_new_n1728_));
OR2X2 OR2X2_3680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6810_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6811_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6812_));
OR2X2 OR2X2_3681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6809_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6812_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6813_));
OR2X2 OR2X2_3682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6806_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6814_));
OR2X2 OR2X2_3683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6814_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6799_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6815_));
OR2X2 OR2X2_3684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6784_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6815_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_19_));
OR2X2 OR2X2_3685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6818_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6817_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6819_));
OR2X2 OR2X2_3686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6820_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6821_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6822_));
OR2X2 OR2X2_3687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6822_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6819_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6823_));
OR2X2 OR2X2_3688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6824_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6825_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6826_));
OR2X2 OR2X2_3689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6827_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6828_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6829_));
OR2X2 OR2X2_369 ( .A(_abc_44694_new_n1694_), .B(pc_q_11_), .Y(_abc_44694_new_n1731_));
OR2X2 OR2X2_3690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6829_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6826_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6830_));
OR2X2 OR2X2_3691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6830_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6823_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6831_));
OR2X2 OR2X2_3692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6833_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6834_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6835_));
OR2X2 OR2X2_3693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6835_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6832_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6836_));
OR2X2 OR2X2_3694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6837_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6838_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6839_));
OR2X2 OR2X2_3695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6841_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6840_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6842_));
OR2X2 OR2X2_3696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6839_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6842_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6843_));
OR2X2 OR2X2_3697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6843_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6836_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6844_));
OR2X2 OR2X2_3698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6844_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6831_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6845_));
OR2X2 OR2X2_3699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6847_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6846_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6848_));
OR2X2 OR2X2_37 ( .A(_abc_44694_new_n752_), .B(_abc_44694_new_n753_), .Y(_abc_44694_new_n754_));
OR2X2 OR2X2_370 ( .A(_abc_44694_new_n1734_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n1735_));
OR2X2 OR2X2_3700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6849_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6850_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6851_));
OR2X2 OR2X2_3701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6851_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6848_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6852_));
OR2X2 OR2X2_3702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6853_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6854_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6855_));
OR2X2 OR2X2_3703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6856_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6857_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6858_));
OR2X2 OR2X2_3704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6855_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6858_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6859_));
OR2X2 OR2X2_3705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6859_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6852_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6860_));
OR2X2 OR2X2_3706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6861_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6862_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6863_));
OR2X2 OR2X2_3707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6864_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6865_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6866_));
OR2X2 OR2X2_3708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6863_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6866_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6867_));
OR2X2 OR2X2_3709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6868_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6869_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6870_));
OR2X2 OR2X2_371 ( .A(_abc_44694_new_n1399__bF_buf4), .B(_abc_44694_new_n1734_), .Y(_abc_44694_new_n1737_));
OR2X2 OR2X2_3710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6871_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6872_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6873_));
OR2X2 OR2X2_3711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6870_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6873_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6874_));
OR2X2 OR2X2_3712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6867_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6874_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6875_));
OR2X2 OR2X2_3713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6875_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6860_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6876_));
OR2X2 OR2X2_3714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6845_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6876_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_20_));
OR2X2 OR2X2_3715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6879_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6878_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6880_));
OR2X2 OR2X2_3716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6881_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6882_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6883_));
OR2X2 OR2X2_3717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6883_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6880_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6884_));
OR2X2 OR2X2_3718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6885_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6886_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6887_));
OR2X2 OR2X2_3719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6888_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6889_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6890_));
OR2X2 OR2X2_372 ( .A(alu_op_r_7_), .B(pc_q_11_), .Y(_abc_44694_new_n1740_));
OR2X2 OR2X2_3720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6890_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6887_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6891_));
OR2X2 OR2X2_3721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6891_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6884_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6892_));
OR2X2 OR2X2_3722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6894_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6895_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6896_));
OR2X2 OR2X2_3723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6896_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6893_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6897_));
OR2X2 OR2X2_3724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6898_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6899_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6900_));
OR2X2 OR2X2_3725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6902_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6901_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6903_));
OR2X2 OR2X2_3726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6900_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6903_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6904_));
OR2X2 OR2X2_3727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6904_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6897_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6905_));
OR2X2 OR2X2_3728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6905_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6892_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6906_));
OR2X2 OR2X2_3729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6908_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6907_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6909_));
OR2X2 OR2X2_373 ( .A(_abc_44694_new_n1747_), .B(_abc_44694_new_n1744_), .Y(_abc_44694_new_n1748_));
OR2X2 OR2X2_3730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6910_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6911_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6912_));
OR2X2 OR2X2_3731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6912_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6909_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6913_));
OR2X2 OR2X2_3732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6914_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6915_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6916_));
OR2X2 OR2X2_3733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6917_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6918_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6919_));
OR2X2 OR2X2_3734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6916_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6919_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6920_));
OR2X2 OR2X2_3735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6920_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6921_));
OR2X2 OR2X2_3736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6922_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6923_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6924_));
OR2X2 OR2X2_3737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6925_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6926_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6927_));
OR2X2 OR2X2_3738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6924_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6927_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6928_));
OR2X2 OR2X2_3739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6929_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6930_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6931_));
OR2X2 OR2X2_374 ( .A(_abc_44694_new_n1749_), .B(_abc_44694_new_n1738_), .Y(_abc_44694_new_n1750_));
OR2X2 OR2X2_3740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6932_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6933_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6934_));
OR2X2 OR2X2_3741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6931_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6934_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6935_));
OR2X2 OR2X2_3742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6928_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6935_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6936_));
OR2X2 OR2X2_3743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6936_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6921_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6937_));
OR2X2 OR2X2_3744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6906_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6937_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_21_));
OR2X2 OR2X2_3745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6940_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6939_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6941_));
OR2X2 OR2X2_3746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6942_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6943_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6944_));
OR2X2 OR2X2_3747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6944_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6941_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6945_));
OR2X2 OR2X2_3748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6946_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6947_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6948_));
OR2X2 OR2X2_3749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6949_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6950_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6951_));
OR2X2 OR2X2_375 ( .A(_abc_44694_new_n1400__bF_buf0), .B(_abc_44694_new_n1752_), .Y(_abc_44694_new_n1753_));
OR2X2 OR2X2_3750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6951_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6948_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6952_));
OR2X2 OR2X2_3751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6952_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6945_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6953_));
OR2X2 OR2X2_3752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6955_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6956_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6957_));
OR2X2 OR2X2_3753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6957_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6954_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6958_));
OR2X2 OR2X2_3754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6959_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6961_));
OR2X2 OR2X2_3755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6963_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6962_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6964_));
OR2X2 OR2X2_3756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6961_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6964_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6965_));
OR2X2 OR2X2_3757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6965_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6966_));
OR2X2 OR2X2_3758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6966_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6953_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6967_));
OR2X2 OR2X2_3759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6969_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6968_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6970_));
OR2X2 OR2X2_376 ( .A(_abc_44694_new_n1751_), .B(_abc_44694_new_n1753_), .Y(_abc_44694_new_n1754_));
OR2X2 OR2X2_3760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6971_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6972_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6973_));
OR2X2 OR2X2_3761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6973_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6970_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6974_));
OR2X2 OR2X2_3762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6975_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6976_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6977_));
OR2X2 OR2X2_3763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6978_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6979_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6980_));
OR2X2 OR2X2_3764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6977_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6980_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6981_));
OR2X2 OR2X2_3765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6981_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6974_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6982_));
OR2X2 OR2X2_3766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6983_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6984_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6985_));
OR2X2 OR2X2_3767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6986_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6988_));
OR2X2 OR2X2_3768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6985_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6988_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6989_));
OR2X2 OR2X2_3769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6990_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6991_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6992_));
OR2X2 OR2X2_377 ( .A(_abc_44694_new_n1755_), .B(_abc_44694_new_n1278__bF_buf3), .Y(_abc_44694_new_n1756_));
OR2X2 OR2X2_3770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6993_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6994_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6995_));
OR2X2 OR2X2_3771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6992_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6995_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6996_));
OR2X2 OR2X2_3772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6989_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6996_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6997_));
OR2X2 OR2X2_3773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6997_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6982_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n6998_));
OR2X2 OR2X2_3774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n6967_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n6998_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_22_));
OR2X2 OR2X2_3775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7001_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7000_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7002_));
OR2X2 OR2X2_3776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7003_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7004_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7005_));
OR2X2 OR2X2_3777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7005_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7002_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7006_));
OR2X2 OR2X2_3778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7007_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7008_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7009_));
OR2X2 OR2X2_3779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7010_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7011_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7012_));
OR2X2 OR2X2_378 ( .A(_abc_44694_new_n1757_), .B(_abc_44694_new_n1758_), .Y(_abc_44694_new_n1759_));
OR2X2 OR2X2_3780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7012_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7009_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7013_));
OR2X2 OR2X2_3781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7013_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7006_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7014_));
OR2X2 OR2X2_3782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7016_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7017_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7018_));
OR2X2 OR2X2_3783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7018_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7015_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7019_));
OR2X2 OR2X2_3784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7020_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7021_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7022_));
OR2X2 OR2X2_3785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7024_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7023_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7025_));
OR2X2 OR2X2_3786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7022_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7025_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7026_));
OR2X2 OR2X2_3787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7026_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7019_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7027_));
OR2X2 OR2X2_3788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7027_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7014_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7028_));
OR2X2 OR2X2_3789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7030_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7029_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7031_));
OR2X2 OR2X2_379 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n1759_), .Y(_abc_44694_new_n1760_));
OR2X2 OR2X2_3790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7032_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7033_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7034_));
OR2X2 OR2X2_3791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7034_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7031_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7035_));
OR2X2 OR2X2_3792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7036_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7037_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7038_));
OR2X2 OR2X2_3793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7039_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7040_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7041_));
OR2X2 OR2X2_3794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7038_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7041_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7042_));
OR2X2 OR2X2_3795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7042_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7035_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7043_));
OR2X2 OR2X2_3796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7044_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7045_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7046_));
OR2X2 OR2X2_3797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7047_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7048_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7049_));
OR2X2 OR2X2_3798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7046_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7049_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7050_));
OR2X2 OR2X2_3799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7051_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7052_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7053_));
OR2X2 OR2X2_38 ( .A(_abc_44694_new_n755_), .B(_abc_44694_new_n756_), .Y(_abc_44694_new_n757_));
OR2X2 OR2X2_380 ( .A(_abc_44694_new_n1762_), .B(_abc_44694_new_n1736_), .Y(_abc_44694_new_n1763_));
OR2X2 OR2X2_3800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7055_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7056_));
OR2X2 OR2X2_3801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7053_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7056_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7057_));
OR2X2 OR2X2_3802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7050_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7058_));
OR2X2 OR2X2_3803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7058_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7043_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7059_));
OR2X2 OR2X2_3804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7028_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7059_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_23_));
OR2X2 OR2X2_3805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7062_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7061_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7063_));
OR2X2 OR2X2_3806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7064_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7065_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7066_));
OR2X2 OR2X2_3807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7066_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7063_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7067_));
OR2X2 OR2X2_3808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7068_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7069_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7070_));
OR2X2 OR2X2_3809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7071_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7072_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7073_));
OR2X2 OR2X2_381 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_11_), .Y(_abc_44694_new_n1764_));
OR2X2 OR2X2_3810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7073_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7070_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7074_));
OR2X2 OR2X2_3811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7074_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7067_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7075_));
OR2X2 OR2X2_3812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7077_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7078_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7079_));
OR2X2 OR2X2_3813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7079_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7076_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7080_));
OR2X2 OR2X2_3814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7081_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7082_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7083_));
OR2X2 OR2X2_3815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7085_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7084_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7086_));
OR2X2 OR2X2_3816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7083_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7086_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7087_));
OR2X2 OR2X2_3817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7087_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7080_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7088_));
OR2X2 OR2X2_3818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7088_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7075_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7089_));
OR2X2 OR2X2_3819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7091_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7090_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7092_));
OR2X2 OR2X2_382 ( .A(_abc_44694_new_n1732_), .B(pc_q_12_), .Y(_abc_44694_new_n1767_));
OR2X2 OR2X2_3820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7093_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7094_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7095_));
OR2X2 OR2X2_3821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7095_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7092_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7096_));
OR2X2 OR2X2_3822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7097_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7098_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7099_));
OR2X2 OR2X2_3823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7100_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7101_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7102_));
OR2X2 OR2X2_3824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7099_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7103_));
OR2X2 OR2X2_3825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7103_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7096_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7104_));
OR2X2 OR2X2_3826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7105_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7106_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7107_));
OR2X2 OR2X2_3827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7108_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7109_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7110_));
OR2X2 OR2X2_3828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7107_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7111_));
OR2X2 OR2X2_3829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7112_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7113_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7114_));
OR2X2 OR2X2_383 ( .A(_abc_44694_new_n1770_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n1771_));
OR2X2 OR2X2_3830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7115_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7117_));
OR2X2 OR2X2_3831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7114_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7117_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7118_));
OR2X2 OR2X2_3832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7111_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7118_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7119_));
OR2X2 OR2X2_3833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7119_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7104_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7120_));
OR2X2 OR2X2_3834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7089_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7120_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_24_));
OR2X2 OR2X2_3835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7123_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7122_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7124_));
OR2X2 OR2X2_3836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7125_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7126_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7127_));
OR2X2 OR2X2_3837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7127_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7124_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7128_));
OR2X2 OR2X2_3838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7129_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7131_));
OR2X2 OR2X2_3839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7132_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7133_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7134_));
OR2X2 OR2X2_384 ( .A(_abc_44694_new_n1770_), .B(_abc_44694_new_n1399__bF_buf3), .Y(_abc_44694_new_n1773_));
OR2X2 OR2X2_3840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7134_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7131_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7135_));
OR2X2 OR2X2_3841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7135_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7128_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7136_));
OR2X2 OR2X2_3842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7138_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7139_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7140_));
OR2X2 OR2X2_3843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7140_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7137_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7141_));
OR2X2 OR2X2_3844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7142_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7143_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7144_));
OR2X2 OR2X2_3845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7146_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7145_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7147_));
OR2X2 OR2X2_3846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7144_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7147_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7148_));
OR2X2 OR2X2_3847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7148_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7141_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7149_));
OR2X2 OR2X2_3848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7149_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7136_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7150_));
OR2X2 OR2X2_3849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7152_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7151_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7153_));
OR2X2 OR2X2_385 ( .A(_abc_44694_new_n1777_), .B(_abc_44694_new_n1741_), .Y(_abc_44694_new_n1778_));
OR2X2 OR2X2_3850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7154_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7156_));
OR2X2 OR2X2_3851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7156_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7153_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7157_));
OR2X2 OR2X2_3852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7158_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7159_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7160_));
OR2X2 OR2X2_3853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7161_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7162_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7163_));
OR2X2 OR2X2_3854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7160_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7163_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7164_));
OR2X2 OR2X2_3855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7164_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7157_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7165_));
OR2X2 OR2X2_3856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7166_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7167_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7168_));
OR2X2 OR2X2_3857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7169_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7171_));
OR2X2 OR2X2_3858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7168_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7171_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7172_));
OR2X2 OR2X2_3859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7173_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7174_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7175_));
OR2X2 OR2X2_386 ( .A(_abc_44694_new_n1776_), .B(_abc_44694_new_n1778_), .Y(_abc_44694_new_n1779_));
OR2X2 OR2X2_3860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7176_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7177_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7178_));
OR2X2 OR2X2_3861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7175_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7178_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7179_));
OR2X2 OR2X2_3862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7172_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7179_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7180_));
OR2X2 OR2X2_3863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7180_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7181_));
OR2X2 OR2X2_3864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7150_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7181_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_25_));
OR2X2 OR2X2_3865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7184_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7183_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7185_));
OR2X2 OR2X2_3866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7186_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7187_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7188_));
OR2X2 OR2X2_3867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7188_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7189_));
OR2X2 OR2X2_3868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7190_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7191_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7192_));
OR2X2 OR2X2_3869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7193_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7194_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7195_));
OR2X2 OR2X2_387 ( .A(_abc_44694_new_n1781_), .B(_abc_44694_new_n1779_), .Y(_abc_44694_new_n1782_));
OR2X2 OR2X2_3870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7195_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7192_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7196_));
OR2X2 OR2X2_3871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7196_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7189_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7197_));
OR2X2 OR2X2_3872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7199_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7200_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7201_));
OR2X2 OR2X2_3873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7201_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7198_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7202_));
OR2X2 OR2X2_3874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7203_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7204_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7205_));
OR2X2 OR2X2_3875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7207_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7206_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7208_));
OR2X2 OR2X2_3876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7205_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7208_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7209_));
OR2X2 OR2X2_3877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7209_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7202_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7210_));
OR2X2 OR2X2_3878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7210_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7197_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7211_));
OR2X2 OR2X2_3879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7213_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7212_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7214_));
OR2X2 OR2X2_388 ( .A(int32_r_10_), .B(pc_q_12_), .Y(_abc_44694_new_n1783_));
OR2X2 OR2X2_3880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7215_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7216_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7217_));
OR2X2 OR2X2_3881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7217_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7214_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7218_));
OR2X2 OR2X2_3882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7219_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7220_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7221_));
OR2X2 OR2X2_3883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7222_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7223_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7224_));
OR2X2 OR2X2_3884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7221_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7224_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7225_));
OR2X2 OR2X2_3885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7225_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7218_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7226_));
OR2X2 OR2X2_3886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7228_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7229_));
OR2X2 OR2X2_3887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7230_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7231_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7232_));
OR2X2 OR2X2_3888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7229_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7232_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7233_));
OR2X2 OR2X2_3889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7234_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7235_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7236_));
OR2X2 OR2X2_389 ( .A(_abc_44694_new_n1782_), .B(_abc_44694_new_n1786_), .Y(_abc_44694_new_n1787_));
OR2X2 OR2X2_3890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7237_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7238_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7239_));
OR2X2 OR2X2_3891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7236_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7239_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7240_));
OR2X2 OR2X2_3892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7233_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7241_));
OR2X2 OR2X2_3893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7241_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7226_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7242_));
OR2X2 OR2X2_3894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7211_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7242_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_26_));
OR2X2 OR2X2_3895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7245_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7244_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7246_));
OR2X2 OR2X2_3896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7247_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7248_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7249_));
OR2X2 OR2X2_3897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7249_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7246_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7250_));
OR2X2 OR2X2_3898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7251_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7252_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7253_));
OR2X2 OR2X2_3899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7254_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7255_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7256_));
OR2X2 OR2X2_39 ( .A(_abc_44694_new_n754_), .B(_abc_44694_new_n757_), .Y(_abc_44694_new_n758_));
OR2X2 OR2X2_390 ( .A(_abc_44694_new_n1791_), .B(_abc_44694_new_n1774_), .Y(_abc_44694_new_n1792_));
OR2X2 OR2X2_3900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7256_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7253_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7257_));
OR2X2 OR2X2_3901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7258_));
OR2X2 OR2X2_3902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7260_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7261_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7262_));
OR2X2 OR2X2_3903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7262_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7259_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7263_));
OR2X2 OR2X2_3904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7264_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7265_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7266_));
OR2X2 OR2X2_3905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7268_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7267_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7269_));
OR2X2 OR2X2_3906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7266_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7270_));
OR2X2 OR2X2_3907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7270_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7263_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7271_));
OR2X2 OR2X2_3908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7271_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7258_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7272_));
OR2X2 OR2X2_3909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7274_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7273_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7275_));
OR2X2 OR2X2_391 ( .A(_abc_44694_new_n1400__bF_buf4), .B(_abc_44694_new_n1794_), .Y(_abc_44694_new_n1795_));
OR2X2 OR2X2_3910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7276_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7277_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7278_));
OR2X2 OR2X2_3911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7278_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7275_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7279_));
OR2X2 OR2X2_3912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7280_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7281_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7282_));
OR2X2 OR2X2_3913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7283_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7284_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7285_));
OR2X2 OR2X2_3914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7282_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7285_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7286_));
OR2X2 OR2X2_3915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7286_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7279_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7287_));
OR2X2 OR2X2_3916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7288_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7289_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7290_));
OR2X2 OR2X2_3917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7291_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7292_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7293_));
OR2X2 OR2X2_3918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7290_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7293_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7294_));
OR2X2 OR2X2_3919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7295_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7296_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7297_));
OR2X2 OR2X2_392 ( .A(_abc_44694_new_n1793_), .B(_abc_44694_new_n1795_), .Y(_abc_44694_new_n1796_));
OR2X2 OR2X2_3920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7298_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7299_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7300_));
OR2X2 OR2X2_3921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7297_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7300_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7301_));
OR2X2 OR2X2_3922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7294_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7301_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7302_));
OR2X2 OR2X2_3923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7302_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7287_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7303_));
OR2X2 OR2X2_3924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7272_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7303_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_27_));
OR2X2 OR2X2_3925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7306_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7305_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7307_));
OR2X2 OR2X2_3926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7308_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7309_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7310_));
OR2X2 OR2X2_3927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7310_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7307_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7311_));
OR2X2 OR2X2_3928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7312_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7313_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7314_));
OR2X2 OR2X2_3929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7315_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7316_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7317_));
OR2X2 OR2X2_393 ( .A(_abc_44694_new_n1797_), .B(_abc_44694_new_n1278__bF_buf2), .Y(_abc_44694_new_n1798_));
OR2X2 OR2X2_3930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7317_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7314_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7318_));
OR2X2 OR2X2_3931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7318_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7311_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7319_));
OR2X2 OR2X2_3932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7321_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7322_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7323_));
OR2X2 OR2X2_3933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7323_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7320_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7324_));
OR2X2 OR2X2_3934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7325_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7326_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7327_));
OR2X2 OR2X2_3935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7329_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7328_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7330_));
OR2X2 OR2X2_3936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7327_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7330_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7331_));
OR2X2 OR2X2_3937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7331_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7324_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7332_));
OR2X2 OR2X2_3938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7332_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7319_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7333_));
OR2X2 OR2X2_3939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7335_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7334_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7336_));
OR2X2 OR2X2_394 ( .A(_abc_44694_new_n1799_), .B(_abc_44694_new_n1800_), .Y(_abc_44694_new_n1801_));
OR2X2 OR2X2_3940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7337_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7338_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7339_));
OR2X2 OR2X2_3941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7339_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7336_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7340_));
OR2X2 OR2X2_3942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7341_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7342_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7343_));
OR2X2 OR2X2_3943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7344_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7346_));
OR2X2 OR2X2_3944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7343_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7346_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7347_));
OR2X2 OR2X2_3945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7347_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7340_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7348_));
OR2X2 OR2X2_3946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7349_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7350_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7351_));
OR2X2 OR2X2_3947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7352_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7353_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7354_));
OR2X2 OR2X2_3948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7351_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7354_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7355_));
OR2X2 OR2X2_3949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7356_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7357_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7358_));
OR2X2 OR2X2_395 ( .A(_abc_44694_new_n1334__bF_buf2), .B(_abc_44694_new_n1801_), .Y(_abc_44694_new_n1802_));
OR2X2 OR2X2_3950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7359_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7360_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7361_));
OR2X2 OR2X2_3951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7358_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7361_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7362_));
OR2X2 OR2X2_3952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7355_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7362_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7363_));
OR2X2 OR2X2_3953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7363_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7348_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7364_));
OR2X2 OR2X2_3954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7333_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7364_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_28_));
OR2X2 OR2X2_3955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7366_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7368_));
OR2X2 OR2X2_3956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7369_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7371_));
OR2X2 OR2X2_3957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7371_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7372_));
OR2X2 OR2X2_3958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7373_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7374_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7375_));
OR2X2 OR2X2_3959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7376_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7377_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7378_));
OR2X2 OR2X2_396 ( .A(_abc_44694_new_n1804_), .B(_abc_44694_new_n1772_), .Y(_abc_44694_new_n1805_));
OR2X2 OR2X2_3960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7378_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7375_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7379_));
OR2X2 OR2X2_3961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7379_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7372_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7380_));
OR2X2 OR2X2_3962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7382_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7383_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7384_));
OR2X2 OR2X2_3963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7384_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7381_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7385_));
OR2X2 OR2X2_3964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7386_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7387_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7388_));
OR2X2 OR2X2_3965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7390_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7389_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7391_));
OR2X2 OR2X2_3966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7388_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7391_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7392_));
OR2X2 OR2X2_3967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7392_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7385_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7393_));
OR2X2 OR2X2_3968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7393_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7380_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7394_));
OR2X2 OR2X2_3969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7396_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7395_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7397_));
OR2X2 OR2X2_397 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_12_), .Y(_abc_44694_new_n1806_));
OR2X2 OR2X2_3970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7398_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7399_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7400_));
OR2X2 OR2X2_3971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7400_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7397_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7401_));
OR2X2 OR2X2_3972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7402_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7403_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7404_));
OR2X2 OR2X2_3973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7405_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7406_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7407_));
OR2X2 OR2X2_3974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7404_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7407_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7408_));
OR2X2 OR2X2_3975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7408_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7401_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7409_));
OR2X2 OR2X2_3976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7410_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7411_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7412_));
OR2X2 OR2X2_3977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7413_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7414_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7415_));
OR2X2 OR2X2_3978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7412_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7415_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7416_));
OR2X2 OR2X2_3979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7417_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7418_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7419_));
OR2X2 OR2X2_398 ( .A(_abc_44694_new_n1768_), .B(pc_q_13_), .Y(_abc_44694_new_n1809_));
OR2X2 OR2X2_3980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7420_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7421_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7422_));
OR2X2 OR2X2_3981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7419_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7422_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7423_));
OR2X2 OR2X2_3982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7416_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7423_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7424_));
OR2X2 OR2X2_3983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7424_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7409_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7425_));
OR2X2 OR2X2_3984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7394_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7425_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_29_));
OR2X2 OR2X2_3985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7428_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7427_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7429_));
OR2X2 OR2X2_3986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7430_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7431_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7432_));
OR2X2 OR2X2_3987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7432_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7429_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7433_));
OR2X2 OR2X2_3988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7434_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7436_));
OR2X2 OR2X2_3989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7437_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7438_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7439_));
OR2X2 OR2X2_399 ( .A(_abc_44694_new_n1812_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n1813_));
OR2X2 OR2X2_3990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7439_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7436_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7440_));
OR2X2 OR2X2_3991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7440_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7433_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7441_));
OR2X2 OR2X2_3992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7443_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7444_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7445_));
OR2X2 OR2X2_3993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7445_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7442_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7446_));
OR2X2 OR2X2_3994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7447_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7448_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7449_));
OR2X2 OR2X2_3995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7451_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7450_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7452_));
OR2X2 OR2X2_3996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7449_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7452_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7453_));
OR2X2 OR2X2_3997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7453_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7446_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7454_));
OR2X2 OR2X2_3998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7454_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7455_));
OR2X2 OR2X2_3999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7457_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7456_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7458_));
OR2X2 OR2X2_4 ( .A(state_q_4_), .B(state_q_0_), .Y(_abc_44694_new_n661_));
OR2X2 OR2X2_40 ( .A(_abc_44694_new_n751_), .B(_abc_44694_new_n759_), .Y(_abc_44694_new_n760_));
OR2X2 OR2X2_400 ( .A(_abc_44694_new_n1812_), .B(_abc_44694_new_n1399__bF_buf2), .Y(_abc_44694_new_n1815_));
OR2X2 OR2X2_4000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7459_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7460_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7461_));
OR2X2 OR2X2_4001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7461_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7458_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7462_));
OR2X2 OR2X2_4002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7463_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7464_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7465_));
OR2X2 OR2X2_4003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7466_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7467_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7468_));
OR2X2 OR2X2_4004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7465_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7469_));
OR2X2 OR2X2_4005 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7469_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7462_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7470_));
OR2X2 OR2X2_4006 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7472_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7473_));
OR2X2 OR2X2_4007 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7474_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7475_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7476_));
OR2X2 OR2X2_4008 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7473_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7476_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7477_));
OR2X2 OR2X2_4009 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7478_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7479_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7480_));
OR2X2 OR2X2_401 ( .A(pc_q_13_), .B(REGFILE_SIM_reg_bank_rb_i_0_), .Y(_abc_44694_new_n1817_));
OR2X2 OR2X2_4010 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7481_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7482_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7483_));
OR2X2 OR2X2_4011 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7480_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7483_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7484_));
OR2X2 OR2X2_4012 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7477_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7484_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7485_));
OR2X2 OR2X2_4013 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7485_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7470_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7486_));
OR2X2 OR2X2_4014 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7455_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7486_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_30_));
OR2X2 OR2X2_4015 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7489_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7488_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7490_));
OR2X2 OR2X2_4016 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7491_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7492_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7493_));
OR2X2 OR2X2_4017 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7493_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7490_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7494_));
OR2X2 OR2X2_4018 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7496_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7497_));
OR2X2 OR2X2_4019 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7498_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7499_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7500_));
OR2X2 OR2X2_402 ( .A(_abc_44694_new_n1820_), .B(_abc_44694_new_n1784_), .Y(_abc_44694_new_n1821_));
OR2X2 OR2X2_4020 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7500_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7497_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7501_));
OR2X2 OR2X2_4021 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7501_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7494_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7502_));
OR2X2 OR2X2_4022 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7504_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7505_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7506_));
OR2X2 OR2X2_4023 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7506_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7503_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7507_));
OR2X2 OR2X2_4024 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7508_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7509_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7510_));
OR2X2 OR2X2_4025 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7512_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7511_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7513_));
OR2X2 OR2X2_4026 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7510_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7513_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7514_));
OR2X2 OR2X2_4027 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7514_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7507_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7515_));
OR2X2 OR2X2_4028 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7502_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7516_));
OR2X2 OR2X2_4029 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7518_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7519_));
OR2X2 OR2X2_403 ( .A(_abc_44694_new_n1788_), .B(_abc_44694_new_n1821_), .Y(_abc_44694_new_n1822_));
OR2X2 OR2X2_4030 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7520_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7521_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7522_));
OR2X2 OR2X2_4031 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7522_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7523_));
OR2X2 OR2X2_4032 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7524_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7525_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7526_));
OR2X2 OR2X2_4033 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7527_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7528_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7529_));
OR2X2 OR2X2_4034 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7526_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7529_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7530_));
OR2X2 OR2X2_4035 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7530_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7523_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7531_));
OR2X2 OR2X2_4036 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7532_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7533_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7534_));
OR2X2 OR2X2_4037 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7535_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7536_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7537_));
OR2X2 OR2X2_4038 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7534_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7537_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7538_));
OR2X2 OR2X2_4039 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7539_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7540_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7541_));
OR2X2 OR2X2_404 ( .A(_abc_44694_new_n1830_), .B(_abc_44694_new_n1816_), .Y(_abc_44694_new_n1831_));
OR2X2 OR2X2_4040 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7542_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7544_));
OR2X2 OR2X2_4041 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7541_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7544_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7545_));
OR2X2 OR2X2_4042 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7538_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7545_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7546_));
OR2X2 OR2X2_4043 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7546_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7531_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7547_));
OR2X2 OR2X2_4044 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7516_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7547_), .Y(REGFILE_SIM_reg_bank_reg_rb_o_31_));
OR2X2 OR2X2_4045 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7559_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7560_));
OR2X2 OR2X2_4046 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7565_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7569_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7570_));
OR2X2 OR2X2_4047 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7570_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7560_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7571_));
OR2X2 OR2X2_4048 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7576_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7579_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7580_));
OR2X2 OR2X2_4049 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7583_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7586_));
OR2X2 OR2X2_405 ( .A(_abc_44694_new_n1400__bF_buf3), .B(_abc_44694_new_n1833_), .Y(_abc_44694_new_n1834_));
OR2X2 OR2X2_4050 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7586_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7580_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7587_));
OR2X2 OR2X2_4051 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7587_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7571_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7588_));
OR2X2 OR2X2_4052 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7596_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7599_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7600_));
OR2X2 OR2X2_4053 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7600_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7593_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7601_));
OR2X2 OR2X2_4054 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7605_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7607_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7608_));
OR2X2 OR2X2_4055 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7614_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7611_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7615_));
OR2X2 OR2X2_4056 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7608_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7615_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7616_));
OR2X2 OR2X2_4057 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7616_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7601_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7617_));
OR2X2 OR2X2_4058 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7617_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7588_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7618_));
OR2X2 OR2X2_4059 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7622_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7620_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7623_));
OR2X2 OR2X2_406 ( .A(_abc_44694_new_n1832_), .B(_abc_44694_new_n1834_), .Y(_abc_44694_new_n1835_));
OR2X2 OR2X2_4060 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7626_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7629_));
OR2X2 OR2X2_4061 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7629_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7630_));
OR2X2 OR2X2_4062 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7632_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7634_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7635_));
OR2X2 OR2X2_4063 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7637_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7639_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7640_));
OR2X2 OR2X2_4064 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7635_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7641_));
OR2X2 OR2X2_4065 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7641_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7630_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7642_));
OR2X2 OR2X2_4066 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7644_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7647_));
OR2X2 OR2X2_4067 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7649_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7651_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7652_));
OR2X2 OR2X2_4068 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7647_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7652_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7653_));
OR2X2 OR2X2_4069 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7655_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7657_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7658_));
OR2X2 OR2X2_407 ( .A(_abc_44694_new_n1836_), .B(_abc_44694_new_n1278__bF_buf1), .Y(_abc_44694_new_n1837_));
OR2X2 OR2X2_4070 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7660_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7662_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7663_));
OR2X2 OR2X2_4071 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7658_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7663_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7664_));
OR2X2 OR2X2_4072 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7653_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7664_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7665_));
OR2X2 OR2X2_4073 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7665_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7642_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7666_));
OR2X2 OR2X2_4074 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7618_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7666_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_0_));
OR2X2 OR2X2_4075 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7669_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7668_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7670_));
OR2X2 OR2X2_4076 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7671_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7672_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7673_));
OR2X2 OR2X2_4077 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7673_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7670_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7674_));
OR2X2 OR2X2_4078 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7675_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7676_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7677_));
OR2X2 OR2X2_4079 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7678_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7679_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7680_));
OR2X2 OR2X2_408 ( .A(_abc_44694_new_n1838_), .B(_abc_44694_new_n1839_), .Y(_abc_44694_new_n1840_));
OR2X2 OR2X2_4080 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7680_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7677_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7681_));
OR2X2 OR2X2_4081 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7681_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7674_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7682_));
OR2X2 OR2X2_4082 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7684_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7685_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7686_));
OR2X2 OR2X2_4083 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7686_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7683_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7687_));
OR2X2 OR2X2_4084 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7688_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7689_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7690_));
OR2X2 OR2X2_4085 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7692_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7691_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7693_));
OR2X2 OR2X2_4086 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7690_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7693_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7694_));
OR2X2 OR2X2_4087 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7694_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7687_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7695_));
OR2X2 OR2X2_4088 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7695_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7682_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7696_));
OR2X2 OR2X2_4089 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7698_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7697_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7699_));
OR2X2 OR2X2_409 ( .A(_abc_44694_new_n1334__bF_buf1), .B(_abc_44694_new_n1840_), .Y(_abc_44694_new_n1841_));
OR2X2 OR2X2_4090 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7700_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7701_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7702_));
OR2X2 OR2X2_4091 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7702_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7703_));
OR2X2 OR2X2_4092 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7704_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7705_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7706_));
OR2X2 OR2X2_4093 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7707_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7708_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7709_));
OR2X2 OR2X2_4094 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7706_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7709_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7710_));
OR2X2 OR2X2_4095 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7710_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7703_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7711_));
OR2X2 OR2X2_4096 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7712_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7713_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7714_));
OR2X2 OR2X2_4097 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7715_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7716_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7717_));
OR2X2 OR2X2_4098 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7714_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7717_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7718_));
OR2X2 OR2X2_4099 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7719_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7720_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7721_));
OR2X2 OR2X2_41 ( .A(_abc_44694_new_n761_), .B(_abc_44694_new_n747_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_4_));
OR2X2 OR2X2_410 ( .A(_abc_44694_new_n1843_), .B(_abc_44694_new_n1814_), .Y(_abc_44694_new_n1844_));
OR2X2 OR2X2_4100 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7722_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7723_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7724_));
OR2X2 OR2X2_4101 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7721_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7724_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7725_));
OR2X2 OR2X2_4102 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7718_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7725_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7726_));
OR2X2 OR2X2_4103 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7726_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7711_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7727_));
OR2X2 OR2X2_4104 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7696_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7727_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_1_));
OR2X2 OR2X2_4105 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7730_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7729_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7731_));
OR2X2 OR2X2_4106 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7732_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7733_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7734_));
OR2X2 OR2X2_4107 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7734_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7731_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7735_));
OR2X2 OR2X2_4108 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7736_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7737_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7738_));
OR2X2 OR2X2_4109 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7739_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7740_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7741_));
OR2X2 OR2X2_411 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_13_), .Y(_abc_44694_new_n1845_));
OR2X2 OR2X2_4110 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7741_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7738_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7742_));
OR2X2 OR2X2_4111 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7742_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7735_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7743_));
OR2X2 OR2X2_4112 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7745_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7746_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7747_));
OR2X2 OR2X2_4113 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7747_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7744_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7748_));
OR2X2 OR2X2_4114 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7749_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7750_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7751_));
OR2X2 OR2X2_4115 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7753_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7752_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7754_));
OR2X2 OR2X2_4116 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7751_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7754_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7755_));
OR2X2 OR2X2_4117 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7755_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7748_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7756_));
OR2X2 OR2X2_4118 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7756_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7743_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7757_));
OR2X2 OR2X2_4119 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7759_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7758_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7760_));
OR2X2 OR2X2_412 ( .A(_abc_44694_new_n1810_), .B(pc_q_14_), .Y(_abc_44694_new_n1848_));
OR2X2 OR2X2_4120 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7761_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7762_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7763_));
OR2X2 OR2X2_4121 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7763_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7760_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7764_));
OR2X2 OR2X2_4122 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7765_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7766_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7767_));
OR2X2 OR2X2_4123 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7768_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7769_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7770_));
OR2X2 OR2X2_4124 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7767_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7770_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7771_));
OR2X2 OR2X2_4125 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7771_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7764_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7772_));
OR2X2 OR2X2_4126 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7773_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7774_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7775_));
OR2X2 OR2X2_4127 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7776_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7777_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7778_));
OR2X2 OR2X2_4128 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7775_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7778_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7779_));
OR2X2 OR2X2_4129 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7780_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7781_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7782_));
OR2X2 OR2X2_413 ( .A(_abc_44694_new_n1851_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n1852_));
OR2X2 OR2X2_4130 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7783_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7784_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7785_));
OR2X2 OR2X2_4131 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7782_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7785_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7786_));
OR2X2 OR2X2_4132 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7779_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7786_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7787_));
OR2X2 OR2X2_4133 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7787_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7772_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7788_));
OR2X2 OR2X2_4134 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7757_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7788_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_2_));
OR2X2 OR2X2_4135 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7791_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7790_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7792_));
OR2X2 OR2X2_4136 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7793_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7794_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7795_));
OR2X2 OR2X2_4137 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7795_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7792_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7796_));
OR2X2 OR2X2_4138 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7797_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7798_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7799_));
OR2X2 OR2X2_4139 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7800_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7801_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7802_));
OR2X2 OR2X2_414 ( .A(_abc_44694_new_n1851_), .B(_abc_44694_new_n1399__bF_buf1), .Y(_abc_44694_new_n1854_));
OR2X2 OR2X2_4140 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7802_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7799_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7803_));
OR2X2 OR2X2_4141 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7803_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7796_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7804_));
OR2X2 OR2X2_4142 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7806_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7807_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7808_));
OR2X2 OR2X2_4143 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7808_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7805_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7809_));
OR2X2 OR2X2_4144 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7810_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7811_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7812_));
OR2X2 OR2X2_4145 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7814_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7813_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7815_));
OR2X2 OR2X2_4146 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7812_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7816_));
OR2X2 OR2X2_4147 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7816_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7809_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7817_));
OR2X2 OR2X2_4148 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7817_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7804_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7818_));
OR2X2 OR2X2_4149 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7820_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7819_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7821_));
OR2X2 OR2X2_415 ( .A(pc_q_14_), .B(REGFILE_SIM_reg_bank_rb_i_1_), .Y(_abc_44694_new_n1859_));
OR2X2 OR2X2_4150 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7822_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7823_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7824_));
OR2X2 OR2X2_4151 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7824_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7821_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7825_));
OR2X2 OR2X2_4152 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7826_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7827_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7828_));
OR2X2 OR2X2_4153 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7829_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7830_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7831_));
OR2X2 OR2X2_4154 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7828_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7831_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7832_));
OR2X2 OR2X2_4155 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7832_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7825_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7833_));
OR2X2 OR2X2_4156 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7834_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7835_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7836_));
OR2X2 OR2X2_4157 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7837_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7838_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7839_));
OR2X2 OR2X2_4158 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7836_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7839_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7840_));
OR2X2 OR2X2_4159 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7841_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7842_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7843_));
OR2X2 OR2X2_416 ( .A(_abc_44694_new_n1858_), .B(_abc_44694_new_n1862_), .Y(_abc_44694_new_n1865_));
OR2X2 OR2X2_4160 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7844_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7845_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7846_));
OR2X2 OR2X2_4161 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7843_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7846_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7847_));
OR2X2 OR2X2_4162 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7840_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7847_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7848_));
OR2X2 OR2X2_4163 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7848_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7833_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7849_));
OR2X2 OR2X2_4164 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7818_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7849_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_3_));
OR2X2 OR2X2_4165 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7852_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7851_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7853_));
OR2X2 OR2X2_4166 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7854_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7855_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7856_));
OR2X2 OR2X2_4167 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7856_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7853_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7857_));
OR2X2 OR2X2_4168 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7858_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7859_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7860_));
OR2X2 OR2X2_4169 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7861_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7862_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7863_));
OR2X2 OR2X2_417 ( .A(_abc_44694_new_n1867_), .B(_abc_44694_new_n1855_), .Y(_abc_44694_new_n1868_));
OR2X2 OR2X2_4170 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7863_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7860_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7864_));
OR2X2 OR2X2_4171 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7864_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7857_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7865_));
OR2X2 OR2X2_4172 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7867_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7868_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7869_));
OR2X2 OR2X2_4173 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7869_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7866_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7870_));
OR2X2 OR2X2_4174 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7871_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7872_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7873_));
OR2X2 OR2X2_4175 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7875_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7874_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7876_));
OR2X2 OR2X2_4176 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7873_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7876_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7877_));
OR2X2 OR2X2_4177 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7877_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7870_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7878_));
OR2X2 OR2X2_4178 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7878_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7865_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7879_));
OR2X2 OR2X2_4179 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7881_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7880_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7882_));
OR2X2 OR2X2_418 ( .A(_abc_44694_new_n1400__bF_buf2), .B(_abc_44694_new_n1870_), .Y(_abc_44694_new_n1871_));
OR2X2 OR2X2_4180 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7883_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7884_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7885_));
OR2X2 OR2X2_4181 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7885_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7882_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7886_));
OR2X2 OR2X2_4182 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7887_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7888_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7889_));
OR2X2 OR2X2_4183 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7890_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7891_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7892_));
OR2X2 OR2X2_4184 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7889_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7892_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7893_));
OR2X2 OR2X2_4185 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7893_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7886_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7894_));
OR2X2 OR2X2_4186 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7895_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7896_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7897_));
OR2X2 OR2X2_4187 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7898_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7899_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7900_));
OR2X2 OR2X2_4188 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7897_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7900_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7901_));
OR2X2 OR2X2_4189 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7902_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7903_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7904_));
OR2X2 OR2X2_419 ( .A(_abc_44694_new_n1869_), .B(_abc_44694_new_n1871_), .Y(_abc_44694_new_n1872_));
OR2X2 OR2X2_4190 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7905_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7906_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7907_));
OR2X2 OR2X2_4191 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7904_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7907_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7908_));
OR2X2 OR2X2_4192 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7901_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7908_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7909_));
OR2X2 OR2X2_4193 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7909_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7894_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7910_));
OR2X2 OR2X2_4194 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7879_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7910_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_4_));
OR2X2 OR2X2_4195 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7913_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7912_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7914_));
OR2X2 OR2X2_4196 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7915_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7916_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7917_));
OR2X2 OR2X2_4197 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7917_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7914_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7918_));
OR2X2 OR2X2_4198 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7919_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7920_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7921_));
OR2X2 OR2X2_4199 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7922_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7923_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7924_));
OR2X2 OR2X2_42 ( .A(_abc_44694_new_n764_), .B(_abc_44694_new_n765_), .Y(_abc_44694_new_n766_));
OR2X2 OR2X2_420 ( .A(_abc_44694_new_n1873_), .B(_abc_44694_new_n1278__bF_buf0), .Y(_abc_44694_new_n1874_));
OR2X2 OR2X2_4200 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7924_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7921_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7925_));
OR2X2 OR2X2_4201 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7925_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7918_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7926_));
OR2X2 OR2X2_4202 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7928_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7929_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7930_));
OR2X2 OR2X2_4203 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7930_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7927_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7931_));
OR2X2 OR2X2_4204 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7932_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7933_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7934_));
OR2X2 OR2X2_4205 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7936_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7935_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7937_));
OR2X2 OR2X2_4206 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7934_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7937_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7938_));
OR2X2 OR2X2_4207 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7938_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7931_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7939_));
OR2X2 OR2X2_4208 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7939_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7926_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7940_));
OR2X2 OR2X2_4209 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7942_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7941_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7943_));
OR2X2 OR2X2_421 ( .A(_abc_44694_new_n1875_), .B(_abc_44694_new_n1876_), .Y(_abc_44694_new_n1877_));
OR2X2 OR2X2_4210 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7944_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7945_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7946_));
OR2X2 OR2X2_4211 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7946_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7943_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7947_));
OR2X2 OR2X2_4212 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7948_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7949_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7950_));
OR2X2 OR2X2_4213 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7951_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7952_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7953_));
OR2X2 OR2X2_4214 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7950_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7953_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7954_));
OR2X2 OR2X2_4215 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7954_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7947_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7955_));
OR2X2 OR2X2_4216 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7956_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7957_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7958_));
OR2X2 OR2X2_4217 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7959_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7961_));
OR2X2 OR2X2_4218 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7958_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7961_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7962_));
OR2X2 OR2X2_4219 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7963_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7964_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7965_));
OR2X2 OR2X2_422 ( .A(_abc_44694_new_n1334__bF_buf0), .B(_abc_44694_new_n1877_), .Y(_abc_44694_new_n1878_));
OR2X2 OR2X2_4220 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7966_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7967_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7968_));
OR2X2 OR2X2_4221 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7965_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7968_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7969_));
OR2X2 OR2X2_4222 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7962_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7969_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7970_));
OR2X2 OR2X2_4223 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7970_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7955_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7971_));
OR2X2 OR2X2_4224 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7940_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7971_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_5_));
OR2X2 OR2X2_4225 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7974_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7973_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7975_));
OR2X2 OR2X2_4226 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7976_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7977_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7978_));
OR2X2 OR2X2_4227 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7978_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7975_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7979_));
OR2X2 OR2X2_4228 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7980_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7981_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7982_));
OR2X2 OR2X2_4229 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7983_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7984_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7985_));
OR2X2 OR2X2_423 ( .A(_abc_44694_new_n1880_), .B(_abc_44694_new_n1853_), .Y(_abc_44694_new_n1881_));
OR2X2 OR2X2_4230 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7985_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7982_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7986_));
OR2X2 OR2X2_4231 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7986_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7979_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7987_));
OR2X2 OR2X2_4232 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7989_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7990_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7991_));
OR2X2 OR2X2_4233 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7991_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7988_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7992_));
OR2X2 OR2X2_4234 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7993_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7994_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7995_));
OR2X2 OR2X2_4235 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7997_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7996_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7998_));
OR2X2 OR2X2_4236 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7995_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7998_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n7999_));
OR2X2 OR2X2_4237 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n7999_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7992_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8000_));
OR2X2 OR2X2_4238 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8000_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n7987_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8001_));
OR2X2 OR2X2_4239 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8003_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8002_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8004_));
OR2X2 OR2X2_424 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_14_), .Y(_abc_44694_new_n1882_));
OR2X2 OR2X2_4240 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8005_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8006_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8007_));
OR2X2 OR2X2_4241 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8007_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8004_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8008_));
OR2X2 OR2X2_4242 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8009_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8010_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8011_));
OR2X2 OR2X2_4243 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8012_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8013_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8014_));
OR2X2 OR2X2_4244 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8011_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8014_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8015_));
OR2X2 OR2X2_4245 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8015_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8008_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8016_));
OR2X2 OR2X2_4246 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8017_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8018_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8019_));
OR2X2 OR2X2_4247 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8020_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8021_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8022_));
OR2X2 OR2X2_4248 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8019_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8022_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8023_));
OR2X2 OR2X2_4249 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8024_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8025_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8026_));
OR2X2 OR2X2_425 ( .A(_abc_44694_new_n1849_), .B(pc_q_15_), .Y(_abc_44694_new_n1885_));
OR2X2 OR2X2_4250 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8027_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8028_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8029_));
OR2X2 OR2X2_4251 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8026_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8029_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8030_));
OR2X2 OR2X2_4252 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8023_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8030_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8031_));
OR2X2 OR2X2_4253 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8031_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8016_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8032_));
OR2X2 OR2X2_4254 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8001_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8032_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_6_));
OR2X2 OR2X2_4255 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8035_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8034_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8036_));
OR2X2 OR2X2_4256 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8037_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8038_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8039_));
OR2X2 OR2X2_4257 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8039_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8036_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8040_));
OR2X2 OR2X2_4258 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8041_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8042_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8043_));
OR2X2 OR2X2_4259 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8044_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8045_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8046_));
OR2X2 OR2X2_426 ( .A(_abc_44694_new_n1888_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n1889_));
OR2X2 OR2X2_4260 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8046_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8043_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8047_));
OR2X2 OR2X2_4261 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8047_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8040_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8048_));
OR2X2 OR2X2_4262 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8050_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8051_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8052_));
OR2X2 OR2X2_4263 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8052_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8049_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8053_));
OR2X2 OR2X2_4264 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8055_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8056_));
OR2X2 OR2X2_4265 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8058_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8057_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8059_));
OR2X2 OR2X2_4266 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8056_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8060_));
OR2X2 OR2X2_4267 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8060_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8053_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8061_));
OR2X2 OR2X2_4268 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8061_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8048_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8062_));
OR2X2 OR2X2_4269 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8064_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8063_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8065_));
OR2X2 OR2X2_427 ( .A(_abc_44694_new_n1888_), .B(_abc_44694_new_n1399__bF_buf0), .Y(_abc_44694_new_n1891_));
OR2X2 OR2X2_4270 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8066_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8067_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8068_));
OR2X2 OR2X2_4271 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8068_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8065_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8069_));
OR2X2 OR2X2_4272 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8070_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8071_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8072_));
OR2X2 OR2X2_4273 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8073_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8074_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8075_));
OR2X2 OR2X2_4274 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8072_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8075_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8076_));
OR2X2 OR2X2_4275 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8076_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8069_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8077_));
OR2X2 OR2X2_4276 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8078_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8079_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8080_));
OR2X2 OR2X2_4277 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8081_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8082_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8083_));
OR2X2 OR2X2_4278 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8080_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8083_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8084_));
OR2X2 OR2X2_4279 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8085_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8086_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8087_));
OR2X2 OR2X2_428 ( .A(pc_q_15_), .B(REGFILE_SIM_reg_bank_rb_i_2_), .Y(_abc_44694_new_n1895_));
OR2X2 OR2X2_4280 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8088_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8089_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8090_));
OR2X2 OR2X2_4281 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8087_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8090_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8091_));
OR2X2 OR2X2_4282 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8084_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8091_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8092_));
OR2X2 OR2X2_4283 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8092_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8077_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8093_));
OR2X2 OR2X2_4284 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8062_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8093_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_7_));
OR2X2 OR2X2_4285 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8096_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8095_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8097_));
OR2X2 OR2X2_4286 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8098_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8099_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8100_));
OR2X2 OR2X2_4287 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8100_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8097_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8101_));
OR2X2 OR2X2_4288 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8102_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8103_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8104_));
OR2X2 OR2X2_4289 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8105_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8106_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8107_));
OR2X2 OR2X2_429 ( .A(_abc_44694_new_n1894_), .B(_abc_44694_new_n1898_), .Y(_abc_44694_new_n1899_));
OR2X2 OR2X2_4290 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8107_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8104_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8108_));
OR2X2 OR2X2_4291 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8108_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8101_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8109_));
OR2X2 OR2X2_4292 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8111_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8112_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8113_));
OR2X2 OR2X2_4293 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8113_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8110_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8114_));
OR2X2 OR2X2_4294 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8115_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8117_));
OR2X2 OR2X2_4295 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8119_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8118_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8120_));
OR2X2 OR2X2_4296 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8117_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8121_));
OR2X2 OR2X2_4297 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8121_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8114_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8122_));
OR2X2 OR2X2_4298 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8122_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8109_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8123_));
OR2X2 OR2X2_4299 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8125_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8124_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8126_));
OR2X2 OR2X2_43 ( .A(_abc_44694_new_n768_), .B(_abc_44694_new_n769_), .Y(_abc_44694_new_n770_));
OR2X2 OR2X2_430 ( .A(_abc_44694_new_n1893_), .B(_abc_44694_new_n1900_), .Y(_abc_44694_new_n1901_));
OR2X2 OR2X2_4300 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8127_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8128_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8129_));
OR2X2 OR2X2_4301 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8129_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8126_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8130_));
OR2X2 OR2X2_4302 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8131_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8132_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8133_));
OR2X2 OR2X2_4303 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8134_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8135_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8136_));
OR2X2 OR2X2_4304 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8133_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8136_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8137_));
OR2X2 OR2X2_4305 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8137_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8130_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8138_));
OR2X2 OR2X2_4306 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8139_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8141_));
OR2X2 OR2X2_4307 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8142_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8143_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8144_));
OR2X2 OR2X2_4308 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8141_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8144_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8145_));
OR2X2 OR2X2_4309 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8146_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8147_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8148_));
OR2X2 OR2X2_431 ( .A(_abc_44694_new_n1903_), .B(_abc_44694_new_n1892_), .Y(_abc_44694_new_n1904_));
OR2X2 OR2X2_4310 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8149_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8150_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8151_));
OR2X2 OR2X2_4311 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8148_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8151_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8152_));
OR2X2 OR2X2_4312 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8145_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8152_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8153_));
OR2X2 OR2X2_4313 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8153_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8138_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8154_));
OR2X2 OR2X2_4314 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8123_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8154_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_8_));
OR2X2 OR2X2_4315 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8157_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8156_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8158_));
OR2X2 OR2X2_4316 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8159_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8160_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8161_));
OR2X2 OR2X2_4317 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8161_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8158_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8162_));
OR2X2 OR2X2_4318 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8163_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8164_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8165_));
OR2X2 OR2X2_4319 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8166_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8167_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8168_));
OR2X2 OR2X2_432 ( .A(_abc_44694_new_n1400__bF_buf1), .B(_abc_44694_new_n1906_), .Y(_abc_44694_new_n1907_));
OR2X2 OR2X2_4320 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8168_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8169_));
OR2X2 OR2X2_4321 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8169_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8162_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8170_));
OR2X2 OR2X2_4322 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8172_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8173_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8174_));
OR2X2 OR2X2_4323 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8174_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8171_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8175_));
OR2X2 OR2X2_4324 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8176_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8177_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8178_));
OR2X2 OR2X2_4325 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8180_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8179_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8181_));
OR2X2 OR2X2_4326 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8178_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8181_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8182_));
OR2X2 OR2X2_4327 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8182_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8183_));
OR2X2 OR2X2_4328 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8183_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8170_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8184_));
OR2X2 OR2X2_4329 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8186_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8185_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8187_));
OR2X2 OR2X2_433 ( .A(_abc_44694_new_n1905_), .B(_abc_44694_new_n1907_), .Y(_abc_44694_new_n1908_));
OR2X2 OR2X2_4330 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8188_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8189_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8190_));
OR2X2 OR2X2_4331 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8190_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8187_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8191_));
OR2X2 OR2X2_4332 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8192_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8193_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8194_));
OR2X2 OR2X2_4333 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8195_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8196_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8197_));
OR2X2 OR2X2_4334 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8194_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8197_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8198_));
OR2X2 OR2X2_4335 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8198_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8191_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8199_));
OR2X2 OR2X2_4336 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8200_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8201_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8202_));
OR2X2 OR2X2_4337 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8203_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8204_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8205_));
OR2X2 OR2X2_4338 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8202_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8205_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8206_));
OR2X2 OR2X2_4339 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8207_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8208_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8209_));
OR2X2 OR2X2_434 ( .A(_abc_44694_new_n1909_), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n1910_));
OR2X2 OR2X2_4340 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8210_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8211_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8212_));
OR2X2 OR2X2_4341 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8209_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8212_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8213_));
OR2X2 OR2X2_4342 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8206_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8213_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8214_));
OR2X2 OR2X2_4343 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8214_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8199_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8215_));
OR2X2 OR2X2_4344 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8184_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8215_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_9_));
OR2X2 OR2X2_4345 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8218_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8217_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8219_));
OR2X2 OR2X2_4346 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8220_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8221_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8222_));
OR2X2 OR2X2_4347 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8222_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8219_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8223_));
OR2X2 OR2X2_4348 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8224_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8225_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8226_));
OR2X2 OR2X2_4349 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8228_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8229_));
OR2X2 OR2X2_435 ( .A(_abc_44694_new_n1911_), .B(_abc_44694_new_n1912_), .Y(_abc_44694_new_n1913_));
OR2X2 OR2X2_4350 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8229_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8226_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8230_));
OR2X2 OR2X2_4351 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8230_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8223_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8231_));
OR2X2 OR2X2_4352 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8233_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8234_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8235_));
OR2X2 OR2X2_4353 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8235_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8232_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8236_));
OR2X2 OR2X2_4354 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8237_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8238_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8239_));
OR2X2 OR2X2_4355 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8241_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8240_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8242_));
OR2X2 OR2X2_4356 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8239_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8242_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8243_));
OR2X2 OR2X2_4357 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8243_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8236_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8244_));
OR2X2 OR2X2_4358 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8244_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8231_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8245_));
OR2X2 OR2X2_4359 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8247_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8246_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8248_));
OR2X2 OR2X2_436 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n1913_), .Y(_abc_44694_new_n1914_));
OR2X2 OR2X2_4360 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8249_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8251_));
OR2X2 OR2X2_4361 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8251_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8248_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8252_));
OR2X2 OR2X2_4362 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8253_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8254_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8255_));
OR2X2 OR2X2_4363 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8256_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8257_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8258_));
OR2X2 OR2X2_4364 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8255_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8258_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8259_));
OR2X2 OR2X2_4365 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8259_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8252_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8260_));
OR2X2 OR2X2_4366 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8261_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8262_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8263_));
OR2X2 OR2X2_4367 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8264_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8265_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8266_));
OR2X2 OR2X2_4368 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8263_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8266_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8267_));
OR2X2 OR2X2_4369 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8268_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8270_));
OR2X2 OR2X2_437 ( .A(_abc_44694_new_n1916_), .B(_abc_44694_new_n1890_), .Y(_abc_44694_new_n1917_));
OR2X2 OR2X2_4370 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8271_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8272_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8273_));
OR2X2 OR2X2_4371 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8270_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8273_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8274_));
OR2X2 OR2X2_4372 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8267_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8274_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8275_));
OR2X2 OR2X2_4373 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8275_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8276_));
OR2X2 OR2X2_4374 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8245_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8276_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_10_));
OR2X2 OR2X2_4375 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8279_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8278_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8280_));
OR2X2 OR2X2_4376 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8281_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8282_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8283_));
OR2X2 OR2X2_4377 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8283_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8280_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8284_));
OR2X2 OR2X2_4378 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8285_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8286_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8287_));
OR2X2 OR2X2_4379 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8288_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8289_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8290_));
OR2X2 OR2X2_438 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_15_), .Y(_abc_44694_new_n1918_));
OR2X2 OR2X2_4380 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8290_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8287_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8291_));
OR2X2 OR2X2_4381 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8291_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8284_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8292_));
OR2X2 OR2X2_4382 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8294_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8295_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8296_));
OR2X2 OR2X2_4383 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8296_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8293_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8297_));
OR2X2 OR2X2_4384 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8298_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8299_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8300_));
OR2X2 OR2X2_4385 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8302_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8301_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8303_));
OR2X2 OR2X2_4386 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8300_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8303_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8304_));
OR2X2 OR2X2_4387 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8304_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8297_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8305_));
OR2X2 OR2X2_4388 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8305_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8292_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8306_));
OR2X2 OR2X2_4389 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8308_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8307_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8309_));
OR2X2 OR2X2_439 ( .A(_abc_44694_new_n1886_), .B(pc_q_16_), .Y(_abc_44694_new_n1921_));
OR2X2 OR2X2_4390 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8310_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8311_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8312_));
OR2X2 OR2X2_4391 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8312_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8309_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8313_));
OR2X2 OR2X2_4392 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8314_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8315_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8316_));
OR2X2 OR2X2_4393 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8317_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8318_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8319_));
OR2X2 OR2X2_4394 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8316_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8319_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8320_));
OR2X2 OR2X2_4395 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8320_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8313_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8321_));
OR2X2 OR2X2_4396 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8322_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8323_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8324_));
OR2X2 OR2X2_4397 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8325_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8326_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8327_));
OR2X2 OR2X2_4398 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8324_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8327_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8328_));
OR2X2 OR2X2_4399 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8329_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8330_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8331_));
OR2X2 OR2X2_44 ( .A(_abc_44694_new_n771_), .B(_abc_44694_new_n772_), .Y(_abc_44694_new_n773_));
OR2X2 OR2X2_440 ( .A(_abc_44694_new_n1924_), .B(_abc_44694_new_n1210__bF_buf1), .Y(_abc_44694_new_n1925_));
OR2X2 OR2X2_4400 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8332_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8333_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8334_));
OR2X2 OR2X2_4401 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8331_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8334_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8335_));
OR2X2 OR2X2_4402 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8328_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8335_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8336_));
OR2X2 OR2X2_4403 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8336_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8321_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8337_));
OR2X2 OR2X2_4404 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8306_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8337_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_11_));
OR2X2 OR2X2_4405 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8340_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8339_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8341_));
OR2X2 OR2X2_4406 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8342_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8343_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8344_));
OR2X2 OR2X2_4407 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8344_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8341_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8345_));
OR2X2 OR2X2_4408 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8346_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8347_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8348_));
OR2X2 OR2X2_4409 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8349_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8350_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8351_));
OR2X2 OR2X2_441 ( .A(_abc_44694_new_n1924_), .B(_abc_44694_new_n1399__bF_buf4), .Y(_abc_44694_new_n1927_));
OR2X2 OR2X2_4410 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8351_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8348_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8352_));
OR2X2 OR2X2_4411 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8352_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8345_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8353_));
OR2X2 OR2X2_4412 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8355_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8356_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8357_));
OR2X2 OR2X2_4413 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8357_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8354_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8358_));
OR2X2 OR2X2_4414 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8359_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8360_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8361_));
OR2X2 OR2X2_4415 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8363_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8362_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8364_));
OR2X2 OR2X2_4416 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8361_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8364_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8365_));
OR2X2 OR2X2_4417 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8365_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8358_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8366_));
OR2X2 OR2X2_4418 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8366_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8353_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8367_));
OR2X2 OR2X2_4419 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8369_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8368_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8370_));
OR2X2 OR2X2_442 ( .A(_abc_44694_new_n1932_), .B(_abc_44694_new_n1896_), .Y(_abc_44694_new_n1933_));
OR2X2 OR2X2_4420 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8371_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8372_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8373_));
OR2X2 OR2X2_4421 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8373_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8374_));
OR2X2 OR2X2_4422 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8375_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8376_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8377_));
OR2X2 OR2X2_4423 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8378_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8379_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8380_));
OR2X2 OR2X2_4424 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8377_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8380_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8381_));
OR2X2 OR2X2_4425 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8381_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8374_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8382_));
OR2X2 OR2X2_4426 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8383_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8384_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8385_));
OR2X2 OR2X2_4427 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8386_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8387_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8388_));
OR2X2 OR2X2_4428 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8385_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8388_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8389_));
OR2X2 OR2X2_4429 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8390_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8391_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8392_));
OR2X2 OR2X2_443 ( .A(_abc_44694_new_n1935_), .B(_abc_44694_new_n1933_), .Y(_abc_44694_new_n1936_));
OR2X2 OR2X2_4430 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8393_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8394_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8395_));
OR2X2 OR2X2_4431 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8392_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8395_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8396_));
OR2X2 OR2X2_4432 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8389_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8396_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8397_));
OR2X2 OR2X2_4433 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8397_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8382_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8398_));
OR2X2 OR2X2_4434 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8367_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8398_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_12_));
OR2X2 OR2X2_4435 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8401_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8400_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8402_));
OR2X2 OR2X2_4436 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8403_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8404_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8405_));
OR2X2 OR2X2_4437 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8405_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8402_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8406_));
OR2X2 OR2X2_4438 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8407_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8408_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8409_));
OR2X2 OR2X2_4439 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8410_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8411_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8412_));
OR2X2 OR2X2_444 ( .A(_abc_44694_new_n1936_), .B(_abc_44694_new_n1931_), .Y(_abc_44694_new_n1937_));
OR2X2 OR2X2_4440 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8412_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8409_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8413_));
OR2X2 OR2X2_4441 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8413_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8406_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8414_));
OR2X2 OR2X2_4442 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8416_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8418_));
OR2X2 OR2X2_4443 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8418_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8415_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8419_));
OR2X2 OR2X2_4444 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8420_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8421_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8422_));
OR2X2 OR2X2_4445 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8424_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8423_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8425_));
OR2X2 OR2X2_4446 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8422_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8425_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8426_));
OR2X2 OR2X2_4447 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8426_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8427_));
OR2X2 OR2X2_4448 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8427_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8414_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8428_));
OR2X2 OR2X2_4449 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8430_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8429_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8431_));
OR2X2 OR2X2_445 ( .A(_abc_44694_new_n1939_), .B(_abc_44694_new_n1937_), .Y(_abc_44694_new_n1940_));
OR2X2 OR2X2_4450 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8432_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8433_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8434_));
OR2X2 OR2X2_4451 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8434_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8431_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8435_));
OR2X2 OR2X2_4452 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8436_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8437_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8438_));
OR2X2 OR2X2_4453 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8439_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8440_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8441_));
OR2X2 OR2X2_4454 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8438_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8442_));
OR2X2 OR2X2_4455 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8442_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8435_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8443_));
OR2X2 OR2X2_4456 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8444_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8445_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8446_));
OR2X2 OR2X2_4457 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8447_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8448_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8449_));
OR2X2 OR2X2_4458 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8446_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8449_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8450_));
OR2X2 OR2X2_4459 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8451_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8452_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8453_));
OR2X2 OR2X2_446 ( .A(pc_q_16_), .B(REGFILE_SIM_reg_bank_rb_i_3_), .Y(_abc_44694_new_n1941_));
OR2X2 OR2X2_4460 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8454_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8455_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8456_));
OR2X2 OR2X2_4461 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8453_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8456_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8457_));
OR2X2 OR2X2_4462 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8450_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8457_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8458_));
OR2X2 OR2X2_4463 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8458_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8459_));
OR2X2 OR2X2_4464 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8428_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8459_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_13_));
OR2X2 OR2X2_4465 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8462_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8461_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8463_));
OR2X2 OR2X2_4466 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8464_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8465_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8466_));
OR2X2 OR2X2_4467 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8466_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8463_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8467_));
OR2X2 OR2X2_4468 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8468_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8469_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8470_));
OR2X2 OR2X2_4469 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8472_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8473_));
OR2X2 OR2X2_447 ( .A(_abc_44694_new_n1940_), .B(_abc_44694_new_n1944_), .Y(_abc_44694_new_n1945_));
OR2X2 OR2X2_4470 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8473_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8470_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8474_));
OR2X2 OR2X2_4471 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8474_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8467_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8475_));
OR2X2 OR2X2_4472 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8477_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8478_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8479_));
OR2X2 OR2X2_4473 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8479_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8476_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8480_));
OR2X2 OR2X2_4474 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8481_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8482_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8483_));
OR2X2 OR2X2_4475 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8485_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8484_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8486_));
OR2X2 OR2X2_4476 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8483_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8486_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8487_));
OR2X2 OR2X2_4477 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8487_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8480_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8488_));
OR2X2 OR2X2_4478 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8488_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8475_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8489_));
OR2X2 OR2X2_4479 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8491_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8490_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8492_));
OR2X2 OR2X2_448 ( .A(_abc_44694_new_n1949_), .B(_abc_44694_new_n1928_), .Y(_abc_44694_new_n1950_));
OR2X2 OR2X2_4480 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8493_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8494_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8495_));
OR2X2 OR2X2_4481 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8492_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8496_));
OR2X2 OR2X2_4482 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8497_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8498_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8499_));
OR2X2 OR2X2_4483 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8500_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8501_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8502_));
OR2X2 OR2X2_4484 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8499_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8502_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8503_));
OR2X2 OR2X2_4485 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8503_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8496_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8504_));
OR2X2 OR2X2_4486 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8505_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8506_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8507_));
OR2X2 OR2X2_4487 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8508_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8509_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8510_));
OR2X2 OR2X2_4488 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8507_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8510_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8511_));
OR2X2 OR2X2_4489 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8512_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8513_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8514_));
OR2X2 OR2X2_449 ( .A(_abc_44694_new_n1400__bF_buf0), .B(_abc_44694_new_n1952_), .Y(_abc_44694_new_n1953_));
OR2X2 OR2X2_4490 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8515_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8516_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8517_));
OR2X2 OR2X2_4491 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8514_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8518_));
OR2X2 OR2X2_4492 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8511_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8518_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8519_));
OR2X2 OR2X2_4493 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8519_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8504_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8520_));
OR2X2 OR2X2_4494 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8489_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8520_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_14_));
OR2X2 OR2X2_4495 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8523_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8522_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8524_));
OR2X2 OR2X2_4496 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8525_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8526_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8527_));
OR2X2 OR2X2_4497 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8527_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8524_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8528_));
OR2X2 OR2X2_4498 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8529_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8530_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8531_));
OR2X2 OR2X2_4499 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8532_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8533_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8534_));
OR2X2 OR2X2_45 ( .A(_abc_44694_new_n770_), .B(_abc_44694_new_n773_), .Y(_abc_44694_new_n774_));
OR2X2 OR2X2_450 ( .A(_abc_44694_new_n1951_), .B(_abc_44694_new_n1953_), .Y(_abc_44694_new_n1954_));
OR2X2 OR2X2_4500 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8534_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8531_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8535_));
OR2X2 OR2X2_4501 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8535_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8528_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8536_));
OR2X2 OR2X2_4502 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8538_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8540_));
OR2X2 OR2X2_4503 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8540_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8537_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8541_));
OR2X2 OR2X2_4504 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8542_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8544_));
OR2X2 OR2X2_4505 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8546_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8545_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8547_));
OR2X2 OR2X2_4506 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8544_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8547_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8548_));
OR2X2 OR2X2_4507 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8548_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8549_));
OR2X2 OR2X2_4508 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8549_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8536_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8550_));
OR2X2 OR2X2_4509 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8552_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8551_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8553_));
OR2X2 OR2X2_451 ( .A(_abc_44694_new_n1955_), .B(_abc_44694_new_n1278__bF_buf4), .Y(_abc_44694_new_n1956_));
OR2X2 OR2X2_4510 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8554_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8555_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8556_));
OR2X2 OR2X2_4511 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8557_));
OR2X2 OR2X2_4512 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8558_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8559_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8560_));
OR2X2 OR2X2_4513 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8561_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8562_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8563_));
OR2X2 OR2X2_4514 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8560_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8563_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8564_));
OR2X2 OR2X2_4515 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8564_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8557_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8565_));
OR2X2 OR2X2_4516 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8566_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8567_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8568_));
OR2X2 OR2X2_4517 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8569_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8570_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8571_));
OR2X2 OR2X2_4518 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8568_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8571_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8572_));
OR2X2 OR2X2_4519 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8573_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8574_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8575_));
OR2X2 OR2X2_452 ( .A(_abc_44694_new_n1957_), .B(_abc_44694_new_n1958_), .Y(_abc_44694_new_n1959_));
OR2X2 OR2X2_4520 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8576_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8577_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8578_));
OR2X2 OR2X2_4521 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8575_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8578_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8579_));
OR2X2 OR2X2_4522 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8572_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8579_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8580_));
OR2X2 OR2X2_4523 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8580_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8565_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8581_));
OR2X2 OR2X2_4524 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8550_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8581_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_15_));
OR2X2 OR2X2_4525 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8584_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8583_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8585_));
OR2X2 OR2X2_4526 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8586_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8587_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8588_));
OR2X2 OR2X2_4527 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8588_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8585_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8589_));
OR2X2 OR2X2_4528 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8590_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8591_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8592_));
OR2X2 OR2X2_4529 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8593_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8594_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8595_));
OR2X2 OR2X2_453 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n1959_), .Y(_abc_44694_new_n1960_));
OR2X2 OR2X2_4530 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8595_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8592_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8596_));
OR2X2 OR2X2_4531 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8596_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8589_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8597_));
OR2X2 OR2X2_4532 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8599_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8600_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8601_));
OR2X2 OR2X2_4533 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8601_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8598_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8602_));
OR2X2 OR2X2_4534 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8603_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8604_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8605_));
OR2X2 OR2X2_4535 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8607_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8606_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8608_));
OR2X2 OR2X2_4536 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8605_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8608_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8609_));
OR2X2 OR2X2_4537 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8609_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8602_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8610_));
OR2X2 OR2X2_4538 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8610_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8597_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8611_));
OR2X2 OR2X2_4539 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8613_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8612_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8614_));
OR2X2 OR2X2_454 ( .A(_abc_44694_new_n1962_), .B(_abc_44694_new_n1926_), .Y(_abc_44694_new_n1963_));
OR2X2 OR2X2_4540 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8615_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8616_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8617_));
OR2X2 OR2X2_4541 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8617_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8614_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8618_));
OR2X2 OR2X2_4542 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8619_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8620_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8621_));
OR2X2 OR2X2_4543 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8622_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8623_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8624_));
OR2X2 OR2X2_4544 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8621_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8624_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8625_));
OR2X2 OR2X2_4545 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8625_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8618_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8626_));
OR2X2 OR2X2_4546 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8627_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8628_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8629_));
OR2X2 OR2X2_4547 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8630_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8631_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8632_));
OR2X2 OR2X2_4548 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8629_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8632_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8633_));
OR2X2 OR2X2_4549 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8634_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8635_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8636_));
OR2X2 OR2X2_455 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_16_), .Y(_abc_44694_new_n1964_));
OR2X2 OR2X2_4550 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8637_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8638_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8639_));
OR2X2 OR2X2_4551 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8636_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8639_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8640_));
OR2X2 OR2X2_4552 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8633_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8640_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8641_));
OR2X2 OR2X2_4553 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8641_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8626_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8642_));
OR2X2 OR2X2_4554 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8611_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8642_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_16_));
OR2X2 OR2X2_4555 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8645_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8644_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8646_));
OR2X2 OR2X2_4556 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8647_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8648_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8649_));
OR2X2 OR2X2_4557 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8649_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8646_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8650_));
OR2X2 OR2X2_4558 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8651_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8652_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8653_));
OR2X2 OR2X2_4559 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8654_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8655_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8656_));
OR2X2 OR2X2_456 ( .A(_abc_44694_new_n1922_), .B(pc_q_17_), .Y(_abc_44694_new_n1967_));
OR2X2 OR2X2_4560 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8656_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8653_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8657_));
OR2X2 OR2X2_4561 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8657_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8650_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8658_));
OR2X2 OR2X2_4562 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8660_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8661_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8662_));
OR2X2 OR2X2_4563 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8662_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8659_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8663_));
OR2X2 OR2X2_4564 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8664_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8665_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8666_));
OR2X2 OR2X2_4565 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8668_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8667_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8669_));
OR2X2 OR2X2_4566 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8666_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8669_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8670_));
OR2X2 OR2X2_4567 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8670_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8663_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8671_));
OR2X2 OR2X2_4568 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8671_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8658_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8672_));
OR2X2 OR2X2_4569 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8674_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8673_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8675_));
OR2X2 OR2X2_457 ( .A(_abc_44694_new_n1970_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n1971_));
OR2X2 OR2X2_4570 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8676_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8677_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8678_));
OR2X2 OR2X2_4571 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8678_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8675_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8679_));
OR2X2 OR2X2_4572 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8680_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8681_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8682_));
OR2X2 OR2X2_4573 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8683_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8684_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8685_));
OR2X2 OR2X2_4574 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8682_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8685_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8686_));
OR2X2 OR2X2_4575 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8686_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8679_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8687_));
OR2X2 OR2X2_4576 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8688_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8689_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8690_));
OR2X2 OR2X2_4577 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8691_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8692_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8693_));
OR2X2 OR2X2_4578 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8690_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8693_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8694_));
OR2X2 OR2X2_4579 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8695_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8696_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8697_));
OR2X2 OR2X2_458 ( .A(_abc_44694_new_n1970_), .B(_abc_44694_new_n1399__bF_buf3), .Y(_abc_44694_new_n1973_));
OR2X2 OR2X2_4580 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8698_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8699_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8700_));
OR2X2 OR2X2_4581 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8697_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8700_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8701_));
OR2X2 OR2X2_4582 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8694_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8701_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8702_));
OR2X2 OR2X2_4583 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8702_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8687_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8703_));
OR2X2 OR2X2_4584 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8672_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8703_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_17_));
OR2X2 OR2X2_4585 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8706_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8705_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8707_));
OR2X2 OR2X2_4586 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8708_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8709_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8710_));
OR2X2 OR2X2_4587 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8710_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8707_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8711_));
OR2X2 OR2X2_4588 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8712_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8713_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8714_));
OR2X2 OR2X2_4589 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8715_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8716_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8717_));
OR2X2 OR2X2_459 ( .A(pc_q_17_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf5_), .Y(_abc_44694_new_n1975_));
OR2X2 OR2X2_4590 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8717_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8714_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8718_));
OR2X2 OR2X2_4591 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8718_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8711_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8719_));
OR2X2 OR2X2_4592 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8721_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8722_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8723_));
OR2X2 OR2X2_4593 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8723_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8720_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8724_));
OR2X2 OR2X2_4594 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8725_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8726_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8727_));
OR2X2 OR2X2_4595 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8729_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8728_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8730_));
OR2X2 OR2X2_4596 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8727_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8730_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8731_));
OR2X2 OR2X2_4597 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8731_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8724_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8732_));
OR2X2 OR2X2_4598 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8732_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8719_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8733_));
OR2X2 OR2X2_4599 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8735_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8734_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8736_));
OR2X2 OR2X2_46 ( .A(_abc_44694_new_n767_), .B(_abc_44694_new_n775_), .Y(_abc_44694_new_n776_));
OR2X2 OR2X2_460 ( .A(_abc_44694_new_n1980_), .B(_abc_44694_new_n1978_), .Y(_abc_44694_new_n1983_));
OR2X2 OR2X2_4600 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8737_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8738_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8739_));
OR2X2 OR2X2_4601 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8739_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8736_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8740_));
OR2X2 OR2X2_4602 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8741_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8742_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8743_));
OR2X2 OR2X2_4603 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8744_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8745_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8746_));
OR2X2 OR2X2_4604 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8743_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8746_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8747_));
OR2X2 OR2X2_4605 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8747_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8740_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8748_));
OR2X2 OR2X2_4606 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8749_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8750_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8751_));
OR2X2 OR2X2_4607 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8752_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8753_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8754_));
OR2X2 OR2X2_4608 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8751_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8754_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8755_));
OR2X2 OR2X2_4609 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8756_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8757_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8758_));
OR2X2 OR2X2_461 ( .A(_abc_44694_new_n1985_), .B(_abc_44694_new_n1974_), .Y(_abc_44694_new_n1986_));
OR2X2 OR2X2_4610 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8759_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8760_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8761_));
OR2X2 OR2X2_4611 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8758_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8761_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8762_));
OR2X2 OR2X2_4612 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8755_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8762_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8763_));
OR2X2 OR2X2_4613 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8763_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8748_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8764_));
OR2X2 OR2X2_4614 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8733_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8764_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_18_));
OR2X2 OR2X2_4615 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8767_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8766_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8768_));
OR2X2 OR2X2_4616 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8769_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8770_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8771_));
OR2X2 OR2X2_4617 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8771_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8768_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8772_));
OR2X2 OR2X2_4618 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8773_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8774_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8775_));
OR2X2 OR2X2_4619 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8776_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8777_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8778_));
OR2X2 OR2X2_462 ( .A(_abc_44694_new_n1400__bF_buf4), .B(_abc_44694_new_n1988_), .Y(_abc_44694_new_n1989_));
OR2X2 OR2X2_4620 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8778_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8775_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8779_));
OR2X2 OR2X2_4621 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8779_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8772_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8780_));
OR2X2 OR2X2_4622 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8782_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8783_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8784_));
OR2X2 OR2X2_4623 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8784_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8781_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8785_));
OR2X2 OR2X2_4624 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8786_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8787_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8788_));
OR2X2 OR2X2_4625 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8790_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8789_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8791_));
OR2X2 OR2X2_4626 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8788_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8791_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8792_));
OR2X2 OR2X2_4627 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8792_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8785_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8793_));
OR2X2 OR2X2_4628 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8793_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8780_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8794_));
OR2X2 OR2X2_4629 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8796_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8795_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8797_));
OR2X2 OR2X2_463 ( .A(_abc_44694_new_n1987_), .B(_abc_44694_new_n1989_), .Y(_abc_44694_new_n1990_));
OR2X2 OR2X2_4630 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8798_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8799_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8800_));
OR2X2 OR2X2_4631 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8800_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8797_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8801_));
OR2X2 OR2X2_4632 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8802_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8803_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8804_));
OR2X2 OR2X2_4633 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8805_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8806_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8807_));
OR2X2 OR2X2_4634 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8804_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8807_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8808_));
OR2X2 OR2X2_4635 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8808_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8801_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8809_));
OR2X2 OR2X2_4636 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8810_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8811_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8812_));
OR2X2 OR2X2_4637 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8813_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8814_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8815_));
OR2X2 OR2X2_4638 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8812_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8815_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8816_));
OR2X2 OR2X2_4639 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8817_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8818_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8819_));
OR2X2 OR2X2_464 ( .A(_abc_44694_new_n1991_), .B(_abc_44694_new_n1278__bF_buf3), .Y(_abc_44694_new_n1992_));
OR2X2 OR2X2_4640 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8820_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8821_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8822_));
OR2X2 OR2X2_4641 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8819_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8822_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8823_));
OR2X2 OR2X2_4642 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8816_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8823_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8824_));
OR2X2 OR2X2_4643 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8824_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8809_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8825_));
OR2X2 OR2X2_4644 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8794_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8825_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_19_));
OR2X2 OR2X2_4645 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8828_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8827_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8829_));
OR2X2 OR2X2_4646 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8830_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8831_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8832_));
OR2X2 OR2X2_4647 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8832_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8829_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8833_));
OR2X2 OR2X2_4648 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8834_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8835_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8836_));
OR2X2 OR2X2_4649 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8837_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8838_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8839_));
OR2X2 OR2X2_465 ( .A(_abc_44694_new_n1993_), .B(_abc_44694_new_n1994_), .Y(_abc_44694_new_n1995_));
OR2X2 OR2X2_4650 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8839_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8836_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8840_));
OR2X2 OR2X2_4651 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8840_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8833_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8841_));
OR2X2 OR2X2_4652 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8843_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8844_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8845_));
OR2X2 OR2X2_4653 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8845_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8842_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8846_));
OR2X2 OR2X2_4654 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8847_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8848_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8849_));
OR2X2 OR2X2_4655 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8851_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8850_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8852_));
OR2X2 OR2X2_4656 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8849_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8852_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8853_));
OR2X2 OR2X2_4657 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8853_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8846_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8854_));
OR2X2 OR2X2_4658 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8854_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8841_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8855_));
OR2X2 OR2X2_4659 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8857_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8856_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8858_));
OR2X2 OR2X2_466 ( .A(_abc_44694_new_n1334__bF_buf2), .B(_abc_44694_new_n1995_), .Y(_abc_44694_new_n1996_));
OR2X2 OR2X2_4660 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8859_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8860_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8861_));
OR2X2 OR2X2_4661 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8861_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8858_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8862_));
OR2X2 OR2X2_4662 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8863_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8864_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8865_));
OR2X2 OR2X2_4663 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8866_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8867_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8868_));
OR2X2 OR2X2_4664 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8865_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8868_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8869_));
OR2X2 OR2X2_4665 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8869_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8862_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8870_));
OR2X2 OR2X2_4666 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8871_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8872_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8873_));
OR2X2 OR2X2_4667 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8874_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8875_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8876_));
OR2X2 OR2X2_4668 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8873_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8876_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8877_));
OR2X2 OR2X2_4669 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8878_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8879_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8880_));
OR2X2 OR2X2_467 ( .A(_abc_44694_new_n1998_), .B(_abc_44694_new_n1972_), .Y(_abc_44694_new_n1999_));
OR2X2 OR2X2_4670 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8881_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8882_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8883_));
OR2X2 OR2X2_4671 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8880_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8883_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8884_));
OR2X2 OR2X2_4672 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8877_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8884_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8885_));
OR2X2 OR2X2_4673 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8885_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8870_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8886_));
OR2X2 OR2X2_4674 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8855_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8886_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_20_));
OR2X2 OR2X2_4675 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8889_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8888_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8890_));
OR2X2 OR2X2_4676 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8891_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8892_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8893_));
OR2X2 OR2X2_4677 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8893_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8890_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8894_));
OR2X2 OR2X2_4678 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8895_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8896_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8897_));
OR2X2 OR2X2_4679 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8898_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8899_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8900_));
OR2X2 OR2X2_468 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(epc_q_17_), .Y(_abc_44694_new_n2000_));
OR2X2 OR2X2_4680 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8900_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8897_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8901_));
OR2X2 OR2X2_4681 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8901_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8894_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8902_));
OR2X2 OR2X2_4682 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8904_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8905_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8906_));
OR2X2 OR2X2_4683 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8906_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8903_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8907_));
OR2X2 OR2X2_4684 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8908_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8909_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8910_));
OR2X2 OR2X2_4685 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8912_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8911_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8913_));
OR2X2 OR2X2_4686 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8910_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8913_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8914_));
OR2X2 OR2X2_4687 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8914_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8907_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8915_));
OR2X2 OR2X2_4688 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8915_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8902_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8916_));
OR2X2 OR2X2_4689 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8918_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8917_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8919_));
OR2X2 OR2X2_469 ( .A(_abc_44694_new_n1968_), .B(pc_q_18_), .Y(_abc_44694_new_n2003_));
OR2X2 OR2X2_4690 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8920_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8921_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8922_));
OR2X2 OR2X2_4691 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8922_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8919_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8923_));
OR2X2 OR2X2_4692 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8924_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8925_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8926_));
OR2X2 OR2X2_4693 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8927_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8928_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8929_));
OR2X2 OR2X2_4694 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8926_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8929_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8930_));
OR2X2 OR2X2_4695 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8930_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8923_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8931_));
OR2X2 OR2X2_4696 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8932_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8933_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8934_));
OR2X2 OR2X2_4697 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8935_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8936_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8937_));
OR2X2 OR2X2_4698 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8934_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8937_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8938_));
OR2X2 OR2X2_4699 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8939_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8940_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8941_));
OR2X2 OR2X2_47 ( .A(_abc_44694_new_n777_), .B(_abc_44694_new_n763_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_5_));
OR2X2 OR2X2_470 ( .A(_abc_44694_new_n2007_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n2008_));
OR2X2 OR2X2_4700 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8942_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8943_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8944_));
OR2X2 OR2X2_4701 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8941_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8944_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8945_));
OR2X2 OR2X2_4702 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8938_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8945_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8946_));
OR2X2 OR2X2_4703 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8946_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8931_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8947_));
OR2X2 OR2X2_4704 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8916_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8947_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_21_));
OR2X2 OR2X2_4705 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8950_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8949_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8951_));
OR2X2 OR2X2_4706 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8952_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8953_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8954_));
OR2X2 OR2X2_4707 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8954_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8951_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8955_));
OR2X2 OR2X2_4708 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8956_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8957_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8958_));
OR2X2 OR2X2_4709 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8959_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8960_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8961_));
OR2X2 OR2X2_471 ( .A(_abc_44694_new_n2006_), .B(_abc_44694_new_n1399__bF_buf2), .Y(_abc_44694_new_n2009_));
OR2X2 OR2X2_4710 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8961_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8958_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8962_));
OR2X2 OR2X2_4711 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8962_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8955_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8963_));
OR2X2 OR2X2_4712 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8965_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8966_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8967_));
OR2X2 OR2X2_4713 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8967_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8964_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8968_));
OR2X2 OR2X2_4714 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8969_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8970_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8971_));
OR2X2 OR2X2_4715 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8973_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8972_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8974_));
OR2X2 OR2X2_4716 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8971_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8974_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8975_));
OR2X2 OR2X2_4717 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8975_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8968_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8976_));
OR2X2 OR2X2_4718 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8976_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8963_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8977_));
OR2X2 OR2X2_4719 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8979_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8978_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8980_));
OR2X2 OR2X2_472 ( .A(pc_q_18_), .B(REGFILE_SIM_reg_bank_ra_i_0_), .Y(_abc_44694_new_n2013_));
OR2X2 OR2X2_4720 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8981_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8982_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8983_));
OR2X2 OR2X2_4721 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8983_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8980_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8984_));
OR2X2 OR2X2_4722 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8985_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8986_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8987_));
OR2X2 OR2X2_4723 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8988_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8989_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8990_));
OR2X2 OR2X2_4724 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8987_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8990_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8991_));
OR2X2 OR2X2_4725 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8991_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8984_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8992_));
OR2X2 OR2X2_4726 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8993_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8994_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8995_));
OR2X2 OR2X2_4727 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8996_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8997_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8998_));
OR2X2 OR2X2_4728 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8995_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8998_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n8999_));
OR2X2 OR2X2_4729 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9000_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9001_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9002_));
OR2X2 OR2X2_473 ( .A(_abc_44694_new_n2012_), .B(_abc_44694_new_n2016_), .Y(_abc_44694_new_n2019_));
OR2X2 OR2X2_4730 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9003_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9004_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9005_));
OR2X2 OR2X2_4731 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9002_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9005_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9006_));
OR2X2 OR2X2_4732 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8999_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9006_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9007_));
OR2X2 OR2X2_4733 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9007_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n8992_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9008_));
OR2X2 OR2X2_4734 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n8977_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9008_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_22_));
OR2X2 OR2X2_4735 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9011_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9010_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9012_));
OR2X2 OR2X2_4736 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9013_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9014_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9015_));
OR2X2 OR2X2_4737 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9015_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9012_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9016_));
OR2X2 OR2X2_4738 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9017_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9018_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9019_));
OR2X2 OR2X2_4739 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9020_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9021_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9022_));
OR2X2 OR2X2_474 ( .A(_abc_44694_new_n2021_), .B(_abc_44694_new_n2010_), .Y(_abc_44694_new_n2022_));
OR2X2 OR2X2_4740 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9022_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9019_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9023_));
OR2X2 OR2X2_4741 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9023_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9016_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9024_));
OR2X2 OR2X2_4742 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9026_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9027_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9028_));
OR2X2 OR2X2_4743 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9028_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9025_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9029_));
OR2X2 OR2X2_4744 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9030_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9031_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9032_));
OR2X2 OR2X2_4745 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9034_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9033_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9035_));
OR2X2 OR2X2_4746 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9032_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9035_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9036_));
OR2X2 OR2X2_4747 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9036_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9029_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9037_));
OR2X2 OR2X2_4748 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9037_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9024_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9038_));
OR2X2 OR2X2_4749 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9040_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9039_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9041_));
OR2X2 OR2X2_475 ( .A(_abc_44694_new_n1400__bF_buf3), .B(_abc_44694_new_n2024_), .Y(_abc_44694_new_n2025_));
OR2X2 OR2X2_4750 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9042_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9043_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9044_));
OR2X2 OR2X2_4751 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9044_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9041_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9045_));
OR2X2 OR2X2_4752 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9046_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9047_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9048_));
OR2X2 OR2X2_4753 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9049_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9050_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9051_));
OR2X2 OR2X2_4754 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9048_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9051_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9052_));
OR2X2 OR2X2_4755 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9052_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9045_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9053_));
OR2X2 OR2X2_4756 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9054_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9055_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9056_));
OR2X2 OR2X2_4757 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9057_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9058_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9059_));
OR2X2 OR2X2_4758 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9056_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9059_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9060_));
OR2X2 OR2X2_4759 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9061_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9062_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9063_));
OR2X2 OR2X2_476 ( .A(_abc_44694_new_n2023_), .B(_abc_44694_new_n2025_), .Y(_abc_44694_new_n2026_));
OR2X2 OR2X2_4760 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9064_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9065_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9066_));
OR2X2 OR2X2_4761 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9063_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9066_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9067_));
OR2X2 OR2X2_4762 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9060_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9067_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9068_));
OR2X2 OR2X2_4763 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9068_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9053_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9069_));
OR2X2 OR2X2_4764 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9038_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9069_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_23_));
OR2X2 OR2X2_4765 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9072_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9071_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9073_));
OR2X2 OR2X2_4766 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9074_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9075_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9076_));
OR2X2 OR2X2_4767 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9076_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9073_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9077_));
OR2X2 OR2X2_4768 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9078_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9079_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9080_));
OR2X2 OR2X2_4769 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9081_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9082_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9083_));
OR2X2 OR2X2_477 ( .A(_abc_44694_new_n2027_), .B(_abc_44694_new_n1278__bF_buf2), .Y(_abc_44694_new_n2028_));
OR2X2 OR2X2_4770 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9083_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9080_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9084_));
OR2X2 OR2X2_4771 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9084_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9077_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9085_));
OR2X2 OR2X2_4772 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9087_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9088_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9089_));
OR2X2 OR2X2_4773 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9089_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9086_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9090_));
OR2X2 OR2X2_4774 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9091_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9092_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9093_));
OR2X2 OR2X2_4775 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9095_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9094_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9096_));
OR2X2 OR2X2_4776 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9093_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9096_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9097_));
OR2X2 OR2X2_4777 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9097_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9090_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9098_));
OR2X2 OR2X2_4778 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9098_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9085_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9099_));
OR2X2 OR2X2_4779 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9101_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9100_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9102_));
OR2X2 OR2X2_478 ( .A(_abc_44694_new_n2029_), .B(_abc_44694_new_n2030_), .Y(_abc_44694_new_n2031_));
OR2X2 OR2X2_4780 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9103_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9104_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9105_));
OR2X2 OR2X2_4781 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9105_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9102_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9106_));
OR2X2 OR2X2_4782 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9107_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9108_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9109_));
OR2X2 OR2X2_4783 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9110_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9111_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9112_));
OR2X2 OR2X2_4784 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9109_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9112_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9113_));
OR2X2 OR2X2_4785 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9113_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9106_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9114_));
OR2X2 OR2X2_4786 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9115_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9116_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9117_));
OR2X2 OR2X2_4787 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9118_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9119_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9120_));
OR2X2 OR2X2_4788 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9117_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9120_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9121_));
OR2X2 OR2X2_4789 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9122_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9123_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9124_));
OR2X2 OR2X2_479 ( .A(_abc_44694_new_n1334__bF_buf1), .B(_abc_44694_new_n2031_), .Y(_abc_44694_new_n2032_));
OR2X2 OR2X2_4790 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9125_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9126_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9127_));
OR2X2 OR2X2_4791 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9124_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9127_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9128_));
OR2X2 OR2X2_4792 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9121_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9128_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9129_));
OR2X2 OR2X2_4793 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9129_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9114_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9130_));
OR2X2 OR2X2_4794 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9099_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9130_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_24_));
OR2X2 OR2X2_4795 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9133_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9132_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9134_));
OR2X2 OR2X2_4796 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9135_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9136_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9137_));
OR2X2 OR2X2_4797 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9137_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9134_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9138_));
OR2X2 OR2X2_4798 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9139_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9140_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9141_));
OR2X2 OR2X2_4799 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9142_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9143_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9144_));
OR2X2 OR2X2_48 ( .A(_abc_44694_new_n781_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n782_));
OR2X2 OR2X2_480 ( .A(_abc_44694_new_n2034_), .B(_abc_44694_new_n2008_), .Y(_abc_44694_new_n2035_));
OR2X2 OR2X2_4800 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9144_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9141_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9145_));
OR2X2 OR2X2_4801 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9145_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9138_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9146_));
OR2X2 OR2X2_4802 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9148_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9149_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9150_));
OR2X2 OR2X2_4803 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9150_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9147_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9151_));
OR2X2 OR2X2_4804 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9152_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9153_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9154_));
OR2X2 OR2X2_4805 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9156_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9155_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9157_));
OR2X2 OR2X2_4806 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9154_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9157_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9158_));
OR2X2 OR2X2_4807 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9158_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9151_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9159_));
OR2X2 OR2X2_4808 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9159_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9146_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9160_));
OR2X2 OR2X2_4809 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9162_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9161_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9163_));
OR2X2 OR2X2_481 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(epc_q_18_), .Y(_abc_44694_new_n2036_));
OR2X2 OR2X2_4810 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9164_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9165_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9166_));
OR2X2 OR2X2_4811 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9166_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9163_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9167_));
OR2X2 OR2X2_4812 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9168_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9169_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9170_));
OR2X2 OR2X2_4813 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9171_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9172_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9173_));
OR2X2 OR2X2_4814 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9170_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9173_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9174_));
OR2X2 OR2X2_4815 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9174_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9167_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9175_));
OR2X2 OR2X2_4816 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9176_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9177_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9178_));
OR2X2 OR2X2_4817 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9179_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9180_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9181_));
OR2X2 OR2X2_4818 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9178_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9181_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9182_));
OR2X2 OR2X2_4819 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9183_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9184_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9185_));
OR2X2 OR2X2_482 ( .A(_abc_44694_new_n2004_), .B(pc_q_19_), .Y(_abc_44694_new_n2039_));
OR2X2 OR2X2_4820 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9186_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9187_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9188_));
OR2X2 OR2X2_4821 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9185_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9188_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9189_));
OR2X2 OR2X2_4822 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9182_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9189_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9190_));
OR2X2 OR2X2_4823 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9190_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9175_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9191_));
OR2X2 OR2X2_4824 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9160_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9191_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_25_));
OR2X2 OR2X2_4825 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9194_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9193_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9195_));
OR2X2 OR2X2_4826 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9196_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9197_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9198_));
OR2X2 OR2X2_4827 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9198_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9195_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9199_));
OR2X2 OR2X2_4828 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9200_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9201_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9202_));
OR2X2 OR2X2_4829 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9203_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9204_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9205_));
OR2X2 OR2X2_483 ( .A(_abc_44694_new_n2043_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n2044_));
OR2X2 OR2X2_4830 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9205_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9202_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9206_));
OR2X2 OR2X2_4831 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9206_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9199_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9207_));
OR2X2 OR2X2_4832 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9209_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9210_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9211_));
OR2X2 OR2X2_4833 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9211_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9208_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9212_));
OR2X2 OR2X2_4834 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9213_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9214_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9215_));
OR2X2 OR2X2_4835 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9217_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9216_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9218_));
OR2X2 OR2X2_4836 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9215_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9218_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9219_));
OR2X2 OR2X2_4837 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9219_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9212_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9220_));
OR2X2 OR2X2_4838 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9220_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9207_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9221_));
OR2X2 OR2X2_4839 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9223_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9222_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9224_));
OR2X2 OR2X2_484 ( .A(_abc_44694_new_n2042_), .B(_abc_44694_new_n1399__bF_buf1), .Y(_abc_44694_new_n2045_));
OR2X2 OR2X2_4840 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9225_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9226_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9227_));
OR2X2 OR2X2_4841 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9227_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9224_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9228_));
OR2X2 OR2X2_4842 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9229_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9230_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9231_));
OR2X2 OR2X2_4843 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9232_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9233_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9234_));
OR2X2 OR2X2_4844 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9231_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9234_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9235_));
OR2X2 OR2X2_4845 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9235_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9228_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9236_));
OR2X2 OR2X2_4846 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9237_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9238_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9239_));
OR2X2 OR2X2_4847 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9240_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9241_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9242_));
OR2X2 OR2X2_4848 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9239_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9242_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9243_));
OR2X2 OR2X2_4849 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9244_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9245_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9246_));
OR2X2 OR2X2_485 ( .A(pc_q_19_), .B(REGFILE_SIM_reg_bank_ra_i_1_), .Y(_abc_44694_new_n2048_));
OR2X2 OR2X2_4850 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9247_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9248_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9249_));
OR2X2 OR2X2_4851 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9246_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9249_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9250_));
OR2X2 OR2X2_4852 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9243_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9250_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9251_));
OR2X2 OR2X2_4853 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9251_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9236_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9252_));
OR2X2 OR2X2_4854 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9221_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9252_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_26_));
OR2X2 OR2X2_4855 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9255_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9254_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9256_));
OR2X2 OR2X2_4856 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9257_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9258_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9259_));
OR2X2 OR2X2_4857 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9259_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9256_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9260_));
OR2X2 OR2X2_4858 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9261_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9262_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9263_));
OR2X2 OR2X2_4859 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9264_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9265_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9266_));
OR2X2 OR2X2_486 ( .A(_abc_44694_new_n2047_), .B(_abc_44694_new_n2052_), .Y(_abc_44694_new_n2053_));
OR2X2 OR2X2_4860 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9266_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9263_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9267_));
OR2X2 OR2X2_4861 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9267_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9260_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9268_));
OR2X2 OR2X2_4862 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9270_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9271_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9272_));
OR2X2 OR2X2_4863 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9272_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9269_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9273_));
OR2X2 OR2X2_4864 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9274_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9275_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9276_));
OR2X2 OR2X2_4865 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9278_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9277_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9279_));
OR2X2 OR2X2_4866 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9276_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9279_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9280_));
OR2X2 OR2X2_4867 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9280_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9273_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9281_));
OR2X2 OR2X2_4868 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9281_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9268_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9282_));
OR2X2 OR2X2_4869 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9284_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9283_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9285_));
OR2X2 OR2X2_487 ( .A(_abc_44694_new_n2054_), .B(_abc_44694_new_n2051_), .Y(_abc_44694_new_n2055_));
OR2X2 OR2X2_4870 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9286_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9287_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9288_));
OR2X2 OR2X2_4871 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9288_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9285_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9289_));
OR2X2 OR2X2_4872 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9290_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9291_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9292_));
OR2X2 OR2X2_4873 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9293_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9294_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9295_));
OR2X2 OR2X2_4874 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9292_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9295_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9296_));
OR2X2 OR2X2_4875 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9296_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9289_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9297_));
OR2X2 OR2X2_4876 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9298_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9299_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9300_));
OR2X2 OR2X2_4877 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9301_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9302_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9303_));
OR2X2 OR2X2_4878 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9300_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9303_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9304_));
OR2X2 OR2X2_4879 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9305_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9306_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9307_));
OR2X2 OR2X2_488 ( .A(_abc_44694_new_n2057_), .B(_abc_44694_new_n2046_), .Y(_abc_44694_new_n2058_));
OR2X2 OR2X2_4880 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9308_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9309_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9310_));
OR2X2 OR2X2_4881 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9307_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9310_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9311_));
OR2X2 OR2X2_4882 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9304_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9311_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9312_));
OR2X2 OR2X2_4883 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9312_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9297_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9313_));
OR2X2 OR2X2_4884 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9282_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9313_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_27_));
OR2X2 OR2X2_4885 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9316_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9315_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9317_));
OR2X2 OR2X2_4886 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9318_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9319_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9320_));
OR2X2 OR2X2_4887 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9320_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9317_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9321_));
OR2X2 OR2X2_4888 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9322_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9323_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9324_));
OR2X2 OR2X2_4889 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9325_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9326_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9327_));
OR2X2 OR2X2_489 ( .A(_abc_44694_new_n1400__bF_buf2), .B(_abc_44694_new_n2060_), .Y(_abc_44694_new_n2061_));
OR2X2 OR2X2_4890 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9327_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9324_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9328_));
OR2X2 OR2X2_4891 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9328_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9321_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9329_));
OR2X2 OR2X2_4892 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9331_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9332_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9333_));
OR2X2 OR2X2_4893 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9333_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9330_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9334_));
OR2X2 OR2X2_4894 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9335_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9336_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9337_));
OR2X2 OR2X2_4895 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9339_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9338_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9340_));
OR2X2 OR2X2_4896 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9337_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9340_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9341_));
OR2X2 OR2X2_4897 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9341_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9334_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9342_));
OR2X2 OR2X2_4898 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9342_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9329_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9343_));
OR2X2 OR2X2_4899 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9345_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9344_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9346_));
OR2X2 OR2X2_49 ( .A(_abc_44694_new_n782_), .B(_abc_44694_new_n780_), .Y(_abc_44694_new_n783_));
OR2X2 OR2X2_490 ( .A(_abc_44694_new_n2059_), .B(_abc_44694_new_n2061_), .Y(_abc_44694_new_n2062_));
OR2X2 OR2X2_4900 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9347_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9348_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9349_));
OR2X2 OR2X2_4901 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9349_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9346_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9350_));
OR2X2 OR2X2_4902 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9351_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9352_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9353_));
OR2X2 OR2X2_4903 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9354_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9355_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9356_));
OR2X2 OR2X2_4904 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9353_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9356_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9357_));
OR2X2 OR2X2_4905 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9357_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9350_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9358_));
OR2X2 OR2X2_4906 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9359_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9360_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9361_));
OR2X2 OR2X2_4907 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9362_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9363_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9364_));
OR2X2 OR2X2_4908 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9361_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9364_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9365_));
OR2X2 OR2X2_4909 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9366_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9367_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9368_));
OR2X2 OR2X2_491 ( .A(_abc_44694_new_n2063_), .B(_abc_44694_new_n1278__bF_buf1), .Y(_abc_44694_new_n2064_));
OR2X2 OR2X2_4910 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9369_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9370_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9371_));
OR2X2 OR2X2_4911 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9368_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9371_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9372_));
OR2X2 OR2X2_4912 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9365_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9372_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9373_));
OR2X2 OR2X2_4913 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9373_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9358_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9374_));
OR2X2 OR2X2_4914 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9343_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9374_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_28_));
OR2X2 OR2X2_4915 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9377_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9376_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9378_));
OR2X2 OR2X2_4916 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9379_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9380_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9381_));
OR2X2 OR2X2_4917 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9381_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9378_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9382_));
OR2X2 OR2X2_4918 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9383_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9384_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9385_));
OR2X2 OR2X2_4919 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9386_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9387_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9388_));
OR2X2 OR2X2_492 ( .A(_abc_44694_new_n2065_), .B(_abc_44694_new_n2066_), .Y(_abc_44694_new_n2067_));
OR2X2 OR2X2_4920 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9388_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9385_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9389_));
OR2X2 OR2X2_4921 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9389_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9382_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9390_));
OR2X2 OR2X2_4922 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9392_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9393_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9394_));
OR2X2 OR2X2_4923 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9394_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9391_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9395_));
OR2X2 OR2X2_4924 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9396_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9397_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9398_));
OR2X2 OR2X2_4925 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9400_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9399_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9401_));
OR2X2 OR2X2_4926 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9398_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9401_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9402_));
OR2X2 OR2X2_4927 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9402_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9395_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9403_));
OR2X2 OR2X2_4928 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9403_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9390_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9404_));
OR2X2 OR2X2_4929 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9406_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9405_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9407_));
OR2X2 OR2X2_493 ( .A(_abc_44694_new_n1334__bF_buf0), .B(_abc_44694_new_n2067_), .Y(_abc_44694_new_n2068_));
OR2X2 OR2X2_4930 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9408_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9409_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9410_));
OR2X2 OR2X2_4931 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9410_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9407_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9411_));
OR2X2 OR2X2_4932 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9412_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9413_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9414_));
OR2X2 OR2X2_4933 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9415_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9416_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9417_));
OR2X2 OR2X2_4934 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9414_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9417_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9418_));
OR2X2 OR2X2_4935 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9418_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9411_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9419_));
OR2X2 OR2X2_4936 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9420_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9421_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9422_));
OR2X2 OR2X2_4937 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9423_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9424_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9425_));
OR2X2 OR2X2_4938 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9422_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9425_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9426_));
OR2X2 OR2X2_4939 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9427_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9428_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9429_));
OR2X2 OR2X2_494 ( .A(_abc_44694_new_n2070_), .B(_abc_44694_new_n2044_), .Y(_abc_44694_new_n2071_));
OR2X2 OR2X2_4940 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9430_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9431_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9432_));
OR2X2 OR2X2_4941 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9429_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9432_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9433_));
OR2X2 OR2X2_4942 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9426_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9433_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9434_));
OR2X2 OR2X2_4943 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9434_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9419_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9435_));
OR2X2 OR2X2_4944 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9404_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9435_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_29_));
OR2X2 OR2X2_4945 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9438_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9437_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9439_));
OR2X2 OR2X2_4946 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9440_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9441_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9442_));
OR2X2 OR2X2_4947 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9442_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9439_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9443_));
OR2X2 OR2X2_4948 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9444_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9445_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9446_));
OR2X2 OR2X2_4949 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9447_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9448_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9449_));
OR2X2 OR2X2_495 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_19_), .Y(_abc_44694_new_n2072_));
OR2X2 OR2X2_4950 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9449_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9446_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9450_));
OR2X2 OR2X2_4951 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9450_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9443_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9451_));
OR2X2 OR2X2_4952 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9453_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9454_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9455_));
OR2X2 OR2X2_4953 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9455_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9452_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9456_));
OR2X2 OR2X2_4954 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9457_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9458_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9459_));
OR2X2 OR2X2_4955 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9461_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9460_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9462_));
OR2X2 OR2X2_4956 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9459_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9462_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9463_));
OR2X2 OR2X2_4957 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9463_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9456_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9464_));
OR2X2 OR2X2_4958 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9464_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9451_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9465_));
OR2X2 OR2X2_4959 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9467_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9466_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9468_));
OR2X2 OR2X2_496 ( .A(_abc_44694_new_n2040_), .B(pc_q_20_), .Y(_abc_44694_new_n2075_));
OR2X2 OR2X2_4960 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9469_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9470_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9471_));
OR2X2 OR2X2_4961 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9471_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9468_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9472_));
OR2X2 OR2X2_4962 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9473_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9474_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9475_));
OR2X2 OR2X2_4963 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9476_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9477_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9478_));
OR2X2 OR2X2_4964 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9475_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9478_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9479_));
OR2X2 OR2X2_4965 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9479_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9472_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9480_));
OR2X2 OR2X2_4966 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9481_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9482_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9483_));
OR2X2 OR2X2_4967 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9484_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9485_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9486_));
OR2X2 OR2X2_4968 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9483_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9486_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9487_));
OR2X2 OR2X2_4969 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9488_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9489_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9490_));
OR2X2 OR2X2_497 ( .A(_abc_44694_new_n2079_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n2080_));
OR2X2 OR2X2_4970 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9491_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9492_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9493_));
OR2X2 OR2X2_4971 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9490_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9493_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9494_));
OR2X2 OR2X2_4972 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9487_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9494_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9495_));
OR2X2 OR2X2_4973 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9495_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9480_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9496_));
OR2X2 OR2X2_4974 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9465_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9496_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_30_));
OR2X2 OR2X2_4975 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9499_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9498_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9500_));
OR2X2 OR2X2_4976 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9501_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9502_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9503_));
OR2X2 OR2X2_4977 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9503_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9500_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9504_));
OR2X2 OR2X2_4978 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9505_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9506_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9507_));
OR2X2 OR2X2_4979 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9508_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9509_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9510_));
OR2X2 OR2X2_498 ( .A(_abc_44694_new_n2078_), .B(_abc_44694_new_n1399__bF_buf0), .Y(_abc_44694_new_n2081_));
OR2X2 OR2X2_4980 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9510_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9507_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9511_));
OR2X2 OR2X2_4981 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9511_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9504_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9512_));
OR2X2 OR2X2_4982 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9514_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9515_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9516_));
OR2X2 OR2X2_4983 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9516_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9513_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9517_));
OR2X2 OR2X2_4984 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9518_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9519_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9520_));
OR2X2 OR2X2_4985 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9522_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9521_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9523_));
OR2X2 OR2X2_4986 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9520_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9523_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9524_));
OR2X2 OR2X2_4987 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9524_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9517_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9525_));
OR2X2 OR2X2_4988 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9525_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9512_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9526_));
OR2X2 OR2X2_4989 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9528_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9527_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9529_));
OR2X2 OR2X2_499 ( .A(_abc_44694_new_n2083_), .B(_abc_44694_new_n1976_), .Y(_abc_44694_new_n2084_));
OR2X2 OR2X2_4990 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9530_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9531_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9532_));
OR2X2 OR2X2_4991 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9532_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9529_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9533_));
OR2X2 OR2X2_4992 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9534_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9535_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9536_));
OR2X2 OR2X2_4993 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9537_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9538_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9539_));
OR2X2 OR2X2_4994 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9536_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9539_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9540_));
OR2X2 OR2X2_4995 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9540_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9533_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9541_));
OR2X2 OR2X2_4996 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9542_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9543_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9544_));
OR2X2 OR2X2_4997 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9545_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9546_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9547_));
OR2X2 OR2X2_4998 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9544_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9547_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9548_));
OR2X2 OR2X2_4999 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9549_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9550_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9551_));
OR2X2 OR2X2_5 ( .A(_abc_44694_new_n662_), .B(_abc_44694_new_n660_), .Y(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_3_));
OR2X2 OR2X2_50 ( .A(_abc_44694_new_n785_), .B(_abc_44694_new_n784_), .Y(_abc_44694_new_n786_));
OR2X2 OR2X2_500 ( .A(_abc_44694_new_n2087_), .B(_abc_44694_new_n2049_), .Y(_abc_44694_new_n2088_));
OR2X2 OR2X2_5000 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9552_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9553_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9554_));
OR2X2 OR2X2_5001 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9551_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9554_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9555_));
OR2X2 OR2X2_5002 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9548_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9555_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9556_));
OR2X2 OR2X2_5003 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9556_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9541_), .Y(REGFILE_SIM_reg_bank__abc_34819_new_n9557_));
OR2X2 OR2X2_5004 ( .A(REGFILE_SIM_reg_bank__abc_34819_new_n9526_), .B(REGFILE_SIM_reg_bank__abc_34819_new_n9557_), .Y(REGFILE_SIM_reg_bank_reg_ra_o_31_));
OR2X2 OR2X2_5005 ( .A(alu__abc_42281_new_n244_), .B(alu__abc_42281_new_n241_), .Y(alu__abc_42281_new_n245_));
OR2X2 OR2X2_5006 ( .A(alu__abc_42281_new_n261_), .B(alu__abc_42281_new_n258_), .Y(alu__abc_42281_new_n262_));
OR2X2 OR2X2_5007 ( .A(alu__abc_42281_new_n267_), .B(alu__abc_42281_new_n264_), .Y(alu__abc_42281_new_n268_));
OR2X2 OR2X2_5008 ( .A(alu__abc_42281_new_n282_), .B(alu__abc_42281_new_n279_), .Y(alu__abc_42281_new_n283_));
OR2X2 OR2X2_5009 ( .A(alu__abc_42281_new_n295_), .B(alu__abc_42281_new_n292_), .Y(alu__abc_42281_new_n296_));
OR2X2 OR2X2_501 ( .A(_abc_44694_new_n2086_), .B(_abc_44694_new_n2088_), .Y(_abc_44694_new_n2089_));
OR2X2 OR2X2_5010 ( .A(alu__abc_42281_new_n300_), .B(alu__abc_42281_new_n297_), .Y(alu__abc_42281_new_n301_));
OR2X2 OR2X2_5011 ( .A(alu__abc_42281_new_n287_), .B(alu__abc_42281_new_n400_), .Y(alu__abc_42281_new_n401_));
OR2X2 OR2X2_5012 ( .A(alu__abc_42281_new_n402_), .B(alu__abc_42281_new_n399_), .Y(alu__abc_42281_new_n403_));
OR2X2 OR2X2_5013 ( .A(alu__abc_42281_new_n404_), .B(alu__abc_42281_new_n396_), .Y(alu__abc_42281_new_n405_));
OR2X2 OR2X2_5014 ( .A(alu__abc_42281_new_n406_), .B(alu__abc_42281_new_n395_), .Y(alu__abc_42281_new_n407_));
OR2X2 OR2X2_5015 ( .A(alu__abc_42281_new_n408_), .B(alu__abc_42281_new_n392_), .Y(alu__abc_42281_new_n409_));
OR2X2 OR2X2_5016 ( .A(alu__abc_42281_new_n410_), .B(alu__abc_42281_new_n391_), .Y(alu__abc_42281_new_n411_));
OR2X2 OR2X2_5017 ( .A(alu__abc_42281_new_n412_), .B(alu__abc_42281_new_n388_), .Y(alu__abc_42281_new_n413_));
OR2X2 OR2X2_5018 ( .A(alu__abc_42281_new_n418_), .B(alu__abc_42281_new_n419_), .Y(alu__abc_42281_new_n420_));
OR2X2 OR2X2_5019 ( .A(alu__abc_42281_new_n426_), .B(alu__abc_42281_new_n424_), .Y(alu__abc_42281_new_n427_));
OR2X2 OR2X2_502 ( .A(_abc_44694_new_n2091_), .B(_abc_44694_new_n2094_), .Y(_abc_44694_new_n2095_));
OR2X2 OR2X2_5020 ( .A(alu__abc_42281_new_n427_), .B(alu__abc_42281_new_n423_), .Y(alu__abc_42281_new_n428_));
OR2X2 OR2X2_5021 ( .A(alu__abc_42281_new_n433_), .B(alu__abc_42281_new_n434_), .Y(alu__abc_42281_new_n435_));
OR2X2 OR2X2_5022 ( .A(alu__abc_42281_new_n441_), .B(alu__abc_42281_new_n439_), .Y(alu__abc_42281_new_n442_));
OR2X2 OR2X2_5023 ( .A(alu__abc_42281_new_n442_), .B(alu__abc_42281_new_n438_), .Y(alu__abc_42281_new_n443_));
OR2X2 OR2X2_5024 ( .A(alu__abc_42281_new_n429_), .B(alu__abc_42281_new_n443_), .Y(alu__abc_42281_new_n444_));
OR2X2 OR2X2_5025 ( .A(alu__abc_42281_new_n414_), .B(alu__abc_42281_new_n444_), .Y(alu__abc_42281_new_n445_));
OR2X2 OR2X2_5026 ( .A(alu__abc_42281_new_n450_), .B(alu__abc_42281_new_n451_), .Y(alu__abc_42281_new_n452_));
OR2X2 OR2X2_5027 ( .A(alu__abc_42281_new_n458_), .B(alu__abc_42281_new_n456_), .Y(alu__abc_42281_new_n459_));
OR2X2 OR2X2_5028 ( .A(alu__abc_42281_new_n459_), .B(alu__abc_42281_new_n455_), .Y(alu__abc_42281_new_n460_));
OR2X2 OR2X2_5029 ( .A(alu__abc_42281_new_n465_), .B(alu__abc_42281_new_n466_), .Y(alu__abc_42281_new_n467_));
OR2X2 OR2X2_503 ( .A(pc_q_20_), .B(REGFILE_SIM_reg_bank_ra_i_2_), .Y(_abc_44694_new_n2098_));
OR2X2 OR2X2_5030 ( .A(alu__abc_42281_new_n473_), .B(alu__abc_42281_new_n471_), .Y(alu__abc_42281_new_n474_));
OR2X2 OR2X2_5031 ( .A(alu__abc_42281_new_n474_), .B(alu__abc_42281_new_n470_), .Y(alu__abc_42281_new_n475_));
OR2X2 OR2X2_5032 ( .A(alu__abc_42281_new_n461_), .B(alu__abc_42281_new_n475_), .Y(alu__abc_42281_new_n476_));
OR2X2 OR2X2_5033 ( .A(alu__abc_42281_new_n446_), .B(alu__abc_42281_new_n476_), .Y(alu__abc_42281_new_n477_));
OR2X2 OR2X2_5034 ( .A(alu__abc_42281_new_n481_), .B(alu__abc_42281_new_n479_), .Y(alu__abc_42281_new_n482_));
OR2X2 OR2X2_5035 ( .A(alu__abc_42281_new_n490_), .B(alu__abc_42281_new_n485_), .Y(alu__abc_42281_new_n491_));
OR2X2 OR2X2_5036 ( .A(alu__abc_42281_new_n484_), .B(alu__abc_42281_new_n491_), .Y(alu__abc_42281_new_n492_));
OR2X2 OR2X2_5037 ( .A(alu__abc_42281_new_n478_), .B(alu__abc_42281_new_n494_), .Y(alu__abc_42281_new_n495_));
OR2X2 OR2X2_5038 ( .A(alu__abc_42281_new_n502_), .B(alu__abc_42281_new_n497_), .Y(alu__abc_42281_new_n503_));
OR2X2 OR2X2_5039 ( .A(alu__abc_42281_new_n496_), .B(alu__abc_42281_new_n504_), .Y(alu__abc_42281_new_n505_));
OR2X2 OR2X2_504 ( .A(_abc_44694_new_n2097_), .B(_abc_44694_new_n2101_), .Y(_abc_44694_new_n2104_));
OR2X2 OR2X2_5040 ( .A(alu__abc_42281_new_n506_), .B(alu__abc_42281_new_n507_), .Y(alu__abc_42281_new_n508_));
OR2X2 OR2X2_5041 ( .A(alu__abc_42281_new_n510_), .B(alu__abc_42281_new_n387_), .Y(alu_less_than_signed_o));
OR2X2 OR2X2_5042 ( .A(alu__abc_42281_new_n516_), .B(alu__abc_42281_new_n210_), .Y(alu__abc_42281_new_n517_));
OR2X2 OR2X2_5043 ( .A(alu__abc_42281_new_n520_), .B(alu__abc_42281_new_n185_), .Y(alu__abc_42281_new_n521_));
OR2X2 OR2X2_5044 ( .A(alu__abc_42281_new_n523_), .B(alu__abc_42281_new_n518_), .Y(alu__abc_42281_new_n524_));
OR2X2 OR2X2_5045 ( .A(alu__abc_42281_new_n526_), .B(alu__abc_42281_new_n228_), .Y(alu__abc_42281_new_n527_));
OR2X2 OR2X2_5046 ( .A(alu__abc_42281_new_n531_), .B(alu__abc_42281_new_n241_), .Y(alu__abc_42281_new_n532_));
OR2X2 OR2X2_5047 ( .A(alu__abc_42281_new_n529_), .B(alu__abc_42281_new_n532_), .Y(alu__abc_42281_new_n533_));
OR2X2 OR2X2_5048 ( .A(alu__abc_42281_new_n525_), .B(alu__abc_42281_new_n533_), .Y(alu__abc_42281_new_n534_));
OR2X2 OR2X2_5049 ( .A(alu__abc_42281_new_n539_), .B(alu__abc_42281_new_n174_), .Y(alu__abc_42281_new_n540_));
OR2X2 OR2X2_505 ( .A(_abc_44694_new_n2106_), .B(_abc_44694_new_n2082_), .Y(_abc_44694_new_n2107_));
OR2X2 OR2X2_5050 ( .A(alu__abc_42281_new_n543_), .B(alu__abc_42281_new_n153_), .Y(alu__abc_42281_new_n544_));
OR2X2 OR2X2_5051 ( .A(alu__abc_42281_new_n542_), .B(alu__abc_42281_new_n544_), .Y(alu__abc_42281_new_n545_));
OR2X2 OR2X2_5052 ( .A(alu__abc_42281_new_n547_), .B(alu__abc_42281_new_n122_), .Y(alu__abc_42281_new_n548_));
OR2X2 OR2X2_5053 ( .A(alu__abc_42281_new_n551_), .B(alu__abc_42281_new_n135_), .Y(alu__abc_42281_new_n552_));
OR2X2 OR2X2_5054 ( .A(alu__abc_42281_new_n550_), .B(alu__abc_42281_new_n552_), .Y(alu__abc_42281_new_n553_));
OR2X2 OR2X2_5055 ( .A(alu__abc_42281_new_n546_), .B(alu__abc_42281_new_n553_), .Y(alu__abc_42281_new_n554_));
OR2X2 OR2X2_5056 ( .A(alu__abc_42281_new_n555_), .B(alu__abc_42281_new_n330_), .Y(alu__abc_42281_new_n556_));
OR2X2 OR2X2_5057 ( .A(alu__abc_42281_new_n557_), .B(alu__abc_42281_new_n313_), .Y(alu__abc_42281_new_n558_));
OR2X2 OR2X2_5058 ( .A(alu__abc_42281_new_n556_), .B(alu__abc_42281_new_n560_), .Y(alu__abc_42281_new_n561_));
OR2X2 OR2X2_5059 ( .A(alu__abc_42281_new_n563_), .B(alu__abc_42281_new_n369_), .Y(alu__abc_42281_new_n564_));
OR2X2 OR2X2_506 ( .A(_abc_44694_new_n1400__bF_buf1), .B(_abc_44694_new_n2109_), .Y(_abc_44694_new_n2110_));
OR2X2 OR2X2_5060 ( .A(alu__abc_42281_new_n567_), .B(alu__abc_42281_new_n348_), .Y(alu__abc_42281_new_n568_));
OR2X2 OR2X2_5061 ( .A(alu__abc_42281_new_n566_), .B(alu__abc_42281_new_n568_), .Y(alu__abc_42281_new_n569_));
OR2X2 OR2X2_5062 ( .A(alu__abc_42281_new_n572_), .B(alu__abc_42281_new_n561_), .Y(alu__abc_42281_new_n573_));
OR2X2 OR2X2_5063 ( .A(alu_a_i_1_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n575_));
OR2X2 OR2X2_5064 ( .A(alu__abc_42281_new_n578_), .B(alu__abc_42281_new_n279_), .Y(alu__abc_42281_new_n579_));
OR2X2 OR2X2_5065 ( .A(alu__abc_42281_new_n296_), .B(alu__abc_42281_new_n301_), .Y(alu__abc_42281_new_n580_));
OR2X2 OR2X2_5066 ( .A(alu__abc_42281_new_n584_), .B(alu__abc_42281_new_n297_), .Y(alu__abc_42281_new_n585_));
OR2X2 OR2X2_5067 ( .A(alu__abc_42281_new_n582_), .B(alu__abc_42281_new_n585_), .Y(alu__abc_42281_new_n586_));
OR2X2 OR2X2_5068 ( .A(alu__abc_42281_new_n264_), .B(alu__abc_42281_new_n269_), .Y(alu__abc_42281_new_n594_));
OR2X2 OR2X2_5069 ( .A(alu__abc_42281_new_n598_), .B(alu__abc_42281_new_n258_), .Y(alu__abc_42281_new_n599_));
OR2X2 OR2X2_507 ( .A(_abc_44694_new_n2108_), .B(_abc_44694_new_n2110_), .Y(_abc_44694_new_n2111_));
OR2X2 OR2X2_5070 ( .A(alu__abc_42281_new_n596_), .B(alu__abc_42281_new_n599_), .Y(alu__abc_42281_new_n600_));
OR2X2 OR2X2_5071 ( .A(alu__abc_42281_new_n592_), .B(alu__abc_42281_new_n600_), .Y(alu__abc_42281_new_n601_));
OR2X2 OR2X2_5072 ( .A(alu__abc_42281_new_n605_), .B(alu__abc_42281_new_n573_), .Y(alu__abc_42281_new_n606_));
OR2X2 OR2X2_5073 ( .A(alu__abc_42281_new_n610_), .B(alu__abc_42281_new_n554_), .Y(alu__abc_42281_new_n611_));
OR2X2 OR2X2_5074 ( .A(alu__abc_42281_new_n615_), .B(alu__abc_42281_new_n534_), .Y(alu__abc_42281_new_n616_));
OR2X2 OR2X2_5075 ( .A(alu__abc_42281_new_n613_), .B(alu__abc_42281_new_n522_), .Y(alu__abc_42281_new_n617_));
OR2X2 OR2X2_5076 ( .A(alu__abc_42281_new_n618_), .B(alu__abc_42281_new_n518_), .Y(alu__abc_42281_new_n619_));
OR2X2 OR2X2_5077 ( .A(alu__abc_42281_new_n620_), .B(alu__abc_42281_new_n528_), .Y(alu__abc_42281_new_n621_));
OR2X2 OR2X2_5078 ( .A(alu__abc_42281_new_n625_), .B(alu__abc_42281_new_n512_), .Y(alu__abc_42281_new_n626_));
OR2X2 OR2X2_5079 ( .A(alu__abc_42281_new_n624_), .B(alu__abc_42281_new_n245_), .Y(alu__abc_42281_new_n627_));
OR2X2 OR2X2_508 ( .A(_abc_44694_new_n2112_), .B(_abc_44694_new_n1278__bF_buf0), .Y(_abc_44694_new_n2113_));
OR2X2 OR2X2_5080 ( .A(alu__abc_42281_new_n621_), .B(alu__abc_42281_new_n239_), .Y(alu__abc_42281_new_n629_));
OR2X2 OR2X2_5081 ( .A(alu__abc_42281_new_n634_), .B(alu__abc_42281_new_n230_), .Y(alu__abc_42281_new_n635_));
OR2X2 OR2X2_5082 ( .A(alu__abc_42281_new_n633_), .B(alu__abc_42281_new_n231_), .Y(alu__abc_42281_new_n636_));
OR2X2 OR2X2_5083 ( .A(alu__abc_42281_new_n619_), .B(alu__abc_42281_new_n222_), .Y(alu__abc_42281_new_n638_));
OR2X2 OR2X2_5084 ( .A(alu__abc_42281_new_n643_), .B(alu__abc_42281_new_n212_), .Y(alu__abc_42281_new_n644_));
OR2X2 OR2X2_5085 ( .A(alu__abc_42281_new_n642_), .B(alu__abc_42281_new_n213_), .Y(alu__abc_42281_new_n645_));
OR2X2 OR2X2_5086 ( .A(alu__abc_42281_new_n611_), .B(alu__abc_42281_new_n195_), .Y(alu__abc_42281_new_n649_));
OR2X2 OR2X2_5087 ( .A(alu__abc_42281_new_n609_), .B(alu__abc_42281_new_n545_), .Y(alu__abc_42281_new_n651_));
OR2X2 OR2X2_5088 ( .A(alu__abc_42281_new_n655_), .B(alu__abc_42281_new_n124_), .Y(alu__abc_42281_new_n656_));
OR2X2 OR2X2_5089 ( .A(alu__abc_42281_new_n654_), .B(alu__abc_42281_new_n125_), .Y(alu__abc_42281_new_n657_));
OR2X2 OR2X2_509 ( .A(_abc_44694_new_n2114_), .B(_abc_44694_new_n2115_), .Y(_abc_44694_new_n2116_));
OR2X2 OR2X2_5090 ( .A(alu__abc_42281_new_n659_), .B(alu__abc_42281_new_n549_), .Y(alu__abc_42281_new_n660_));
OR2X2 OR2X2_5091 ( .A(alu__abc_42281_new_n660_), .B(alu__abc_42281_new_n133_), .Y(alu__abc_42281_new_n663_));
OR2X2 OR2X2_5092 ( .A(alu__abc_42281_new_n668_), .B(alu__abc_42281_new_n187_), .Y(alu__abc_42281_new_n669_));
OR2X2 OR2X2_5093 ( .A(alu__abc_42281_new_n667_), .B(alu__abc_42281_new_n188_), .Y(alu__abc_42281_new_n670_));
OR2X2 OR2X2_5094 ( .A(alu__abc_42281_new_n651_), .B(alu__abc_42281_new_n116_), .Y(alu__abc_42281_new_n672_));
OR2X2 OR2X2_5095 ( .A(alu__abc_42281_new_n608_), .B(alu__abc_42281_new_n541_), .Y(alu__abc_42281_new_n674_));
OR2X2 OR2X2_5096 ( .A(alu__abc_42281_new_n678_), .B(alu__abc_42281_new_n159_), .Y(alu__abc_42281_new_n679_));
OR2X2 OR2X2_5097 ( .A(alu__abc_42281_new_n677_), .B(alu__abc_42281_new_n160_), .Y(alu__abc_42281_new_n680_));
OR2X2 OR2X2_5098 ( .A(alu__abc_42281_new_n674_), .B(alu__abc_42281_new_n151_), .Y(alu__abc_42281_new_n682_));
OR2X2 OR2X2_5099 ( .A(alu__abc_42281_new_n686_), .B(alu__abc_42281_new_n177_), .Y(alu__abc_42281_new_n689_));
OR2X2 OR2X2_51 ( .A(_abc_44694_new_n787_), .B(_abc_44694_new_n788_), .Y(_abc_44694_new_n789_));
OR2X2 OR2X2_510 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n2116_), .Y(_abc_44694_new_n2117_));
OR2X2 OR2X2_5100 ( .A(alu__abc_42281_new_n606_), .B(alu__abc_42281_new_n168_), .Y(alu__abc_42281_new_n691_));
OR2X2 OR2X2_5101 ( .A(alu__abc_42281_new_n283_), .B(alu__abc_42281_new_n696_), .Y(alu__abc_42281_new_n697_));
OR2X2 OR2X2_5102 ( .A(alu__abc_42281_new_n698_), .B(alu__abc_42281_new_n580_), .Y(alu__abc_42281_new_n699_));
OR2X2 OR2X2_5103 ( .A(alu__abc_42281_new_n701_), .B(alu__abc_42281_new_n702_), .Y(alu__abc_42281_new_n703_));
OR2X2 OR2X2_5104 ( .A(alu__abc_42281_new_n705_), .B(alu__abc_42281_new_n706_), .Y(alu__abc_42281_new_n707_));
OR2X2 OR2X2_5105 ( .A(alu__abc_42281_new_n708_), .B(alu__abc_42281_new_n694_), .Y(alu__abc_42281_new_n709_));
OR2X2 OR2X2_5106 ( .A(alu__abc_42281_new_n710_), .B(alu__abc_42281_new_n329_), .Y(alu__abc_42281_new_n711_));
OR2X2 OR2X2_5107 ( .A(alu__abc_42281_new_n712_), .B(alu__abc_42281_new_n337_), .Y(alu__abc_42281_new_n713_));
OR2X2 OR2X2_5108 ( .A(alu__abc_42281_new_n714_), .B(alu__abc_42281_new_n569_), .Y(alu__abc_42281_new_n715_));
OR2X2 OR2X2_5109 ( .A(alu__abc_42281_new_n716_), .B(alu__abc_42281_new_n558_), .Y(alu__abc_42281_new_n717_));
OR2X2 OR2X2_511 ( .A(_abc_44694_new_n2119_), .B(_abc_44694_new_n2080_), .Y(_abc_44694_new_n2120_));
OR2X2 OR2X2_5110 ( .A(alu__abc_42281_new_n718_), .B(alu__abc_42281_new_n322_), .Y(alu__abc_42281_new_n719_));
OR2X2 OR2X2_5111 ( .A(alu__abc_42281_new_n719_), .B(alu__abc_42281_new_n336_), .Y(alu__abc_42281_new_n720_));
OR2X2 OR2X2_5112 ( .A(alu__abc_42281_new_n725_), .B(alu__abc_42281_new_n371_), .Y(alu__abc_42281_new_n726_));
OR2X2 OR2X2_5113 ( .A(alu__abc_42281_new_n724_), .B(alu__abc_42281_new_n372_), .Y(alu__abc_42281_new_n727_));
OR2X2 OR2X2_5114 ( .A(alu__abc_42281_new_n729_), .B(alu__abc_42281_new_n722_), .Y(alu__abc_42281_new_n730_));
OR2X2 OR2X2_5115 ( .A(alu__abc_42281_new_n732_), .B(alu__abc_42281_new_n595_), .Y(alu__abc_42281_new_n733_));
OR2X2 OR2X2_5116 ( .A(alu__abc_42281_new_n737_), .B(alu__abc_42281_new_n587_), .Y(alu__abc_42281_new_n738_));
OR2X2 OR2X2_5117 ( .A(alu__abc_42281_new_n736_), .B(alu__abc_42281_new_n262_), .Y(alu__abc_42281_new_n739_));
OR2X2 OR2X2_5118 ( .A(alu__abc_42281_new_n733_), .B(alu__abc_42281_new_n256_), .Y(alu__abc_42281_new_n741_));
OR2X2 OR2X2_5119 ( .A(alu__abc_42281_new_n746_), .B(alu__abc_42281_new_n589_), .Y(alu__abc_42281_new_n747_));
OR2X2 OR2X2_512 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_20_), .Y(_abc_44694_new_n2121_));
OR2X2 OR2X2_5120 ( .A(alu__abc_42281_new_n745_), .B(alu__abc_42281_new_n268_), .Y(alu__abc_42281_new_n748_));
OR2X2 OR2X2_5121 ( .A(alu__abc_42281_new_n752_), .B(alu__abc_42281_new_n292_), .Y(alu__abc_42281_new_n753_));
OR2X2 OR2X2_5122 ( .A(alu__abc_42281_new_n753_), .B(alu__abc_42281_new_n750_), .Y(alu__abc_42281_new_n754_));
OR2X2 OR2X2_5123 ( .A(alu__abc_42281_new_n755_), .B(alu__abc_42281_new_n301_), .Y(alu__abc_42281_new_n756_));
OR2X2 OR2X2_5124 ( .A(alu__abc_42281_new_n763_), .B(alu__abc_42281_new_n752_), .Y(alu__abc_42281_new_n764_));
OR2X2 OR2X2_5125 ( .A(alu__abc_42281_new_n586_), .B(alu__abc_42281_new_n275_), .Y(alu__abc_42281_new_n768_));
OR2X2 OR2X2_5126 ( .A(alu__abc_42281_new_n776_), .B(alu__abc_42281_new_n305_), .Y(alu__abc_42281_new_n777_));
OR2X2 OR2X2_5127 ( .A(alu__abc_42281_new_n777_), .B(alu__abc_42281_new_n319_), .Y(alu__abc_42281_new_n778_));
OR2X2 OR2X2_5128 ( .A(alu__abc_42281_new_n708_), .B(alu__abc_42281_new_n312_), .Y(alu__abc_42281_new_n779_));
OR2X2 OR2X2_5129 ( .A(alu__abc_42281_new_n780_), .B(alu__abc_42281_new_n320_), .Y(alu__abc_42281_new_n781_));
OR2X2 OR2X2_513 ( .A(_abc_44694_new_n2076_), .B(pc_q_21_), .Y(_abc_44694_new_n2124_));
OR2X2 OR2X2_5130 ( .A(alu__abc_42281_new_n705_), .B(alu__abc_42281_new_n783_), .Y(alu__abc_42281_new_n784_));
OR2X2 OR2X2_5131 ( .A(alu__abc_42281_new_n785_), .B(alu__abc_42281_new_n347_), .Y(alu__abc_42281_new_n786_));
OR2X2 OR2X2_5132 ( .A(alu__abc_42281_new_n787_), .B(alu__abc_42281_new_n565_), .Y(alu__abc_42281_new_n788_));
OR2X2 OR2X2_5133 ( .A(alu__abc_42281_new_n788_), .B(alu__abc_42281_new_n346_), .Y(alu__abc_42281_new_n789_));
OR2X2 OR2X2_5134 ( .A(alu__abc_42281_new_n715_), .B(alu__abc_42281_new_n311_), .Y(alu__abc_42281_new_n791_));
OR2X2 OR2X2_5135 ( .A(alu__abc_42281_new_n795_), .B(alu__abc_42281_new_n340_), .Y(alu__abc_42281_new_n796_));
OR2X2 OR2X2_5136 ( .A(alu__abc_42281_new_n796_), .B(alu__abc_42281_new_n354_), .Y(alu__abc_42281_new_n797_));
OR2X2 OR2X2_5137 ( .A(alu__abc_42281_new_n798_), .B(alu__abc_42281_new_n355_), .Y(alu__abc_42281_new_n799_));
OR2X2 OR2X2_5138 ( .A(alu__abc_42281_new_n717_), .B(alu__abc_42281_new_n328_), .Y(alu__abc_42281_new_n801_));
OR2X2 OR2X2_5139 ( .A(alu__abc_42281_new_n617_), .B(alu__abc_42281_new_n204_), .Y(alu__abc_42281_new_n814_));
OR2X2 OR2X2_514 ( .A(_abc_44694_new_n2128_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n2129_));
OR2X2 OR2X2_5140 ( .A(alu__abc_42281_new_n817_), .B(alu__abc_42281_new_n141_), .Y(alu__abc_42281_new_n818_));
OR2X2 OR2X2_5141 ( .A(alu__abc_42281_new_n816_), .B(alu__abc_42281_new_n142_), .Y(alu__abc_42281_new_n819_));
OR2X2 OR2X2_5142 ( .A(alu__abc_42281_new_n827_), .B(alu__abc_42281_new_n616_), .Y(alu__abc_42281_new_n828_));
OR2X2 OR2X2_5143 ( .A(alu_a_i_8_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n830_));
OR2X2 OR2X2_5144 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_9_), .Y(alu__abc_42281_new_n831_));
OR2X2 OR2X2_5145 ( .A(alu__abc_42281_new_n832_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n833_));
OR2X2 OR2X2_5146 ( .A(alu_a_i_10_), .B(alu_b_i_0_bF_buf0_), .Y(alu__abc_42281_new_n834_));
OR2X2 OR2X2_5147 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_11_), .Y(alu__abc_42281_new_n835_));
OR2X2 OR2X2_5148 ( .A(alu__abc_42281_new_n836_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n837_));
OR2X2 OR2X2_5149 ( .A(alu__abc_42281_new_n838_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n839_));
OR2X2 OR2X2_515 ( .A(_abc_44694_new_n2127_), .B(_abc_44694_new_n1399__bF_buf4), .Y(_abc_44694_new_n2130_));
OR2X2 OR2X2_5150 ( .A(alu_a_i_12_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n840_));
OR2X2 OR2X2_5151 ( .A(alu__abc_42281_new_n288__bF_buf0), .B(alu_a_i_13_), .Y(alu__abc_42281_new_n841_));
OR2X2 OR2X2_5152 ( .A(alu__abc_42281_new_n842_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n843_));
OR2X2 OR2X2_5153 ( .A(alu_a_i_14_), .B(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n844_));
OR2X2 OR2X2_5154 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_15_), .Y(alu__abc_42281_new_n845_));
OR2X2 OR2X2_5155 ( .A(alu__abc_42281_new_n846_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n847_));
OR2X2 OR2X2_5156 ( .A(alu__abc_42281_new_n848_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n849_));
OR2X2 OR2X2_5157 ( .A(alu__abc_42281_new_n850_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n851_));
OR2X2 OR2X2_5158 ( .A(alu_a_i_4_), .B(alu_b_i_0_bF_buf2_), .Y(alu__abc_42281_new_n852_));
OR2X2 OR2X2_5159 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu_a_i_5_), .Y(alu__abc_42281_new_n853_));
OR2X2 OR2X2_516 ( .A(pc_q_21_), .B(REGFILE_SIM_reg_bank_ra_i_3_), .Y(_abc_44694_new_n2132_));
OR2X2 OR2X2_5160 ( .A(alu__abc_42281_new_n854_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n855_));
OR2X2 OR2X2_5161 ( .A(alu_a_i_6_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n856_));
OR2X2 OR2X2_5162 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_7_), .Y(alu__abc_42281_new_n857_));
OR2X2 OR2X2_5163 ( .A(alu__abc_42281_new_n858_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n859_));
OR2X2 OR2X2_5164 ( .A(alu_a_i_2_), .B(alu_b_i_0_bF_buf0_), .Y(alu__abc_42281_new_n862_));
OR2X2 OR2X2_5165 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_3_), .Y(alu__abc_42281_new_n863_));
OR2X2 OR2X2_5166 ( .A(alu__abc_42281_new_n288__bF_buf0), .B(alu_a_i_1_), .Y(alu__abc_42281_new_n866_));
OR2X2 OR2X2_5167 ( .A(alu__abc_42281_new_n868_), .B(alu__abc_42281_new_n865_), .Y(alu__abc_42281_new_n869_));
OR2X2 OR2X2_5168 ( .A(alu__abc_42281_new_n870_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n871_));
OR2X2 OR2X2_5169 ( .A(alu__abc_42281_new_n871_), .B(alu__abc_42281_new_n861_), .Y(alu__abc_42281_new_n872_));
OR2X2 OR2X2_517 ( .A(_abc_44694_new_n2135_), .B(_abc_44694_new_n2099_), .Y(_abc_44694_new_n2136_));
OR2X2 OR2X2_5170 ( .A(alu__abc_42281_new_n873_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n874_));
OR2X2 OR2X2_5171 ( .A(alu_a_i_24_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n877_));
OR2X2 OR2X2_5172 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_25_), .Y(alu__abc_42281_new_n878_));
OR2X2 OR2X2_5173 ( .A(alu__abc_42281_new_n879_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n880_));
OR2X2 OR2X2_5174 ( .A(alu_a_i_26_), .B(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n881_));
OR2X2 OR2X2_5175 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu_a_i_27_), .Y(alu__abc_42281_new_n882_));
OR2X2 OR2X2_5176 ( .A(alu__abc_42281_new_n883_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n884_));
OR2X2 OR2X2_5177 ( .A(alu__abc_42281_new_n885_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n886_));
OR2X2 OR2X2_5178 ( .A(alu_a_i_28_), .B(alu_b_i_0_bF_buf2_), .Y(alu__abc_42281_new_n887_));
OR2X2 OR2X2_5179 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_29_), .Y(alu__abc_42281_new_n888_));
OR2X2 OR2X2_518 ( .A(_abc_44694_new_n2102_), .B(_abc_44694_new_n2136_), .Y(_abc_44694_new_n2137_));
OR2X2 OR2X2_5180 ( .A(alu__abc_42281_new_n889_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n890_));
OR2X2 OR2X2_5181 ( .A(alu_a_i_30_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n891_));
OR2X2 OR2X2_5182 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_31_), .Y(alu__abc_42281_new_n892_));
OR2X2 OR2X2_5183 ( .A(alu__abc_42281_new_n893_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n894_));
OR2X2 OR2X2_5184 ( .A(alu__abc_42281_new_n895_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n896_));
OR2X2 OR2X2_5185 ( .A(alu__abc_42281_new_n897_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n898_));
OR2X2 OR2X2_5186 ( .A(alu_a_i_16_), .B(alu_b_i_0_bF_buf0_), .Y(alu__abc_42281_new_n899_));
OR2X2 OR2X2_5187 ( .A(alu__abc_42281_new_n288__bF_buf0), .B(alu_a_i_17_), .Y(alu__abc_42281_new_n900_));
OR2X2 OR2X2_5188 ( .A(alu__abc_42281_new_n901_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n902_));
OR2X2 OR2X2_5189 ( .A(alu_a_i_18_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n903_));
OR2X2 OR2X2_519 ( .A(_abc_44694_new_n2145_), .B(_abc_44694_new_n2131_), .Y(_abc_44694_new_n2146_));
OR2X2 OR2X2_5190 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_19_), .Y(alu__abc_42281_new_n904_));
OR2X2 OR2X2_5191 ( .A(alu__abc_42281_new_n905_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n906_));
OR2X2 OR2X2_5192 ( .A(alu__abc_42281_new_n907_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n908_));
OR2X2 OR2X2_5193 ( .A(alu_a_i_20_), .B(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n909_));
OR2X2 OR2X2_5194 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu_a_i_21_), .Y(alu__abc_42281_new_n910_));
OR2X2 OR2X2_5195 ( .A(alu__abc_42281_new_n911_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n912_));
OR2X2 OR2X2_5196 ( .A(alu_a_i_22_), .B(alu_b_i_0_bF_buf2_), .Y(alu__abc_42281_new_n913_));
OR2X2 OR2X2_5197 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_23_), .Y(alu__abc_42281_new_n914_));
OR2X2 OR2X2_5198 ( .A(alu__abc_42281_new_n915_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n916_));
OR2X2 OR2X2_5199 ( .A(alu__abc_42281_new_n917_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n918_));
OR2X2 OR2X2_52 ( .A(_abc_44694_new_n789_), .B(_abc_44694_new_n786_), .Y(_abc_44694_new_n790_));
OR2X2 OR2X2_520 ( .A(_abc_44694_new_n1400__bF_buf0), .B(_abc_44694_new_n2148_), .Y(_abc_44694_new_n2149_));
OR2X2 OR2X2_5200 ( .A(alu__abc_42281_new_n919_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n920_));
OR2X2 OR2X2_5201 ( .A(alu__abc_42281_new_n921_), .B(alu__abc_42281_new_n271__bF_buf2), .Y(alu__abc_42281_new_n922_));
OR2X2 OR2X2_5202 ( .A(alu__abc_42281_new_n927_), .B(alu__abc_42281_new_n929_), .Y(alu__abc_42281_new_n930_));
OR2X2 OR2X2_5203 ( .A(alu__abc_42281_new_n941__bF_buf4), .B(alu__abc_42281_new_n942__bF_buf4), .Y(alu__abc_42281_new_n943_));
OR2X2 OR2X2_5204 ( .A(alu__abc_42281_new_n944_), .B(alu__abc_42281_new_n940_), .Y(alu__abc_42281_new_n945_));
OR2X2 OR2X2_5205 ( .A(alu__abc_42281_new_n945_), .B(alu__abc_42281_new_n937_), .Y(alu__abc_42281_new_n946_));
OR2X2 OR2X2_5206 ( .A(alu_op_i_1_), .B(alu_op_i_2_), .Y(alu__abc_42281_new_n947_));
OR2X2 OR2X2_5207 ( .A(alu__abc_42281_new_n949_), .B(alu__abc_42281_new_n948_), .Y(alu__abc_42281_new_n950_));
OR2X2 OR2X2_5208 ( .A(alu__abc_42281_new_n760_), .B(alu_c_i), .Y(alu__abc_42281_new_n954_));
OR2X2 OR2X2_5209 ( .A(alu__abc_42281_new_n956_), .B(alu__abc_42281_new_n951_), .Y(alu__abc_42281_new_n957_));
OR2X2 OR2X2_521 ( .A(_abc_44694_new_n2147_), .B(_abc_44694_new_n2149_), .Y(_abc_44694_new_n2150_));
OR2X2 OR2X2_5210 ( .A(alu__abc_42281_new_n957_), .B(alu__abc_42281_new_n946_), .Y(alu__abc_42281_new_n958_));
OR2X2 OR2X2_5211 ( .A(alu__abc_42281_new_n958_), .B(alu__abc_42281_new_n930_), .Y(alu__abc_42281_new_n959_));
OR2X2 OR2X2_5212 ( .A(alu__abc_42281_new_n924_), .B(alu__abc_42281_new_n959_), .Y(alu_p_o_0_));
OR2X2 OR2X2_5213 ( .A(alu__abc_42281_new_n962_), .B(alu__abc_42281_new_n963_), .Y(alu__abc_42281_new_n964_));
OR2X2 OR2X2_5214 ( .A(alu__abc_42281_new_n967_), .B(alu__abc_42281_new_n966_), .Y(alu__abc_42281_new_n968_));
OR2X2 OR2X2_5215 ( .A(alu__abc_42281_new_n965_), .B(alu__abc_42281_new_n969_), .Y(alu__abc_42281_new_n970_));
OR2X2 OR2X2_5216 ( .A(alu_a_i_25_), .B(alu_b_i_0_bF_buf0_), .Y(alu__abc_42281_new_n972_));
OR2X2 OR2X2_5217 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_26_), .Y(alu__abc_42281_new_n973_));
OR2X2 OR2X2_5218 ( .A(alu__abc_42281_new_n974_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n975_));
OR2X2 OR2X2_5219 ( .A(alu_a_i_27_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n976_));
OR2X2 OR2X2_522 ( .A(_abc_44694_new_n2151_), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n2152_));
OR2X2 OR2X2_5220 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu_a_i_28_), .Y(alu__abc_42281_new_n977_));
OR2X2 OR2X2_5221 ( .A(alu__abc_42281_new_n978_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n979_));
OR2X2 OR2X2_5222 ( .A(alu__abc_42281_new_n971_), .B(alu__abc_42281_new_n981_), .Y(alu__abc_42281_new_n982_));
OR2X2 OR2X2_5223 ( .A(alu_a_i_17_), .B(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n984_));
OR2X2 OR2X2_5224 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_18_), .Y(alu__abc_42281_new_n985_));
OR2X2 OR2X2_5225 ( .A(alu__abc_42281_new_n986_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n987_));
OR2X2 OR2X2_5226 ( .A(alu_a_i_19_), .B(alu_b_i_0_bF_buf2_), .Y(alu__abc_42281_new_n988_));
OR2X2 OR2X2_5227 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_20_), .Y(alu__abc_42281_new_n989_));
OR2X2 OR2X2_5228 ( .A(alu__abc_42281_new_n990_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n991_));
OR2X2 OR2X2_5229 ( .A(alu__abc_42281_new_n992_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n993_));
OR2X2 OR2X2_523 ( .A(_abc_44694_new_n2153_), .B(_abc_44694_new_n2154_), .Y(_abc_44694_new_n2155_));
OR2X2 OR2X2_5230 ( .A(alu_a_i_21_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n994_));
OR2X2 OR2X2_5231 ( .A(alu__abc_42281_new_n288__bF_buf0), .B(alu_a_i_22_), .Y(alu__abc_42281_new_n995_));
OR2X2 OR2X2_5232 ( .A(alu__abc_42281_new_n996_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n997_));
OR2X2 OR2X2_5233 ( .A(alu_a_i_23_), .B(alu_b_i_0_bF_buf0_), .Y(alu__abc_42281_new_n998_));
OR2X2 OR2X2_5234 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_24_), .Y(alu__abc_42281_new_n999_));
OR2X2 OR2X2_5235 ( .A(alu__abc_42281_new_n1000_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n1001_));
OR2X2 OR2X2_5236 ( .A(alu__abc_42281_new_n1002_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1003_));
OR2X2 OR2X2_5237 ( .A(alu__abc_42281_new_n983_), .B(alu__abc_42281_new_n1005_), .Y(alu__abc_42281_new_n1006_));
OR2X2 OR2X2_5238 ( .A(alu__abc_42281_new_n1006_), .B(alu__abc_42281_new_n271__bF_buf0), .Y(alu__abc_42281_new_n1007_));
OR2X2 OR2X2_5239 ( .A(alu_a_i_3_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n1008_));
OR2X2 OR2X2_524 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n2155_), .Y(_abc_44694_new_n2156_));
OR2X2 OR2X2_5240 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu_a_i_4_), .Y(alu__abc_42281_new_n1009_));
OR2X2 OR2X2_5241 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_2_), .Y(alu__abc_42281_new_n1012_));
OR2X2 OR2X2_5242 ( .A(alu_a_i_1_), .B(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n1013_));
OR2X2 OR2X2_5243 ( .A(alu__abc_42281_new_n1011_), .B(alu__abc_42281_new_n1015_), .Y(alu__abc_42281_new_n1016_));
OR2X2 OR2X2_5244 ( .A(alu__abc_42281_new_n1016_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1017_));
OR2X2 OR2X2_5245 ( .A(alu_a_i_5_), .B(alu_b_i_0_bF_buf2_), .Y(alu__abc_42281_new_n1018_));
OR2X2 OR2X2_5246 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_6_), .Y(alu__abc_42281_new_n1019_));
OR2X2 OR2X2_5247 ( .A(alu__abc_42281_new_n1020_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n1021_));
OR2X2 OR2X2_5248 ( .A(alu_a_i_7_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n1022_));
OR2X2 OR2X2_5249 ( .A(alu__abc_42281_new_n288__bF_buf0), .B(alu_a_i_8_), .Y(alu__abc_42281_new_n1023_));
OR2X2 OR2X2_525 ( .A(_abc_44694_new_n2158_), .B(_abc_44694_new_n2129_), .Y(_abc_44694_new_n2159_));
OR2X2 OR2X2_5250 ( .A(alu__abc_42281_new_n1024_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n1025_));
OR2X2 OR2X2_5251 ( .A(alu__abc_42281_new_n1026_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1027_));
OR2X2 OR2X2_5252 ( .A(alu__abc_42281_new_n1028_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n1029_));
OR2X2 OR2X2_5253 ( .A(alu_a_i_9_), .B(alu_b_i_0_bF_buf0_), .Y(alu__abc_42281_new_n1030_));
OR2X2 OR2X2_5254 ( .A(alu__abc_42281_new_n288__bF_buf4), .B(alu_a_i_10_), .Y(alu__abc_42281_new_n1031_));
OR2X2 OR2X2_5255 ( .A(alu__abc_42281_new_n1032_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n1033_));
OR2X2 OR2X2_5256 ( .A(alu_a_i_11_), .B(alu_b_i_0_bF_buf4_), .Y(alu__abc_42281_new_n1034_));
OR2X2 OR2X2_5257 ( .A(alu__abc_42281_new_n288__bF_buf3), .B(alu_a_i_12_), .Y(alu__abc_42281_new_n1035_));
OR2X2 OR2X2_5258 ( .A(alu__abc_42281_new_n1036_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n1037_));
OR2X2 OR2X2_5259 ( .A(alu__abc_42281_new_n1038_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n1039_));
OR2X2 OR2X2_526 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_21_), .Y(_abc_44694_new_n2160_));
OR2X2 OR2X2_5260 ( .A(alu_a_i_13_), .B(alu_b_i_0_bF_buf3_), .Y(alu__abc_42281_new_n1040_));
OR2X2 OR2X2_5261 ( .A(alu__abc_42281_new_n288__bF_buf2), .B(alu_a_i_14_), .Y(alu__abc_42281_new_n1041_));
OR2X2 OR2X2_5262 ( .A(alu__abc_42281_new_n1042_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n1043_));
OR2X2 OR2X2_5263 ( .A(alu_a_i_15_), .B(alu_b_i_0_bF_buf2_), .Y(alu__abc_42281_new_n1044_));
OR2X2 OR2X2_5264 ( .A(alu__abc_42281_new_n288__bF_buf1), .B(alu_a_i_16_), .Y(alu__abc_42281_new_n1045_));
OR2X2 OR2X2_5265 ( .A(alu__abc_42281_new_n1046_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n1047_));
OR2X2 OR2X2_5266 ( .A(alu__abc_42281_new_n1048_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n1049_));
OR2X2 OR2X2_5267 ( .A(alu__abc_42281_new_n1050_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n1051_));
OR2X2 OR2X2_5268 ( .A(alu__abc_42281_new_n1052_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n1053_));
OR2X2 OR2X2_5269 ( .A(alu__abc_42281_new_n283_), .B(alu__abc_42281_new_n286_), .Y(alu__abc_42281_new_n1056_));
OR2X2 OR2X2_527 ( .A(_abc_44694_new_n2125_), .B(pc_q_22_), .Y(_abc_44694_new_n2163_));
OR2X2 OR2X2_5270 ( .A(alu__abc_42281_new_n576_), .B(alu__abc_42281_new_n577_), .Y(alu__abc_42281_new_n1060_));
OR2X2 OR2X2_5271 ( .A(alu__abc_42281_new_n1064_), .B(alu__abc_42281_new_n1063_), .Y(alu__abc_42281_new_n1065_));
OR2X2 OR2X2_5272 ( .A(alu__abc_42281_new_n1062_), .B(alu__abc_42281_new_n1065_), .Y(alu__abc_42281_new_n1066_));
OR2X2 OR2X2_5273 ( .A(alu__abc_42281_new_n1066_), .B(alu__abc_42281_new_n1059_), .Y(alu__abc_42281_new_n1067_));
OR2X2 OR2X2_5274 ( .A(alu__abc_42281_new_n1061_), .B(alu__abc_42281_new_n761_), .Y(alu__abc_42281_new_n1068_));
OR2X2 OR2X2_5275 ( .A(alu__abc_42281_new_n1076_), .B(alu__abc_42281_new_n1077_), .Y(alu__abc_42281_new_n1078_));
OR2X2 OR2X2_5276 ( .A(alu__abc_42281_new_n1075_), .B(alu__abc_42281_new_n1078_), .Y(alu__abc_42281_new_n1079_));
OR2X2 OR2X2_5277 ( .A(alu__abc_42281_new_n1071_), .B(alu__abc_42281_new_n1079_), .Y(alu__abc_42281_new_n1080_));
OR2X2 OR2X2_5278 ( .A(alu__abc_42281_new_n1080_), .B(alu__abc_42281_new_n1067_), .Y(alu__abc_42281_new_n1081_));
OR2X2 OR2X2_5279 ( .A(alu__abc_42281_new_n1055_), .B(alu__abc_42281_new_n1081_), .Y(alu_p_o_1_));
OR2X2 OR2X2_528 ( .A(_abc_44694_new_n2167_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n2168_));
OR2X2 OR2X2_5280 ( .A(alu__abc_42281_new_n893_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n1083_));
OR2X2 OR2X2_5281 ( .A(alu__abc_42281_new_n962_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n1084_));
OR2X2 OR2X2_5282 ( .A(alu__abc_42281_new_n883_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n1087_));
OR2X2 OR2X2_5283 ( .A(alu__abc_42281_new_n889_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n1088_));
OR2X2 OR2X2_5284 ( .A(alu__abc_42281_new_n1086_), .B(alu__abc_42281_new_n1090_), .Y(alu__abc_42281_new_n1091_));
OR2X2 OR2X2_5285 ( .A(alu__abc_42281_new_n905_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n1093_));
OR2X2 OR2X2_5286 ( .A(alu__abc_42281_new_n911_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n1094_));
OR2X2 OR2X2_5287 ( .A(alu__abc_42281_new_n1095_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n1096_));
OR2X2 OR2X2_5288 ( .A(alu__abc_42281_new_n915_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n1097_));
OR2X2 OR2X2_5289 ( .A(alu__abc_42281_new_n879_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n1098_));
OR2X2 OR2X2_529 ( .A(_abc_44694_new_n2166_), .B(_abc_44694_new_n1399__bF_buf3), .Y(_abc_44694_new_n2169_));
OR2X2 OR2X2_5290 ( .A(alu__abc_42281_new_n1099_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n1100_));
OR2X2 OR2X2_5291 ( .A(alu__abc_42281_new_n1092_), .B(alu__abc_42281_new_n1102_), .Y(alu__abc_42281_new_n1103_));
OR2X2 OR2X2_5292 ( .A(alu__abc_42281_new_n1103_), .B(alu__abc_42281_new_n271__bF_buf4), .Y(alu__abc_42281_new_n1104_));
OR2X2 OR2X2_5293 ( .A(alu__abc_42281_new_n1106_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n1107_));
OR2X2 OR2X2_5294 ( .A(alu__abc_42281_new_n1107_), .B(alu__abc_42281_new_n1105_), .Y(alu__abc_42281_new_n1108_));
OR2X2 OR2X2_5295 ( .A(alu__abc_42281_new_n858_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n1109_));
OR2X2 OR2X2_5296 ( .A(alu__abc_42281_new_n832_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n1110_));
OR2X2 OR2X2_5297 ( .A(alu__abc_42281_new_n1111_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n1112_));
OR2X2 OR2X2_5298 ( .A(alu__abc_42281_new_n836_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n1115_));
OR2X2 OR2X2_5299 ( .A(alu__abc_42281_new_n842_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n1116_));
OR2X2 OR2X2_53 ( .A(_abc_44694_new_n673__bF_buf3), .B(_abc_44694_new_n790_), .Y(_abc_44694_new_n791_));
OR2X2 OR2X2_530 ( .A(pc_q_22_), .B(REGFILE_SIM_reg_bank_ra_i_4_bF_buf3_), .Y(_abc_44694_new_n2174_));
OR2X2 OR2X2_5300 ( .A(alu__abc_42281_new_n1117_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n1118_));
OR2X2 OR2X2_5301 ( .A(alu__abc_42281_new_n846_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n1119_));
OR2X2 OR2X2_5302 ( .A(alu__abc_42281_new_n901_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n1120_));
OR2X2 OR2X2_5303 ( .A(alu__abc_42281_new_n1121_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1122_));
OR2X2 OR2X2_5304 ( .A(alu__abc_42281_new_n1124_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n1125_));
OR2X2 OR2X2_5305 ( .A(alu__abc_42281_new_n1125_), .B(alu__abc_42281_new_n1114_), .Y(alu__abc_42281_new_n1126_));
OR2X2 OR2X2_5306 ( .A(alu__abc_42281_new_n765_), .B(alu__abc_42281_new_n762_), .Y(alu__abc_42281_new_n1130_));
OR2X2 OR2X2_5307 ( .A(alu__abc_42281_new_n1133_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n1134_));
OR2X2 OR2X2_5308 ( .A(alu__abc_42281_new_n1144_), .B(alu__abc_42281_new_n1145_), .Y(alu__abc_42281_new_n1146_));
OR2X2 OR2X2_5309 ( .A(alu__abc_42281_new_n1146_), .B(alu__abc_42281_new_n1143_), .Y(alu__abc_42281_new_n1147_));
OR2X2 OR2X2_531 ( .A(_abc_44694_new_n2173_), .B(_abc_44694_new_n2177_), .Y(_abc_44694_new_n2180_));
OR2X2 OR2X2_5310 ( .A(alu__abc_42281_new_n1147_), .B(alu__abc_42281_new_n1141_), .Y(alu__abc_42281_new_n1148_));
OR2X2 OR2X2_5311 ( .A(alu__abc_42281_new_n1140_), .B(alu__abc_42281_new_n1148_), .Y(alu__abc_42281_new_n1149_));
OR2X2 OR2X2_5312 ( .A(alu__abc_42281_new_n401_), .B(alu__abc_42281_new_n296_), .Y(alu__abc_42281_new_n1151_));
OR2X2 OR2X2_5313 ( .A(alu__abc_42281_new_n1150_), .B(alu__abc_42281_new_n1154_), .Y(alu__abc_42281_new_n1155_));
OR2X2 OR2X2_5314 ( .A(alu__abc_42281_new_n1155_), .B(alu__abc_42281_new_n1149_), .Y(alu__abc_42281_new_n1156_));
OR2X2 OR2X2_5315 ( .A(alu__abc_42281_new_n1132_), .B(alu__abc_42281_new_n1156_), .Y(alu__abc_42281_new_n1157_));
OR2X2 OR2X2_5316 ( .A(alu__abc_42281_new_n1157_), .B(alu__abc_42281_new_n1128_), .Y(alu_p_o_2_));
OR2X2 OR2X2_5317 ( .A(alu__abc_42281_new_n978_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n1161_));
OR2X2 OR2X2_5318 ( .A(alu__abc_42281_new_n968_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n1162_));
OR2X2 OR2X2_5319 ( .A(alu__abc_42281_new_n1160_), .B(alu__abc_42281_new_n1164_), .Y(alu__abc_42281_new_n1165_));
OR2X2 OR2X2_532 ( .A(_abc_44694_new_n2182_), .B(_abc_44694_new_n2170_), .Y(_abc_44694_new_n2183_));
OR2X2 OR2X2_5320 ( .A(alu__abc_42281_new_n990_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n1167_));
OR2X2 OR2X2_5321 ( .A(alu__abc_42281_new_n996_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n1168_));
OR2X2 OR2X2_5322 ( .A(alu__abc_42281_new_n1169_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1170_));
OR2X2 OR2X2_5323 ( .A(alu__abc_42281_new_n1000_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n1171_));
OR2X2 OR2X2_5324 ( .A(alu__abc_42281_new_n974_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n1172_));
OR2X2 OR2X2_5325 ( .A(alu__abc_42281_new_n1173_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n1174_));
OR2X2 OR2X2_5326 ( .A(alu__abc_42281_new_n1166_), .B(alu__abc_42281_new_n1176_), .Y(alu__abc_42281_new_n1177_));
OR2X2 OR2X2_5327 ( .A(alu__abc_42281_new_n1177_), .B(alu__abc_42281_new_n271__bF_buf3), .Y(alu__abc_42281_new_n1178_));
OR2X2 OR2X2_5328 ( .A(alu__abc_42281_new_n1180_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n1181_));
OR2X2 OR2X2_5329 ( .A(alu__abc_42281_new_n1181_), .B(alu__abc_42281_new_n1179_), .Y(alu__abc_42281_new_n1182_));
OR2X2 OR2X2_533 ( .A(_abc_44694_new_n1400__bF_buf4), .B(_abc_44694_new_n2185_), .Y(_abc_44694_new_n2186_));
OR2X2 OR2X2_5330 ( .A(alu__abc_42281_new_n1024_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n1183_));
OR2X2 OR2X2_5331 ( .A(alu__abc_42281_new_n1032_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n1184_));
OR2X2 OR2X2_5332 ( .A(alu__abc_42281_new_n1185_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n1186_));
OR2X2 OR2X2_5333 ( .A(alu__abc_42281_new_n1036_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n1189_));
OR2X2 OR2X2_5334 ( .A(alu__abc_42281_new_n1042_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n1190_));
OR2X2 OR2X2_5335 ( .A(alu__abc_42281_new_n1191_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n1192_));
OR2X2 OR2X2_5336 ( .A(alu__abc_42281_new_n1046_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n1193_));
OR2X2 OR2X2_5337 ( .A(alu__abc_42281_new_n986_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n1194_));
OR2X2 OR2X2_5338 ( .A(alu__abc_42281_new_n1195_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n1196_));
OR2X2 OR2X2_5339 ( .A(alu__abc_42281_new_n1198_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n1199_));
OR2X2 OR2X2_534 ( .A(_abc_44694_new_n2184_), .B(_abc_44694_new_n2186_), .Y(_abc_44694_new_n2187_));
OR2X2 OR2X2_5340 ( .A(alu__abc_42281_new_n1199_), .B(alu__abc_42281_new_n1188_), .Y(alu__abc_42281_new_n1200_));
OR2X2 OR2X2_5341 ( .A(alu__abc_42281_new_n757_), .B(alu__abc_42281_new_n766_), .Y(alu__abc_42281_new_n1203_));
OR2X2 OR2X2_5342 ( .A(alu__abc_42281_new_n1208_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n1209_));
OR2X2 OR2X2_5343 ( .A(alu__abc_42281_new_n1210_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n1211_));
OR2X2 OR2X2_5344 ( .A(alu__abc_42281_new_n1218_), .B(alu__abc_42281_new_n1217_), .Y(alu__abc_42281_new_n1219_));
OR2X2 OR2X2_5345 ( .A(alu__abc_42281_new_n1219_), .B(alu__abc_42281_new_n1216_), .Y(alu__abc_42281_new_n1220_));
OR2X2 OR2X2_5346 ( .A(alu__abc_42281_new_n1215_), .B(alu__abc_42281_new_n1220_), .Y(alu__abc_42281_new_n1221_));
OR2X2 OR2X2_5347 ( .A(alu__abc_42281_new_n1207_), .B(alu__abc_42281_new_n1221_), .Y(alu__abc_42281_new_n1222_));
OR2X2 OR2X2_5348 ( .A(alu__abc_42281_new_n1224_), .B(alu__abc_42281_new_n750_), .Y(alu__abc_42281_new_n1225_));
OR2X2 OR2X2_5349 ( .A(alu__abc_42281_new_n403_), .B(alu__abc_42281_new_n301_), .Y(alu__abc_42281_new_n1226_));
OR2X2 OR2X2_535 ( .A(_abc_44694_new_n2188_), .B(_abc_44694_new_n1278__bF_buf4), .Y(_abc_44694_new_n2189_));
OR2X2 OR2X2_5350 ( .A(alu__abc_42281_new_n1228_), .B(alu__abc_42281_new_n1223_), .Y(alu__abc_42281_new_n1229_));
OR2X2 OR2X2_5351 ( .A(alu__abc_42281_new_n1222_), .B(alu__abc_42281_new_n1229_), .Y(alu__abc_42281_new_n1230_));
OR2X2 OR2X2_5352 ( .A(alu__abc_42281_new_n1206_), .B(alu__abc_42281_new_n1230_), .Y(alu__abc_42281_new_n1231_));
OR2X2 OR2X2_5353 ( .A(alu__abc_42281_new_n1231_), .B(alu__abc_42281_new_n1202_), .Y(alu_p_o_3_));
OR2X2 OR2X2_5354 ( .A(alu__abc_42281_new_n767_), .B(alu__abc_42281_new_n769_), .Y(alu__abc_42281_new_n1234_));
OR2X2 OR2X2_5355 ( .A(alu__abc_42281_new_n405_), .B(alu__abc_42281_new_n276_), .Y(alu__abc_42281_new_n1237_));
OR2X2 OR2X2_5356 ( .A(alu__abc_42281_new_n860_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n1241_));
OR2X2 OR2X2_5357 ( .A(alu__abc_42281_new_n838_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1242_));
OR2X2 OR2X2_5358 ( .A(alu__abc_42281_new_n848_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n1245_));
OR2X2 OR2X2_5359 ( .A(alu__abc_42281_new_n907_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1246_));
OR2X2 OR2X2_536 ( .A(_abc_44694_new_n2190_), .B(_abc_44694_new_n2191_), .Y(_abc_44694_new_n2192_));
OR2X2 OR2X2_5360 ( .A(alu__abc_42281_new_n1248_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n1249_));
OR2X2 OR2X2_5361 ( .A(alu__abc_42281_new_n1249_), .B(alu__abc_42281_new_n1244_), .Y(alu__abc_42281_new_n1250_));
OR2X2 OR2X2_5362 ( .A(alu__abc_42281_new_n917_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n1251_));
OR2X2 OR2X2_5363 ( .A(alu__abc_42281_new_n885_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n1252_));
OR2X2 OR2X2_5364 ( .A(alu__abc_42281_new_n1253_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n1254_));
OR2X2 OR2X2_5365 ( .A(alu__abc_42281_new_n895_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n1255_));
OR2X2 OR2X2_5366 ( .A(alu__abc_42281_new_n962_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n1256_));
OR2X2 OR2X2_5367 ( .A(alu__abc_42281_new_n1257_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n1258_));
OR2X2 OR2X2_5368 ( .A(alu__abc_42281_new_n1259_), .B(alu__abc_42281_new_n271__bF_buf2), .Y(alu__abc_42281_new_n1260_));
OR2X2 OR2X2_5369 ( .A(alu__abc_42281_new_n931_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n1264_));
OR2X2 OR2X2_537 ( .A(_abc_44694_new_n1334__bF_buf2), .B(_abc_44694_new_n2192_), .Y(_abc_44694_new_n2193_));
OR2X2 OR2X2_5370 ( .A(alu__abc_42281_new_n1265_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n1266_));
OR2X2 OR2X2_5371 ( .A(alu__abc_42281_new_n1133_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n1267_));
OR2X2 OR2X2_5372 ( .A(alu__abc_42281_new_n1268_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1269_));
OR2X2 OR2X2_5373 ( .A(alu__abc_42281_new_n1275_), .B(alu__abc_42281_new_n1276_), .Y(alu__abc_42281_new_n1277_));
OR2X2 OR2X2_5374 ( .A(alu__abc_42281_new_n1277_), .B(alu__abc_42281_new_n1274_), .Y(alu__abc_42281_new_n1278_));
OR2X2 OR2X2_5375 ( .A(alu__abc_42281_new_n1278_), .B(alu__abc_42281_new_n1273_), .Y(alu__abc_42281_new_n1279_));
OR2X2 OR2X2_5376 ( .A(alu__abc_42281_new_n1272_), .B(alu__abc_42281_new_n1279_), .Y(alu__abc_42281_new_n1280_));
OR2X2 OR2X2_5377 ( .A(alu__abc_42281_new_n1263_), .B(alu__abc_42281_new_n1280_), .Y(alu__abc_42281_new_n1281_));
OR2X2 OR2X2_5378 ( .A(alu__abc_42281_new_n1262_), .B(alu__abc_42281_new_n1281_), .Y(alu__abc_42281_new_n1282_));
OR2X2 OR2X2_5379 ( .A(alu__abc_42281_new_n1282_), .B(alu__abc_42281_new_n1240_), .Y(alu__abc_42281_new_n1283_));
OR2X2 OR2X2_538 ( .A(_abc_44694_new_n2195_), .B(_abc_44694_new_n2168_), .Y(_abc_44694_new_n2196_));
OR2X2 OR2X2_5380 ( .A(alu__abc_42281_new_n1283_), .B(alu__abc_42281_new_n1236_), .Y(alu_p_o_4_));
OR2X2 OR2X2_5381 ( .A(alu__abc_42281_new_n749_), .B(alu__abc_42281_new_n770_), .Y(alu__abc_42281_new_n1287_));
OR2X2 OR2X2_5382 ( .A(alu__abc_42281_new_n1289_), .B(alu__abc_42281_new_n1285_), .Y(alu__abc_42281_new_n1290_));
OR2X2 OR2X2_5383 ( .A(alu__abc_42281_new_n1291_), .B(alu__abc_42281_new_n589_), .Y(alu__abc_42281_new_n1292_));
OR2X2 OR2X2_5384 ( .A(alu__abc_42281_new_n407_), .B(alu__abc_42281_new_n268_), .Y(alu__abc_42281_new_n1293_));
OR2X2 OR2X2_5385 ( .A(alu__abc_42281_new_n970_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n1296_));
OR2X2 OR2X2_5386 ( .A(alu__abc_42281_new_n1002_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n1299_));
OR2X2 OR2X2_5387 ( .A(alu__abc_42281_new_n980_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n1300_));
OR2X2 OR2X2_5388 ( .A(alu__abc_42281_new_n1298_), .B(alu__abc_42281_new_n1302_), .Y(alu__abc_42281_new_n1303_));
OR2X2 OR2X2_5389 ( .A(alu__abc_42281_new_n1303_), .B(alu__abc_42281_new_n271__bF_buf1), .Y(alu__abc_42281_new_n1304_));
OR2X2 OR2X2_539 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_22_), .Y(_abc_44694_new_n2197_));
OR2X2 OR2X2_5390 ( .A(alu__abc_42281_new_n1306_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n1307_));
OR2X2 OR2X2_5391 ( .A(alu__abc_42281_new_n1307_), .B(alu__abc_42281_new_n1305_), .Y(alu__abc_42281_new_n1308_));
OR2X2 OR2X2_5392 ( .A(alu__abc_42281_new_n1048_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n1309_));
OR2X2 OR2X2_5393 ( .A(alu__abc_42281_new_n992_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1310_));
OR2X2 OR2X2_5394 ( .A(alu__abc_42281_new_n1311_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n1312_));
OR2X2 OR2X2_5395 ( .A(alu__abc_42281_new_n1313_), .B(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n1314_));
OR2X2 OR2X2_5396 ( .A(alu__abc_42281_new_n1072_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1317_));
OR2X2 OR2X2_5397 ( .A(alu__abc_42281_new_n1318_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n1319_));
OR2X2 OR2X2_5398 ( .A(alu__abc_42281_new_n1210_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n1320_));
OR2X2 OR2X2_5399 ( .A(alu__abc_42281_new_n1321_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n1322_));
OR2X2 OR2X2_54 ( .A(_abc_44694_new_n793_), .B(_abc_44694_new_n779_), .Y(REGFILE_SIM_reg_bank_reg_rd_i_6_));
OR2X2 OR2X2_540 ( .A(_abc_44694_new_n2164_), .B(pc_q_23_), .Y(_abc_44694_new_n2200_));
OR2X2 OR2X2_5400 ( .A(alu__abc_42281_new_n1328_), .B(alu__abc_42281_new_n1327_), .Y(alu__abc_42281_new_n1329_));
OR2X2 OR2X2_5401 ( .A(alu__abc_42281_new_n1329_), .B(alu__abc_42281_new_n1330_), .Y(alu__abc_42281_new_n1331_));
OR2X2 OR2X2_5402 ( .A(alu__abc_42281_new_n1331_), .B(alu__abc_42281_new_n1326_), .Y(alu__abc_42281_new_n1332_));
OR2X2 OR2X2_5403 ( .A(alu__abc_42281_new_n1325_), .B(alu__abc_42281_new_n1332_), .Y(alu__abc_42281_new_n1333_));
OR2X2 OR2X2_5404 ( .A(alu__abc_42281_new_n1316_), .B(alu__abc_42281_new_n1333_), .Y(alu__abc_42281_new_n1334_));
OR2X2 OR2X2_5405 ( .A(alu__abc_42281_new_n1295_), .B(alu__abc_42281_new_n1334_), .Y(alu__abc_42281_new_n1335_));
OR2X2 OR2X2_5406 ( .A(alu__abc_42281_new_n1290_), .B(alu__abc_42281_new_n1335_), .Y(alu_p_o_5_));
OR2X2 OR2X2_5407 ( .A(alu__abc_42281_new_n409_), .B(alu__abc_42281_new_n257_), .Y(alu__abc_42281_new_n1337_));
OR2X2 OR2X2_5408 ( .A(alu__abc_42281_new_n771_), .B(alu__abc_42281_new_n742_), .Y(alu__abc_42281_new_n1342_));
OR2X2 OR2X2_5409 ( .A(alu__abc_42281_new_n1085_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n1346_));
OR2X2 OR2X2_541 ( .A(_abc_44694_new_n2204_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n2205_));
OR2X2 OR2X2_5410 ( .A(alu__abc_42281_new_n1099_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1349_));
OR2X2 OR2X2_5411 ( .A(alu__abc_42281_new_n1089_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n1350_));
OR2X2 OR2X2_5412 ( .A(alu__abc_42281_new_n1348_), .B(alu__abc_42281_new_n1352_), .Y(alu__abc_42281_new_n1353_));
OR2X2 OR2X2_5413 ( .A(alu__abc_42281_new_n1353_), .B(alu__abc_42281_new_n271__bF_buf0), .Y(alu__abc_42281_new_n1354_));
OR2X2 OR2X2_5414 ( .A(alu__abc_42281_new_n1111_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n1355_));
OR2X2 OR2X2_5415 ( .A(alu__abc_42281_new_n1117_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n1356_));
OR2X2 OR2X2_5416 ( .A(alu__abc_42281_new_n1121_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n1359_));
OR2X2 OR2X2_5417 ( .A(alu__abc_42281_new_n1095_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n1360_));
OR2X2 OR2X2_5418 ( .A(alu__abc_42281_new_n1362_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n1363_));
OR2X2 OR2X2_5419 ( .A(alu__abc_42281_new_n1363_), .B(alu__abc_42281_new_n1358_), .Y(alu__abc_42281_new_n1364_));
OR2X2 OR2X2_542 ( .A(_abc_44694_new_n2203_), .B(_abc_44694_new_n1399__bF_buf2), .Y(_abc_44694_new_n2206_));
OR2X2 OR2X2_5420 ( .A(alu__abc_42281_new_n1137_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n1367_));
OR2X2 OR2X2_5421 ( .A(alu__abc_42281_new_n1368_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n1369_));
OR2X2 OR2X2_5422 ( .A(alu__abc_42281_new_n1265_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n1370_));
OR2X2 OR2X2_5423 ( .A(alu__abc_42281_new_n1371_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n1372_));
OR2X2 OR2X2_5424 ( .A(alu__abc_42281_new_n1378_), .B(alu__abc_42281_new_n1379_), .Y(alu__abc_42281_new_n1380_));
OR2X2 OR2X2_5425 ( .A(alu__abc_42281_new_n1380_), .B(alu__abc_42281_new_n1377_), .Y(alu__abc_42281_new_n1381_));
OR2X2 OR2X2_5426 ( .A(alu__abc_42281_new_n1381_), .B(alu__abc_42281_new_n1376_), .Y(alu__abc_42281_new_n1382_));
OR2X2 OR2X2_5427 ( .A(alu__abc_42281_new_n1375_), .B(alu__abc_42281_new_n1382_), .Y(alu__abc_42281_new_n1383_));
OR2X2 OR2X2_5428 ( .A(alu__abc_42281_new_n1366_), .B(alu__abc_42281_new_n1383_), .Y(alu__abc_42281_new_n1384_));
OR2X2 OR2X2_5429 ( .A(alu__abc_42281_new_n1384_), .B(alu__abc_42281_new_n1345_), .Y(alu__abc_42281_new_n1385_));
OR2X2 OR2X2_543 ( .A(opcode_q_21_), .B(pc_q_23_), .Y(_abc_44694_new_n2210_));
OR2X2 OR2X2_5430 ( .A(alu__abc_42281_new_n1344_), .B(alu__abc_42281_new_n1385_), .Y(alu__abc_42281_new_n1386_));
OR2X2 OR2X2_5431 ( .A(alu__abc_42281_new_n1386_), .B(alu__abc_42281_new_n1340_), .Y(alu_p_o_6_));
OR2X2 OR2X2_5432 ( .A(alu__abc_42281_new_n411_), .B(alu__abc_42281_new_n262_), .Y(alu__abc_42281_new_n1388_));
OR2X2 OR2X2_5433 ( .A(alu__abc_42281_new_n1389_), .B(alu__abc_42281_new_n587_), .Y(alu__abc_42281_new_n1390_));
OR2X2 OR2X2_5434 ( .A(alu__abc_42281_new_n740_), .B(alu__abc_42281_new_n772_), .Y(alu__abc_42281_new_n1394_));
OR2X2 OR2X2_5435 ( .A(alu__abc_42281_new_n1159_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n1398_));
OR2X2 OR2X2_5436 ( .A(alu__abc_42281_new_n1173_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n1401_));
OR2X2 OR2X2_5437 ( .A(alu__abc_42281_new_n1163_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n1402_));
OR2X2 OR2X2_5438 ( .A(alu__abc_42281_new_n1400_), .B(alu__abc_42281_new_n1404_), .Y(alu__abc_42281_new_n1405_));
OR2X2 OR2X2_5439 ( .A(alu__abc_42281_new_n1405_), .B(alu__abc_42281_new_n271__bF_buf4), .Y(alu__abc_42281_new_n1406_));
OR2X2 OR2X2_544 ( .A(_abc_44694_new_n2209_), .B(_abc_44694_new_n2213_), .Y(_abc_44694_new_n2214_));
OR2X2 OR2X2_5440 ( .A(alu__abc_42281_new_n1195_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n1407_));
OR2X2 OR2X2_5441 ( .A(alu__abc_42281_new_n1169_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1408_));
OR2X2 OR2X2_5442 ( .A(alu__abc_42281_new_n1185_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1411_));
OR2X2 OR2X2_5443 ( .A(alu__abc_42281_new_n1191_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1412_));
OR2X2 OR2X2_5444 ( .A(alu__abc_42281_new_n1414_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n1415_));
OR2X2 OR2X2_5445 ( .A(alu__abc_42281_new_n1415_), .B(alu__abc_42281_new_n1410_), .Y(alu__abc_42281_new_n1416_));
OR2X2 OR2X2_5446 ( .A(alu__abc_42281_new_n1420_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n1421_));
OR2X2 OR2X2_5447 ( .A(alu__abc_42281_new_n1318_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n1422_));
OR2X2 OR2X2_5448 ( .A(alu__abc_42281_new_n1419_), .B(alu__abc_42281_new_n1424_), .Y(alu__abc_42281_new_n1425_));
OR2X2 OR2X2_5449 ( .A(alu__abc_42281_new_n1430_), .B(alu__abc_42281_new_n1431_), .Y(alu__abc_42281_new_n1432_));
OR2X2 OR2X2_545 ( .A(_abc_44694_new_n2208_), .B(_abc_44694_new_n2215_), .Y(_abc_44694_new_n2216_));
OR2X2 OR2X2_5450 ( .A(alu__abc_42281_new_n1432_), .B(alu__abc_42281_new_n1429_), .Y(alu__abc_42281_new_n1433_));
OR2X2 OR2X2_5451 ( .A(alu__abc_42281_new_n1433_), .B(alu__abc_42281_new_n1428_), .Y(alu__abc_42281_new_n1434_));
OR2X2 OR2X2_5452 ( .A(alu__abc_42281_new_n1427_), .B(alu__abc_42281_new_n1434_), .Y(alu__abc_42281_new_n1435_));
OR2X2 OR2X2_5453 ( .A(alu__abc_42281_new_n1418_), .B(alu__abc_42281_new_n1435_), .Y(alu__abc_42281_new_n1436_));
OR2X2 OR2X2_5454 ( .A(alu__abc_42281_new_n1397_), .B(alu__abc_42281_new_n1436_), .Y(alu__abc_42281_new_n1437_));
OR2X2 OR2X2_5455 ( .A(alu__abc_42281_new_n1396_), .B(alu__abc_42281_new_n1437_), .Y(alu__abc_42281_new_n1438_));
OR2X2 OR2X2_5456 ( .A(alu__abc_42281_new_n1392_), .B(alu__abc_42281_new_n1438_), .Y(alu_p_o_7_));
OR2X2 OR2X2_5457 ( .A(alu__abc_42281_new_n413_), .B(alu__abc_42281_new_n364_), .Y(alu__abc_42281_new_n1442_));
OR2X2 OR2X2_5458 ( .A(alu__abc_42281_new_n773_), .B(alu__abc_42281_new_n731_), .Y(alu__abc_42281_new_n1446_));
OR2X2 OR2X2_5459 ( .A(alu__abc_42281_new_n897_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n1450_));
OR2X2 OR2X2_546 ( .A(_abc_44694_new_n2218_), .B(_abc_44694_new_n2207_), .Y(_abc_44694_new_n2219_));
OR2X2 OR2X2_5460 ( .A(alu__abc_42281_new_n962_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1451_));
OR2X2 OR2X2_5461 ( .A(alu__abc_42281_new_n1452_), .B(alu__abc_42281_new_n271__bF_buf3), .Y(alu__abc_42281_new_n1453_));
OR2X2 OR2X2_5462 ( .A(alu__abc_42281_new_n850_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n1454_));
OR2X2 OR2X2_5463 ( .A(alu__abc_42281_new_n919_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n1455_));
OR2X2 OR2X2_5464 ( .A(alu__abc_42281_new_n1456_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n1457_));
OR2X2 OR2X2_5465 ( .A(alu__abc_42281_new_n932_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n1460_));
OR2X2 OR2X2_5466 ( .A(alu__abc_42281_new_n1268_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n1461_));
OR2X2 OR2X2_5467 ( .A(alu__abc_42281_new_n1462_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n1463_));
OR2X2 OR2X2_5468 ( .A(alu__abc_42281_new_n1368_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n1464_));
OR2X2 OR2X2_5469 ( .A(alu__abc_42281_new_n1465_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n1466_));
OR2X2 OR2X2_547 ( .A(_abc_44694_new_n1400__bF_buf3), .B(_abc_44694_new_n2221_), .Y(_abc_44694_new_n2222_));
OR2X2 OR2X2_5470 ( .A(alu__abc_42281_new_n1467_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n1468_));
OR2X2 OR2X2_5471 ( .A(alu__abc_42281_new_n1472_), .B(alu__abc_42281_new_n1473_), .Y(alu__abc_42281_new_n1474_));
OR2X2 OR2X2_5472 ( .A(alu__abc_42281_new_n1474_), .B(alu__abc_42281_new_n1475_), .Y(alu__abc_42281_new_n1476_));
OR2X2 OR2X2_5473 ( .A(alu__abc_42281_new_n1476_), .B(alu__abc_42281_new_n1471_), .Y(alu__abc_42281_new_n1477_));
OR2X2 OR2X2_5474 ( .A(alu__abc_42281_new_n1470_), .B(alu__abc_42281_new_n1477_), .Y(alu__abc_42281_new_n1478_));
OR2X2 OR2X2_5475 ( .A(alu__abc_42281_new_n1459_), .B(alu__abc_42281_new_n1478_), .Y(alu__abc_42281_new_n1479_));
OR2X2 OR2X2_5476 ( .A(alu__abc_42281_new_n1479_), .B(alu__abc_42281_new_n1449_), .Y(alu__abc_42281_new_n1480_));
OR2X2 OR2X2_5477 ( .A(alu__abc_42281_new_n1448_), .B(alu__abc_42281_new_n1480_), .Y(alu__abc_42281_new_n1481_));
OR2X2 OR2X2_5478 ( .A(alu__abc_42281_new_n1444_), .B(alu__abc_42281_new_n1481_), .Y(alu_p_o_8_));
OR2X2 OR2X2_5479 ( .A(alu__abc_42281_new_n1484_), .B(alu__abc_42281_new_n372_), .Y(alu__abc_42281_new_n1485_));
OR2X2 OR2X2_548 ( .A(_abc_44694_new_n2220_), .B(_abc_44694_new_n2222_), .Y(_abc_44694_new_n2223_));
OR2X2 OR2X2_5480 ( .A(alu__abc_42281_new_n1483_), .B(alu__abc_42281_new_n371_), .Y(alu__abc_42281_new_n1486_));
OR2X2 OR2X2_5481 ( .A(alu__abc_42281_new_n774_), .B(alu__abc_42281_new_n728_), .Y(alu__abc_42281_new_n1490_));
OR2X2 OR2X2_5482 ( .A(alu__abc_42281_new_n982_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n1494_));
OR2X2 OR2X2_5483 ( .A(alu__abc_42281_new_n1495_), .B(alu__abc_42281_new_n271__bF_buf2), .Y(alu__abc_42281_new_n1496_));
OR2X2 OR2X2_5484 ( .A(alu__abc_42281_new_n1498_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n1499_));
OR2X2 OR2X2_5485 ( .A(alu__abc_42281_new_n1499_), .B(alu__abc_42281_new_n1497_), .Y(alu__abc_42281_new_n1500_));
OR2X2 OR2X2_5486 ( .A(alu__abc_42281_new_n1504_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n1505_));
OR2X2 OR2X2_5487 ( .A(alu__abc_42281_new_n1420_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n1506_));
OR2X2 OR2X2_5488 ( .A(alu__abc_42281_new_n1507_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n1508_));
OR2X2 OR2X2_5489 ( .A(alu__abc_42281_new_n1321_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n1509_));
OR2X2 OR2X2_549 ( .A(_abc_44694_new_n2224_), .B(_abc_44694_new_n1278__bF_buf3), .Y(_abc_44694_new_n2225_));
OR2X2 OR2X2_5490 ( .A(alu__abc_42281_new_n1511_), .B(alu__abc_42281_new_n1503_), .Y(alu__abc_42281_new_n1512_));
OR2X2 OR2X2_5491 ( .A(alu__abc_42281_new_n1516_), .B(alu__abc_42281_new_n1517_), .Y(alu__abc_42281_new_n1518_));
OR2X2 OR2X2_5492 ( .A(alu__abc_42281_new_n1518_), .B(alu__abc_42281_new_n1515_), .Y(alu__abc_42281_new_n1519_));
OR2X2 OR2X2_5493 ( .A(alu__abc_42281_new_n1519_), .B(alu__abc_42281_new_n1514_), .Y(alu__abc_42281_new_n1520_));
OR2X2 OR2X2_5494 ( .A(alu__abc_42281_new_n1513_), .B(alu__abc_42281_new_n1520_), .Y(alu__abc_42281_new_n1521_));
OR2X2 OR2X2_5495 ( .A(alu__abc_42281_new_n1502_), .B(alu__abc_42281_new_n1521_), .Y(alu__abc_42281_new_n1522_));
OR2X2 OR2X2_5496 ( .A(alu__abc_42281_new_n1493_), .B(alu__abc_42281_new_n1522_), .Y(alu__abc_42281_new_n1523_));
OR2X2 OR2X2_5497 ( .A(alu__abc_42281_new_n1492_), .B(alu__abc_42281_new_n1523_), .Y(alu__abc_42281_new_n1524_));
OR2X2 OR2X2_5498 ( .A(alu__abc_42281_new_n1488_), .B(alu__abc_42281_new_n1524_), .Y(alu_p_o_9_));
OR2X2 OR2X2_5499 ( .A(alu__abc_42281_new_n1526_), .B(alu__abc_42281_new_n422_), .Y(alu__abc_42281_new_n1527_));
OR2X2 OR2X2_55 ( .A(_abc_44694_new_n795_), .B(_abc_44694_new_n796_), .Y(_abc_44694_new_n797_));
OR2X2 OR2X2_550 ( .A(_abc_44694_new_n2226_), .B(_abc_44694_new_n2227_), .Y(_abc_44694_new_n2228_));
OR2X2 OR2X2_5500 ( .A(alu__abc_42281_new_n1527_), .B(alu__abc_42281_new_n347_), .Y(alu__abc_42281_new_n1530_));
OR2X2 OR2X2_5501 ( .A(alu__abc_42281_new_n775_), .B(alu__abc_42281_new_n790_), .Y(alu__abc_42281_new_n1533_));
OR2X2 OR2X2_5502 ( .A(alu__abc_42281_new_n1091_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n1540_));
OR2X2 OR2X2_5503 ( .A(alu__abc_42281_new_n1541_), .B(alu__abc_42281_new_n271__bF_buf1), .Y(alu__abc_42281_new_n1542_));
OR2X2 OR2X2_5504 ( .A(alu__abc_42281_new_n1544_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n1545_));
OR2X2 OR2X2_5505 ( .A(alu__abc_42281_new_n1545_), .B(alu__abc_42281_new_n1543_), .Y(alu__abc_42281_new_n1546_));
OR2X2 OR2X2_5506 ( .A(alu__abc_42281_new_n1550_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n1551_));
OR2X2 OR2X2_5507 ( .A(alu__abc_42281_new_n1462_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n1552_));
OR2X2 OR2X2_5508 ( .A(alu__abc_42281_new_n1553_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n1554_));
OR2X2 OR2X2_5509 ( .A(alu__abc_42281_new_n1371_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n1555_));
OR2X2 OR2X2_551 ( .A(_abc_44694_new_n1334__bF_buf1), .B(_abc_44694_new_n2228_), .Y(_abc_44694_new_n2229_));
OR2X2 OR2X2_5510 ( .A(alu__abc_42281_new_n1557_), .B(alu__abc_42281_new_n1549_), .Y(alu__abc_42281_new_n1558_));
OR2X2 OR2X2_5511 ( .A(alu__abc_42281_new_n1561_), .B(alu__abc_42281_new_n1562_), .Y(alu__abc_42281_new_n1563_));
OR2X2 OR2X2_5512 ( .A(alu__abc_42281_new_n1563_), .B(alu__abc_42281_new_n1560_), .Y(alu__abc_42281_new_n1564_));
OR2X2 OR2X2_5513 ( .A(alu__abc_42281_new_n1559_), .B(alu__abc_42281_new_n1564_), .Y(alu__abc_42281_new_n1565_));
OR2X2 OR2X2_5514 ( .A(alu__abc_42281_new_n1548_), .B(alu__abc_42281_new_n1565_), .Y(alu__abc_42281_new_n1566_));
OR2X2 OR2X2_5515 ( .A(alu__abc_42281_new_n1539_), .B(alu__abc_42281_new_n1566_), .Y(alu__abc_42281_new_n1567_));
OR2X2 OR2X2_5516 ( .A(alu__abc_42281_new_n1567_), .B(alu__abc_42281_new_n1538_), .Y(alu__abc_42281_new_n1568_));
OR2X2 OR2X2_5517 ( .A(alu__abc_42281_new_n1537_), .B(alu__abc_42281_new_n1568_), .Y(alu__abc_42281_new_n1569_));
OR2X2 OR2X2_5518 ( .A(alu__abc_42281_new_n1532_), .B(alu__abc_42281_new_n1569_), .Y(alu_p_o_10_));
OR2X2 OR2X2_5519 ( .A(alu__abc_42281_new_n1528_), .B(alu__abc_42281_new_n425_), .Y(alu__abc_42281_new_n1571_));
OR2X2 OR2X2_552 ( .A(_abc_44694_new_n2231_), .B(_abc_44694_new_n2205_), .Y(_abc_44694_new_n2232_));
OR2X2 OR2X2_5520 ( .A(alu__abc_42281_new_n1571_), .B(alu__abc_42281_new_n355_), .Y(alu__abc_42281_new_n1572_));
OR2X2 OR2X2_5521 ( .A(alu__abc_42281_new_n1573_), .B(alu__abc_42281_new_n354_), .Y(alu__abc_42281_new_n1574_));
OR2X2 OR2X2_5522 ( .A(alu__abc_42281_new_n1534_), .B(alu__abc_42281_new_n800_), .Y(alu__abc_42281_new_n1579_));
OR2X2 OR2X2_5523 ( .A(alu__abc_42281_new_n1165_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n1582_));
OR2X2 OR2X2_5524 ( .A(alu__abc_42281_new_n1583_), .B(alu__abc_42281_new_n271__bF_buf0), .Y(alu__abc_42281_new_n1584_));
OR2X2 OR2X2_5525 ( .A(alu__abc_42281_new_n1197_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n1585_));
OR2X2 OR2X2_5526 ( .A(alu__abc_42281_new_n1175_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1586_));
OR2X2 OR2X2_5527 ( .A(alu__abc_42281_new_n1587_), .B(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n1588_));
OR2X2 OR2X2_5528 ( .A(alu__abc_42281_new_n1593_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n1594_));
OR2X2 OR2X2_5529 ( .A(alu__abc_42281_new_n1504_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n1595_));
OR2X2 OR2X2_553 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_23_), .Y(_abc_44694_new_n2233_));
OR2X2 OR2X2_5530 ( .A(alu__abc_42281_new_n1596_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n1597_));
OR2X2 OR2X2_5531 ( .A(alu__abc_42281_new_n1423_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n1598_));
OR2X2 OR2X2_5532 ( .A(alu__abc_42281_new_n1600_), .B(alu__abc_42281_new_n1592_), .Y(alu__abc_42281_new_n1601_));
OR2X2 OR2X2_5533 ( .A(alu__abc_42281_new_n1604_), .B(alu__abc_42281_new_n1605_), .Y(alu__abc_42281_new_n1606_));
OR2X2 OR2X2_5534 ( .A(alu__abc_42281_new_n1606_), .B(alu__abc_42281_new_n1607_), .Y(alu__abc_42281_new_n1608_));
OR2X2 OR2X2_5535 ( .A(alu__abc_42281_new_n1608_), .B(alu__abc_42281_new_n1603_), .Y(alu__abc_42281_new_n1609_));
OR2X2 OR2X2_5536 ( .A(alu__abc_42281_new_n1602_), .B(alu__abc_42281_new_n1609_), .Y(alu__abc_42281_new_n1610_));
OR2X2 OR2X2_5537 ( .A(alu__abc_42281_new_n1591_), .B(alu__abc_42281_new_n1610_), .Y(alu__abc_42281_new_n1611_));
OR2X2 OR2X2_5538 ( .A(alu__abc_42281_new_n1611_), .B(alu__abc_42281_new_n1590_), .Y(alu__abc_42281_new_n1612_));
OR2X2 OR2X2_5539 ( .A(alu__abc_42281_new_n1581_), .B(alu__abc_42281_new_n1612_), .Y(alu__abc_42281_new_n1613_));
OR2X2 OR2X2_554 ( .A(_abc_44694_new_n2201_), .B(pc_q_24_), .Y(_abc_44694_new_n2236_));
OR2X2 OR2X2_5540 ( .A(alu__abc_42281_new_n1576_), .B(alu__abc_42281_new_n1613_), .Y(alu_p_o_11_));
OR2X2 OR2X2_5541 ( .A(alu__abc_42281_new_n1615_), .B(alu__abc_42281_new_n428_), .Y(alu__abc_42281_new_n1616_));
OR2X2 OR2X2_5542 ( .A(alu__abc_42281_new_n1616_), .B(alu__abc_42281_new_n312_), .Y(alu__abc_42281_new_n1617_));
OR2X2 OR2X2_5543 ( .A(alu__abc_42281_new_n1577_), .B(alu__abc_42281_new_n792_), .Y(alu__abc_42281_new_n1622_));
OR2X2 OR2X2_5544 ( .A(alu__abc_42281_new_n1628_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n1629_));
OR2X2 OR2X2_5545 ( .A(alu__abc_42281_new_n1629_), .B(alu__abc_42281_new_n1627_), .Y(alu__abc_42281_new_n1630_));
OR2X2 OR2X2_5546 ( .A(alu__abc_42281_new_n1257_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n1631_));
OR2X2 OR2X2_5547 ( .A(alu__abc_42281_new_n1632_), .B(alu__abc_42281_new_n271__bF_buf4), .Y(alu__abc_42281_new_n1633_));
OR2X2 OR2X2_5548 ( .A(alu__abc_42281_new_n1637_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n1638_));
OR2X2 OR2X2_5549 ( .A(alu__abc_42281_new_n1550_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n1639_));
OR2X2 OR2X2_555 ( .A(_abc_44694_new_n2240_), .B(_abc_44694_new_n1210__bF_buf1), .Y(_abc_44694_new_n2241_));
OR2X2 OR2X2_5550 ( .A(alu__abc_42281_new_n1640_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n1641_));
OR2X2 OR2X2_5551 ( .A(alu__abc_42281_new_n1465_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1642_));
OR2X2 OR2X2_5552 ( .A(alu__abc_42281_new_n1643_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n1644_));
OR2X2 OR2X2_5553 ( .A(alu__abc_42281_new_n1270_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n1645_));
OR2X2 OR2X2_5554 ( .A(alu__abc_42281_new_n1650_), .B(alu__abc_42281_new_n1651_), .Y(alu__abc_42281_new_n1652_));
OR2X2 OR2X2_5555 ( .A(alu__abc_42281_new_n1652_), .B(alu__abc_42281_new_n1649_), .Y(alu__abc_42281_new_n1653_));
OR2X2 OR2X2_5556 ( .A(alu__abc_42281_new_n1653_), .B(alu__abc_42281_new_n1648_), .Y(alu__abc_42281_new_n1654_));
OR2X2 OR2X2_5557 ( .A(alu__abc_42281_new_n1647_), .B(alu__abc_42281_new_n1654_), .Y(alu__abc_42281_new_n1655_));
OR2X2 OR2X2_5558 ( .A(alu__abc_42281_new_n1636_), .B(alu__abc_42281_new_n1655_), .Y(alu__abc_42281_new_n1656_));
OR2X2 OR2X2_5559 ( .A(alu__abc_42281_new_n1656_), .B(alu__abc_42281_new_n1635_), .Y(alu__abc_42281_new_n1657_));
OR2X2 OR2X2_556 ( .A(_abc_44694_new_n2249_), .B(_abc_44694_new_n2211_), .Y(_abc_44694_new_n2250_));
OR2X2 OR2X2_5560 ( .A(alu__abc_42281_new_n1626_), .B(alu__abc_42281_new_n1657_), .Y(alu__abc_42281_new_n1658_));
OR2X2 OR2X2_5561 ( .A(alu__abc_42281_new_n1658_), .B(alu__abc_42281_new_n1621_), .Y(alu_p_o_12_));
OR2X2 OR2X2_5562 ( .A(alu__abc_42281_new_n1661_), .B(alu__abc_42281_new_n320_), .Y(alu__abc_42281_new_n1662_));
OR2X2 OR2X2_5563 ( .A(alu__abc_42281_new_n1660_), .B(alu__abc_42281_new_n319_), .Y(alu__abc_42281_new_n1663_));
OR2X2 OR2X2_5564 ( .A(alu__abc_42281_new_n1623_), .B(alu__abc_42281_new_n782_), .Y(alu__abc_42281_new_n1668_));
OR2X2 OR2X2_5565 ( .A(alu__abc_42281_new_n1297_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n1671_));
OR2X2 OR2X2_5566 ( .A(alu__abc_42281_new_n1672_), .B(alu__abc_42281_new_n271__bF_buf3), .Y(alu__abc_42281_new_n1673_));
OR2X2 OR2X2_5567 ( .A(alu__abc_42281_new_n1675_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n1676_));
OR2X2 OR2X2_5568 ( .A(alu__abc_42281_new_n1676_), .B(alu__abc_42281_new_n1674_), .Y(alu__abc_42281_new_n1677_));
OR2X2 OR2X2_5569 ( .A(alu__abc_42281_new_n1681_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n1682_));
OR2X2 OR2X2_557 ( .A(_abc_44694_new_n2248_), .B(_abc_44694_new_n2250_), .Y(_abc_44694_new_n2251_));
OR2X2 OR2X2_5570 ( .A(alu__abc_42281_new_n1593_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n1683_));
OR2X2 OR2X2_5571 ( .A(alu__abc_42281_new_n1684_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1685_));
OR2X2 OR2X2_5572 ( .A(alu__abc_42281_new_n1507_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1686_));
OR2X2 OR2X2_5573 ( .A(alu__abc_42281_new_n1687_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n1688_));
OR2X2 OR2X2_5574 ( .A(alu__abc_42281_new_n1323_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n1689_));
OR2X2 OR2X2_5575 ( .A(alu__abc_42281_new_n1693_), .B(alu__abc_42281_new_n1694_), .Y(alu__abc_42281_new_n1695_));
OR2X2 OR2X2_5576 ( .A(alu__abc_42281_new_n1695_), .B(alu__abc_42281_new_n1696_), .Y(alu__abc_42281_new_n1697_));
OR2X2 OR2X2_5577 ( .A(alu__abc_42281_new_n1697_), .B(alu__abc_42281_new_n1692_), .Y(alu__abc_42281_new_n1698_));
OR2X2 OR2X2_5578 ( .A(alu__abc_42281_new_n1691_), .B(alu__abc_42281_new_n1698_), .Y(alu__abc_42281_new_n1699_));
OR2X2 OR2X2_5579 ( .A(alu__abc_42281_new_n1680_), .B(alu__abc_42281_new_n1699_), .Y(alu__abc_42281_new_n1700_));
OR2X2 OR2X2_558 ( .A(_abc_44694_new_n2251_), .B(_abc_44694_new_n2247_), .Y(_abc_44694_new_n2252_));
OR2X2 OR2X2_5580 ( .A(alu__abc_42281_new_n1700_), .B(alu__abc_42281_new_n1679_), .Y(alu__abc_42281_new_n1701_));
OR2X2 OR2X2_5581 ( .A(alu__abc_42281_new_n1670_), .B(alu__abc_42281_new_n1701_), .Y(alu__abc_42281_new_n1702_));
OR2X2 OR2X2_5582 ( .A(alu__abc_42281_new_n1665_), .B(alu__abc_42281_new_n1702_), .Y(alu_p_o_13_));
OR2X2 OR2X2_5583 ( .A(alu__abc_42281_new_n1704_), .B(alu__abc_42281_new_n437_), .Y(alu__abc_42281_new_n1705_));
OR2X2 OR2X2_5584 ( .A(alu__abc_42281_new_n1705_), .B(alu__abc_42281_new_n329_), .Y(alu__abc_42281_new_n1706_));
OR2X2 OR2X2_5585 ( .A(alu__abc_42281_new_n1666_), .B(alu__abc_42281_new_n802_), .Y(alu__abc_42281_new_n1711_));
OR2X2 OR2X2_5586 ( .A(alu__abc_42281_new_n1347_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n1717_));
OR2X2 OR2X2_5587 ( .A(alu__abc_42281_new_n1718_), .B(alu__abc_42281_new_n271__bF_buf2), .Y(alu__abc_42281_new_n1719_));
OR2X2 OR2X2_5588 ( .A(alu__abc_42281_new_n1721_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n1722_));
OR2X2 OR2X2_5589 ( .A(alu__abc_42281_new_n1722_), .B(alu__abc_42281_new_n1720_), .Y(alu__abc_42281_new_n1723_));
OR2X2 OR2X2_559 ( .A(_abc_44694_new_n2245_), .B(_abc_44694_new_n2252_), .Y(_abc_44694_new_n2253_));
OR2X2 OR2X2_5590 ( .A(alu__abc_42281_new_n1726_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n1727_));
OR2X2 OR2X2_5591 ( .A(alu__abc_42281_new_n1637_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n1728_));
OR2X2 OR2X2_5592 ( .A(alu__abc_42281_new_n1729_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n1730_));
OR2X2 OR2X2_5593 ( .A(alu__abc_42281_new_n1553_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n1731_));
OR2X2 OR2X2_5594 ( .A(alu__abc_42281_new_n1732_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n1733_));
OR2X2 OR2X2_5595 ( .A(alu__abc_42281_new_n1373_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n1734_));
OR2X2 OR2X2_5596 ( .A(alu__abc_42281_new_n1739_), .B(alu__abc_42281_new_n1738_), .Y(alu__abc_42281_new_n1740_));
OR2X2 OR2X2_5597 ( .A(alu__abc_42281_new_n1740_), .B(alu__abc_42281_new_n1741_), .Y(alu__abc_42281_new_n1742_));
OR2X2 OR2X2_5598 ( .A(alu__abc_42281_new_n1742_), .B(alu__abc_42281_new_n1737_), .Y(alu__abc_42281_new_n1743_));
OR2X2 OR2X2_5599 ( .A(alu__abc_42281_new_n1736_), .B(alu__abc_42281_new_n1743_), .Y(alu__abc_42281_new_n1744_));
OR2X2 OR2X2_56 ( .A(_abc_44694_new_n798_), .B(_abc_44694_new_n799_), .Y(_abc_44694_new_n800_));
OR2X2 OR2X2_560 ( .A(opcode_q_22_), .B(pc_q_24_), .Y(_abc_44694_new_n2254_));
OR2X2 OR2X2_5600 ( .A(alu__abc_42281_new_n1725_), .B(alu__abc_42281_new_n1744_), .Y(alu__abc_42281_new_n1745_));
OR2X2 OR2X2_5601 ( .A(alu__abc_42281_new_n1716_), .B(alu__abc_42281_new_n1745_), .Y(alu__abc_42281_new_n1746_));
OR2X2 OR2X2_5602 ( .A(alu__abc_42281_new_n1715_), .B(alu__abc_42281_new_n1746_), .Y(alu__abc_42281_new_n1747_));
OR2X2 OR2X2_5603 ( .A(alu__abc_42281_new_n1747_), .B(alu__abc_42281_new_n1710_), .Y(alu_p_o_14_));
OR2X2 OR2X2_5604 ( .A(alu__abc_42281_new_n1707_), .B(alu__abc_42281_new_n440_), .Y(alu__abc_42281_new_n1749_));
OR2X2 OR2X2_5605 ( .A(alu__abc_42281_new_n1750_), .B(alu__abc_42281_new_n336_), .Y(alu__abc_42281_new_n1751_));
OR2X2 OR2X2_5606 ( .A(alu__abc_42281_new_n1749_), .B(alu__abc_42281_new_n337_), .Y(alu__abc_42281_new_n1752_));
OR2X2 OR2X2_5607 ( .A(alu__abc_42281_new_n1712_), .B(alu__abc_42281_new_n721_), .Y(alu__abc_42281_new_n1755_));
OR2X2 OR2X2_5608 ( .A(alu__abc_42281_new_n1758_), .B(alu__abc_42281_new_n1756_), .Y(alu__abc_42281_new_n1759_));
OR2X2 OR2X2_5609 ( .A(alu__abc_42281_new_n1399_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n1761_));
OR2X2 OR2X2_561 ( .A(_abc_44694_new_n2253_), .B(_abc_44694_new_n2257_), .Y(_abc_44694_new_n2258_));
OR2X2 OR2X2_5610 ( .A(alu__abc_42281_new_n1762_), .B(alu__abc_42281_new_n271__bF_buf1), .Y(alu__abc_42281_new_n1763_));
OR2X2 OR2X2_5611 ( .A(alu__abc_42281_new_n1765_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n1766_));
OR2X2 OR2X2_5612 ( .A(alu__abc_42281_new_n1766_), .B(alu__abc_42281_new_n1764_), .Y(alu__abc_42281_new_n1767_));
OR2X2 OR2X2_5613 ( .A(alu__abc_42281_new_n1771_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n1772_));
OR2X2 OR2X2_5614 ( .A(alu__abc_42281_new_n1681_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n1773_));
OR2X2 OR2X2_5615 ( .A(alu__abc_42281_new_n1774_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n1775_));
OR2X2 OR2X2_5616 ( .A(alu__abc_42281_new_n1596_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n1776_));
OR2X2 OR2X2_5617 ( .A(alu__abc_42281_new_n1770_), .B(alu__abc_42281_new_n1778_), .Y(alu__abc_42281_new_n1779_));
OR2X2 OR2X2_5618 ( .A(alu__abc_42281_new_n1782_), .B(alu__abc_42281_new_n1781_), .Y(alu__abc_42281_new_n1783_));
OR2X2 OR2X2_5619 ( .A(alu__abc_42281_new_n1784_), .B(alu__abc_42281_new_n1785_), .Y(alu__abc_42281_new_n1786_));
OR2X2 OR2X2_562 ( .A(_abc_44694_new_n2262_), .B(_abc_44694_new_n2263_), .Y(_abc_44694_new_n2264_));
OR2X2 OR2X2_5620 ( .A(alu__abc_42281_new_n1786_), .B(alu__abc_42281_new_n1783_), .Y(alu__abc_42281_new_n1787_));
OR2X2 OR2X2_5621 ( .A(alu__abc_42281_new_n1780_), .B(alu__abc_42281_new_n1787_), .Y(alu__abc_42281_new_n1788_));
OR2X2 OR2X2_5622 ( .A(alu__abc_42281_new_n1769_), .B(alu__abc_42281_new_n1788_), .Y(alu__abc_42281_new_n1789_));
OR2X2 OR2X2_5623 ( .A(alu__abc_42281_new_n1760_), .B(alu__abc_42281_new_n1789_), .Y(alu__abc_42281_new_n1790_));
OR2X2 OR2X2_5624 ( .A(alu__abc_42281_new_n1754_), .B(alu__abc_42281_new_n1790_), .Y(alu_p_o_15_));
OR2X2 OR2X2_5625 ( .A(alu__abc_42281_new_n806_), .B(alu__abc_42281_new_n692_), .Y(alu__abc_42281_new_n1792_));
OR2X2 OR2X2_5626 ( .A(alu__abc_42281_new_n445_), .B(alu__abc_42281_new_n169_), .Y(alu__abc_42281_new_n1796_));
OR2X2 OR2X2_5627 ( .A(alu__abc_42281_new_n961_), .B(alu__abc_42281_new_n271__bF_buf0), .Y(alu__abc_42281_new_n1802_));
OR2X2 OR2X2_5628 ( .A(alu__abc_42281_new_n921_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n1804_));
OR2X2 OR2X2_5629 ( .A(alu__abc_42281_new_n1640_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n1806_));
OR2X2 OR2X2_563 ( .A(_abc_44694_new_n2265_), .B(_abc_44694_new_n2266_), .Y(_abc_44694_new_n2267_));
OR2X2 OR2X2_5630 ( .A(alu__abc_42281_new_n1807_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n1808_));
OR2X2 OR2X2_5631 ( .A(alu__abc_42281_new_n1726_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n1809_));
OR2X2 OR2X2_5632 ( .A(alu__abc_42281_new_n1810_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n1811_));
OR2X2 OR2X2_5633 ( .A(alu__abc_42281_new_n1813_), .B(alu__abc_42281_new_n1814_), .Y(alu__abc_42281_new_n1815_));
OR2X2 OR2X2_5634 ( .A(alu__abc_42281_new_n1819_), .B(alu__abc_42281_new_n1817_), .Y(alu__abc_42281_new_n1820_));
OR2X2 OR2X2_5635 ( .A(alu__abc_42281_new_n1823_), .B(alu__abc_42281_new_n1822_), .Y(alu__abc_42281_new_n1824_));
OR2X2 OR2X2_5636 ( .A(alu__abc_42281_new_n1824_), .B(alu__abc_42281_new_n1821_), .Y(alu__abc_42281_new_n1825_));
OR2X2 OR2X2_5637 ( .A(alu__abc_42281_new_n1820_), .B(alu__abc_42281_new_n1825_), .Y(alu__abc_42281_new_n1826_));
OR2X2 OR2X2_5638 ( .A(alu__abc_42281_new_n1816_), .B(alu__abc_42281_new_n1826_), .Y(alu__abc_42281_new_n1827_));
OR2X2 OR2X2_5639 ( .A(alu__abc_42281_new_n1827_), .B(alu__abc_42281_new_n1805_), .Y(alu__abc_42281_new_n1828_));
OR2X2 OR2X2_564 ( .A(_abc_44694_new_n2267_), .B(_abc_44694_new_n1400__bF_buf2), .Y(_abc_44694_new_n2268_));
OR2X2 OR2X2_5640 ( .A(alu__abc_42281_new_n1801_), .B(alu__abc_42281_new_n1828_), .Y(alu__abc_42281_new_n1829_));
OR2X2 OR2X2_5641 ( .A(alu__abc_42281_new_n1800_), .B(alu__abc_42281_new_n1829_), .Y(alu__abc_42281_new_n1830_));
OR2X2 OR2X2_5642 ( .A(alu__abc_42281_new_n1830_), .B(alu__abc_42281_new_n1795_), .Y(alu_p_o_16_));
OR2X2 OR2X2_5643 ( .A(alu__abc_42281_new_n807_), .B(alu__abc_42281_new_n690_), .Y(alu__abc_42281_new_n1838_));
OR2X2 OR2X2_5644 ( .A(alu__abc_42281_new_n1841_), .B(alu__abc_42281_new_n176_), .Y(alu__abc_42281_new_n1842_));
OR2X2 OR2X2_5645 ( .A(alu__abc_42281_new_n1843_), .B(alu__abc_42281_new_n177_), .Y(alu__abc_42281_new_n1844_));
OR2X2 OR2X2_5646 ( .A(alu__abc_42281_new_n1006_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n1848_));
OR2X2 OR2X2_5647 ( .A(alu__abc_42281_new_n1851_), .B(alu__abc_42281_new_n1852_), .Y(alu__abc_42281_new_n1853_));
OR2X2 OR2X2_5648 ( .A(alu__abc_42281_new_n1853_), .B(alu__abc_42281_new_n1854_), .Y(alu__abc_42281_new_n1855_));
OR2X2 OR2X2_5649 ( .A(alu__abc_42281_new_n1855_), .B(alu__abc_42281_new_n1850_), .Y(alu__abc_42281_new_n1856_));
OR2X2 OR2X2_565 ( .A(_abc_44694_new_n2239_), .B(_abc_44694_new_n1399__bF_buf1), .Y(_abc_44694_new_n2269_));
OR2X2 OR2X2_5650 ( .A(alu__abc_42281_new_n1857_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n1858_));
OR2X2 OR2X2_5651 ( .A(alu__abc_42281_new_n1771_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n1859_));
OR2X2 OR2X2_5652 ( .A(alu__abc_42281_new_n1860_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n1861_));
OR2X2 OR2X2_5653 ( .A(alu__abc_42281_new_n1684_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n1862_));
OR2X2 OR2X2_5654 ( .A(alu__abc_42281_new_n1865_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n1866_));
OR2X2 OR2X2_5655 ( .A(alu__abc_42281_new_n1866_), .B(alu__abc_42281_new_n1864_), .Y(alu__abc_42281_new_n1867_));
OR2X2 OR2X2_5656 ( .A(alu__abc_42281_new_n1074_), .B(alu__abc_42281_new_n271__bF_buf4), .Y(alu__abc_42281_new_n1868_));
OR2X2 OR2X2_5657 ( .A(alu__abc_42281_new_n1870_), .B(alu__abc_42281_new_n1856_), .Y(alu__abc_42281_new_n1871_));
OR2X2 OR2X2_5658 ( .A(alu__abc_42281_new_n1849_), .B(alu__abc_42281_new_n1871_), .Y(alu__abc_42281_new_n1872_));
OR2X2 OR2X2_5659 ( .A(alu__abc_42281_new_n1847_), .B(alu__abc_42281_new_n1872_), .Y(alu__abc_42281_new_n1873_));
OR2X2 OR2X2_566 ( .A(_abc_44694_new_n2270_), .B(_abc_44694_new_n1278__bF_buf2), .Y(_abc_44694_new_n2271_));
OR2X2 OR2X2_5660 ( .A(alu__abc_42281_new_n1846_), .B(alu__abc_42281_new_n1873_), .Y(alu__abc_42281_new_n1874_));
OR2X2 OR2X2_5661 ( .A(alu__abc_42281_new_n1874_), .B(alu__abc_42281_new_n1840_), .Y(alu_p_o_17_));
OR2X2 OR2X2_5662 ( .A(alu__abc_42281_new_n808_), .B(alu__abc_42281_new_n683_), .Y(alu__abc_42281_new_n1878_));
OR2X2 OR2X2_5663 ( .A(alu__abc_42281_new_n1881_), .B(alu__abc_42281_new_n454_), .Y(alu__abc_42281_new_n1882_));
OR2X2 OR2X2_5664 ( .A(alu__abc_42281_new_n1882_), .B(alu__abc_42281_new_n152_), .Y(alu__abc_42281_new_n1883_));
OR2X2 OR2X2_5665 ( .A(alu__abc_42281_new_n1103_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n1889_));
OR2X2 OR2X2_5666 ( .A(alu__abc_42281_new_n1891_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n1892_));
OR2X2 OR2X2_5667 ( .A(alu__abc_42281_new_n1807_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n1893_));
OR2X2 OR2X2_5668 ( .A(alu__abc_42281_new_n1894_), .B(alu_b_i_2_bF_buf0_), .Y(alu__abc_42281_new_n1895_));
OR2X2 OR2X2_5669 ( .A(alu__abc_42281_new_n1729_), .B(alu__abc_42281_new_n294__bF_buf6), .Y(alu__abc_42281_new_n1896_));
OR2X2 OR2X2_567 ( .A(_abc_44694_new_n2272_), .B(_abc_44694_new_n2273_), .Y(_abc_44694_new_n2274_));
OR2X2 OR2X2_5670 ( .A(alu__abc_42281_new_n1899_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n1900_));
OR2X2 OR2X2_5671 ( .A(alu__abc_42281_new_n1900_), .B(alu__abc_42281_new_n1898_), .Y(alu__abc_42281_new_n1901_));
OR2X2 OR2X2_5672 ( .A(alu__abc_42281_new_n1139_), .B(alu__abc_42281_new_n271__bF_buf3), .Y(alu__abc_42281_new_n1902_));
OR2X2 OR2X2_5673 ( .A(alu__abc_42281_new_n1908_), .B(alu__abc_42281_new_n1907_), .Y(alu__abc_42281_new_n1909_));
OR2X2 OR2X2_5674 ( .A(alu__abc_42281_new_n1909_), .B(alu__abc_42281_new_n1906_), .Y(alu__abc_42281_new_n1910_));
OR2X2 OR2X2_5675 ( .A(alu__abc_42281_new_n1910_), .B(alu__abc_42281_new_n1905_), .Y(alu__abc_42281_new_n1911_));
OR2X2 OR2X2_5676 ( .A(alu__abc_42281_new_n1904_), .B(alu__abc_42281_new_n1911_), .Y(alu__abc_42281_new_n1912_));
OR2X2 OR2X2_5677 ( .A(alu__abc_42281_new_n1912_), .B(alu__abc_42281_new_n1890_), .Y(alu__abc_42281_new_n1913_));
OR2X2 OR2X2_5678 ( .A(alu__abc_42281_new_n1888_), .B(alu__abc_42281_new_n1913_), .Y(alu__abc_42281_new_n1914_));
OR2X2 OR2X2_5679 ( .A(alu__abc_42281_new_n1887_), .B(alu__abc_42281_new_n1914_), .Y(alu__abc_42281_new_n1915_));
OR2X2 OR2X2_568 ( .A(_abc_44694_new_n1334__bF_buf0), .B(_abc_44694_new_n2274_), .Y(_abc_44694_new_n2275_));
OR2X2 OR2X2_5680 ( .A(alu__abc_42281_new_n1915_), .B(alu__abc_42281_new_n1880_), .Y(alu_p_o_18_));
OR2X2 OR2X2_5681 ( .A(alu__abc_42281_new_n809_), .B(alu__abc_42281_new_n681_), .Y(alu__abc_42281_new_n1917_));
OR2X2 OR2X2_5682 ( .A(alu__abc_42281_new_n1884_), .B(alu__abc_42281_new_n457_), .Y(alu__abc_42281_new_n1922_));
OR2X2 OR2X2_5683 ( .A(alu__abc_42281_new_n1922_), .B(alu__abc_42281_new_n160_), .Y(alu__abc_42281_new_n1923_));
OR2X2 OR2X2_5684 ( .A(alu__abc_42281_new_n1924_), .B(alu__abc_42281_new_n159_), .Y(alu__abc_42281_new_n1925_));
OR2X2 OR2X2_5685 ( .A(alu__abc_42281_new_n1929_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n1930_));
OR2X2 OR2X2_5686 ( .A(alu__abc_42281_new_n1857_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n1931_));
OR2X2 OR2X2_5687 ( .A(alu__abc_42281_new_n1932_), .B(alu_b_i_2_bF_buf6_), .Y(alu__abc_42281_new_n1933_));
OR2X2 OR2X2_5688 ( .A(alu__abc_42281_new_n1774_), .B(alu__abc_42281_new_n294__bF_buf5), .Y(alu__abc_42281_new_n1934_));
OR2X2 OR2X2_5689 ( .A(alu__abc_42281_new_n1937_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n1938_));
OR2X2 OR2X2_569 ( .A(_abc_44694_new_n2277_), .B(_abc_44694_new_n2241_), .Y(_abc_44694_new_n2278_));
OR2X2 OR2X2_5690 ( .A(alu__abc_42281_new_n1938_), .B(alu__abc_42281_new_n1936_), .Y(alu__abc_42281_new_n1939_));
OR2X2 OR2X2_5691 ( .A(alu__abc_42281_new_n1214_), .B(alu__abc_42281_new_n271__bF_buf2), .Y(alu__abc_42281_new_n1940_));
OR2X2 OR2X2_5692 ( .A(alu__abc_42281_new_n1177_), .B(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n1943_));
OR2X2 OR2X2_5693 ( .A(alu__abc_42281_new_n1948_), .B(alu__abc_42281_new_n1947_), .Y(alu__abc_42281_new_n1949_));
OR2X2 OR2X2_5694 ( .A(alu__abc_42281_new_n1949_), .B(alu__abc_42281_new_n1946_), .Y(alu__abc_42281_new_n1950_));
OR2X2 OR2X2_5695 ( .A(alu__abc_42281_new_n1950_), .B(alu__abc_42281_new_n1945_), .Y(alu__abc_42281_new_n1951_));
OR2X2 OR2X2_5696 ( .A(alu__abc_42281_new_n1944_), .B(alu__abc_42281_new_n1951_), .Y(alu__abc_42281_new_n1952_));
OR2X2 OR2X2_5697 ( .A(alu__abc_42281_new_n1952_), .B(alu__abc_42281_new_n1942_), .Y(alu__abc_42281_new_n1953_));
OR2X2 OR2X2_5698 ( .A(alu__abc_42281_new_n1928_), .B(alu__abc_42281_new_n1953_), .Y(alu__abc_42281_new_n1954_));
OR2X2 OR2X2_5699 ( .A(alu__abc_42281_new_n1927_), .B(alu__abc_42281_new_n1954_), .Y(alu__abc_42281_new_n1955_));
OR2X2 OR2X2_57 ( .A(_abc_44694_new_n797_), .B(_abc_44694_new_n800_), .Y(_abc_44694_new_n801_));
OR2X2 OR2X2_570 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(epc_q_24_), .Y(_abc_44694_new_n2279_));
OR2X2 OR2X2_5700 ( .A(alu__abc_42281_new_n1955_), .B(alu__abc_42281_new_n1921_), .Y(alu_p_o_19_));
OR2X2 OR2X2_5701 ( .A(alu__abc_42281_new_n810_), .B(alu__abc_42281_new_n673_), .Y(alu__abc_42281_new_n1957_));
OR2X2 OR2X2_5702 ( .A(alu__abc_42281_new_n1961_), .B(alu__abc_42281_new_n460_), .Y(alu__abc_42281_new_n1962_));
OR2X2 OR2X2_5703 ( .A(alu__abc_42281_new_n1962_), .B(alu__abc_42281_new_n117_), .Y(alu__abc_42281_new_n1965_));
OR2X2 OR2X2_5704 ( .A(alu__abc_42281_new_n1969_), .B(alu_b_i_1_bF_buf2_), .Y(alu__abc_42281_new_n1970_));
OR2X2 OR2X2_5705 ( .A(alu__abc_42281_new_n1891_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n1971_));
OR2X2 OR2X2_5706 ( .A(alu__abc_42281_new_n1972_), .B(alu_b_i_2_bF_buf5_), .Y(alu__abc_42281_new_n1973_));
OR2X2 OR2X2_5707 ( .A(alu__abc_42281_new_n1810_), .B(alu__abc_42281_new_n294__bF_buf4), .Y(alu__abc_42281_new_n1974_));
OR2X2 OR2X2_5708 ( .A(alu__abc_42281_new_n1977_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n1978_));
OR2X2 OR2X2_5709 ( .A(alu__abc_42281_new_n1978_), .B(alu__abc_42281_new_n1976_), .Y(alu__abc_42281_new_n1979_));
OR2X2 OR2X2_571 ( .A(_abc_44694_new_n2237_), .B(pc_q_25_), .Y(_abc_44694_new_n2282_));
OR2X2 OR2X2_5710 ( .A(alu__abc_42281_new_n1271_), .B(alu__abc_42281_new_n271__bF_buf1), .Y(alu__abc_42281_new_n1980_));
OR2X2 OR2X2_5711 ( .A(alu__abc_42281_new_n1259_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n1983_));
OR2X2 OR2X2_5712 ( .A(alu__abc_42281_new_n1986_), .B(alu__abc_42281_new_n1985_), .Y(alu__abc_42281_new_n1987_));
OR2X2 OR2X2_5713 ( .A(alu__abc_42281_new_n1988_), .B(alu__abc_42281_new_n1989_), .Y(alu__abc_42281_new_n1990_));
OR2X2 OR2X2_5714 ( .A(alu__abc_42281_new_n1990_), .B(alu__abc_42281_new_n1987_), .Y(alu__abc_42281_new_n1991_));
OR2X2 OR2X2_5715 ( .A(alu__abc_42281_new_n1984_), .B(alu__abc_42281_new_n1991_), .Y(alu__abc_42281_new_n1992_));
OR2X2 OR2X2_5716 ( .A(alu__abc_42281_new_n1992_), .B(alu__abc_42281_new_n1982_), .Y(alu__abc_42281_new_n1993_));
OR2X2 OR2X2_5717 ( .A(alu__abc_42281_new_n1968_), .B(alu__abc_42281_new_n1993_), .Y(alu__abc_42281_new_n1994_));
OR2X2 OR2X2_5718 ( .A(alu__abc_42281_new_n1967_), .B(alu__abc_42281_new_n1994_), .Y(alu__abc_42281_new_n1995_));
OR2X2 OR2X2_5719 ( .A(alu__abc_42281_new_n1960_), .B(alu__abc_42281_new_n1995_), .Y(alu_p_o_20_));
OR2X2 OR2X2_572 ( .A(_abc_44694_new_n2286_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n2287_));
OR2X2 OR2X2_5720 ( .A(alu__abc_42281_new_n811_), .B(alu__abc_42281_new_n658_), .Y(alu__abc_42281_new_n1997_));
OR2X2 OR2X2_5721 ( .A(alu__abc_42281_new_n2004_), .B(alu__abc_42281_new_n125_), .Y(alu__abc_42281_new_n2005_));
OR2X2 OR2X2_5722 ( .A(alu__abc_42281_new_n2003_), .B(alu__abc_42281_new_n124_), .Y(alu__abc_42281_new_n2006_));
OR2X2 OR2X2_5723 ( .A(alu__abc_42281_new_n1303_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n2010_));
OR2X2 OR2X2_5724 ( .A(alu__abc_42281_new_n2012_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n2013_));
OR2X2 OR2X2_5725 ( .A(alu__abc_42281_new_n1929_), .B(alu__abc_42281_new_n281__bF_buf3), .Y(alu__abc_42281_new_n2014_));
OR2X2 OR2X2_5726 ( .A(alu__abc_42281_new_n2015_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n2016_));
OR2X2 OR2X2_5727 ( .A(alu__abc_42281_new_n1860_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n2017_));
OR2X2 OR2X2_5728 ( .A(alu__abc_42281_new_n2020_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n2021_));
OR2X2 OR2X2_5729 ( .A(alu__abc_42281_new_n2021_), .B(alu__abc_42281_new_n2019_), .Y(alu__abc_42281_new_n2022_));
OR2X2 OR2X2_573 ( .A(opcode_q_23_), .B(pc_q_25_), .Y(_abc_44694_new_n2288_));
OR2X2 OR2X2_5730 ( .A(alu__abc_42281_new_n1324_), .B(alu__abc_42281_new_n271__bF_buf0), .Y(alu__abc_42281_new_n2023_));
OR2X2 OR2X2_5731 ( .A(alu__abc_42281_new_n2029_), .B(alu__abc_42281_new_n2028_), .Y(alu__abc_42281_new_n2030_));
OR2X2 OR2X2_5732 ( .A(alu__abc_42281_new_n2030_), .B(alu__abc_42281_new_n2027_), .Y(alu__abc_42281_new_n2031_));
OR2X2 OR2X2_5733 ( .A(alu__abc_42281_new_n2031_), .B(alu__abc_42281_new_n2026_), .Y(alu__abc_42281_new_n2032_));
OR2X2 OR2X2_5734 ( .A(alu__abc_42281_new_n2025_), .B(alu__abc_42281_new_n2032_), .Y(alu__abc_42281_new_n2033_));
OR2X2 OR2X2_5735 ( .A(alu__abc_42281_new_n2011_), .B(alu__abc_42281_new_n2033_), .Y(alu__abc_42281_new_n2034_));
OR2X2 OR2X2_5736 ( .A(alu__abc_42281_new_n2009_), .B(alu__abc_42281_new_n2034_), .Y(alu__abc_42281_new_n2035_));
OR2X2 OR2X2_5737 ( .A(alu__abc_42281_new_n2008_), .B(alu__abc_42281_new_n2035_), .Y(alu__abc_42281_new_n2036_));
OR2X2 OR2X2_5738 ( .A(alu__abc_42281_new_n2036_), .B(alu__abc_42281_new_n2002_), .Y(alu_p_o_21_));
OR2X2 OR2X2_5739 ( .A(alu__abc_42281_new_n2038_), .B(alu__abc_42281_new_n469_), .Y(alu__abc_42281_new_n2039_));
OR2X2 OR2X2_574 ( .A(_abc_44694_new_n2291_), .B(_abc_44694_new_n2255_), .Y(_abc_44694_new_n2292_));
OR2X2 OR2X2_5740 ( .A(alu__abc_42281_new_n2039_), .B(alu__abc_42281_new_n134_), .Y(alu__abc_42281_new_n2040_));
OR2X2 OR2X2_5741 ( .A(alu__abc_42281_new_n1999_), .B(alu__abc_42281_new_n664_), .Y(alu__abc_42281_new_n2045_));
OR2X2 OR2X2_5742 ( .A(alu__abc_42281_new_n2051_), .B(alu_b_i_1_bF_buf0_), .Y(alu__abc_42281_new_n2052_));
OR2X2 OR2X2_5743 ( .A(alu__abc_42281_new_n1969_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n2053_));
OR2X2 OR2X2_5744 ( .A(alu__abc_42281_new_n2054_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n2055_));
OR2X2 OR2X2_5745 ( .A(alu__abc_42281_new_n1894_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n2056_));
OR2X2 OR2X2_5746 ( .A(alu__abc_42281_new_n2059_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n2060_));
OR2X2 OR2X2_5747 ( .A(alu__abc_42281_new_n2060_), .B(alu__abc_42281_new_n2058_), .Y(alu__abc_42281_new_n2061_));
OR2X2 OR2X2_5748 ( .A(alu__abc_42281_new_n1374_), .B(alu__abc_42281_new_n271__bF_buf4), .Y(alu__abc_42281_new_n2062_));
OR2X2 OR2X2_5749 ( .A(alu__abc_42281_new_n1353_), .B(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n2065_));
OR2X2 OR2X2_575 ( .A(_abc_44694_new_n2259_), .B(_abc_44694_new_n2292_), .Y(_abc_44694_new_n2293_));
OR2X2 OR2X2_5750 ( .A(alu__abc_42281_new_n2068_), .B(alu__abc_42281_new_n2069_), .Y(alu__abc_42281_new_n2070_));
OR2X2 OR2X2_5751 ( .A(alu__abc_42281_new_n2070_), .B(alu__abc_42281_new_n2071_), .Y(alu__abc_42281_new_n2072_));
OR2X2 OR2X2_5752 ( .A(alu__abc_42281_new_n2072_), .B(alu__abc_42281_new_n2067_), .Y(alu__abc_42281_new_n2073_));
OR2X2 OR2X2_5753 ( .A(alu__abc_42281_new_n2066_), .B(alu__abc_42281_new_n2073_), .Y(alu__abc_42281_new_n2074_));
OR2X2 OR2X2_5754 ( .A(alu__abc_42281_new_n2074_), .B(alu__abc_42281_new_n2064_), .Y(alu__abc_42281_new_n2075_));
OR2X2 OR2X2_5755 ( .A(alu__abc_42281_new_n2050_), .B(alu__abc_42281_new_n2075_), .Y(alu__abc_42281_new_n2076_));
OR2X2 OR2X2_5756 ( .A(alu__abc_42281_new_n2049_), .B(alu__abc_42281_new_n2076_), .Y(alu__abc_42281_new_n2077_));
OR2X2 OR2X2_5757 ( .A(alu__abc_42281_new_n2077_), .B(alu__abc_42281_new_n2044_), .Y(alu_p_o_22_));
OR2X2 OR2X2_5758 ( .A(alu__abc_42281_new_n2046_), .B(alu__abc_42281_new_n820_), .Y(alu__abc_42281_new_n2079_));
OR2X2 OR2X2_5759 ( .A(alu__abc_42281_new_n2041_), .B(alu__abc_42281_new_n472_), .Y(alu__abc_42281_new_n2085_));
OR2X2 OR2X2_576 ( .A(_abc_44694_new_n2301_), .B(_abc_44694_new_n2302_), .Y(_abc_44694_new_n2303_));
OR2X2 OR2X2_5760 ( .A(alu__abc_42281_new_n2086_), .B(alu__abc_42281_new_n141_), .Y(alu__abc_42281_new_n2087_));
OR2X2 OR2X2_5761 ( .A(alu__abc_42281_new_n2085_), .B(alu__abc_42281_new_n142_), .Y(alu__abc_42281_new_n2088_));
OR2X2 OR2X2_5762 ( .A(alu__abc_42281_new_n2092_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n2093_));
OR2X2 OR2X2_5763 ( .A(alu__abc_42281_new_n2012_), .B(alu__abc_42281_new_n281__bF_buf1), .Y(alu__abc_42281_new_n2094_));
OR2X2 OR2X2_5764 ( .A(alu__abc_42281_new_n2095_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n2096_));
OR2X2 OR2X2_5765 ( .A(alu__abc_42281_new_n1932_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n2097_));
OR2X2 OR2X2_5766 ( .A(alu__abc_42281_new_n2100_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n2101_));
OR2X2 OR2X2_5767 ( .A(alu__abc_42281_new_n2101_), .B(alu__abc_42281_new_n2099_), .Y(alu__abc_42281_new_n2102_));
OR2X2 OR2X2_5768 ( .A(alu__abc_42281_new_n1426_), .B(alu__abc_42281_new_n271__bF_buf3), .Y(alu__abc_42281_new_n2103_));
OR2X2 OR2X2_5769 ( .A(alu__abc_42281_new_n1405_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n2106_));
OR2X2 OR2X2_577 ( .A(_abc_44694_new_n2304_), .B(_abc_44694_new_n2305_), .Y(_abc_44694_new_n2306_));
OR2X2 OR2X2_5770 ( .A(alu__abc_42281_new_n2109_), .B(alu__abc_42281_new_n2110_), .Y(alu__abc_42281_new_n2111_));
OR2X2 OR2X2_5771 ( .A(alu__abc_42281_new_n2111_), .B(alu__abc_42281_new_n2112_), .Y(alu__abc_42281_new_n2113_));
OR2X2 OR2X2_5772 ( .A(alu__abc_42281_new_n2113_), .B(alu__abc_42281_new_n2108_), .Y(alu__abc_42281_new_n2114_));
OR2X2 OR2X2_5773 ( .A(alu__abc_42281_new_n2107_), .B(alu__abc_42281_new_n2114_), .Y(alu__abc_42281_new_n2115_));
OR2X2 OR2X2_5774 ( .A(alu__abc_42281_new_n2115_), .B(alu__abc_42281_new_n2105_), .Y(alu__abc_42281_new_n2116_));
OR2X2 OR2X2_5775 ( .A(alu__abc_42281_new_n2091_), .B(alu__abc_42281_new_n2116_), .Y(alu__abc_42281_new_n2117_));
OR2X2 OR2X2_5776 ( .A(alu__abc_42281_new_n2090_), .B(alu__abc_42281_new_n2117_), .Y(alu__abc_42281_new_n2118_));
OR2X2 OR2X2_5777 ( .A(alu__abc_42281_new_n2118_), .B(alu__abc_42281_new_n2084_), .Y(alu_p_o_23_));
OR2X2 OR2X2_5778 ( .A(alu__abc_42281_new_n2120_), .B(alu__abc_42281_new_n650_), .Y(alu__abc_42281_new_n2121_));
OR2X2 OR2X2_5779 ( .A(alu__abc_42281_new_n477_), .B(alu__abc_42281_new_n196_), .Y(alu__abc_42281_new_n2126_));
OR2X2 OR2X2_578 ( .A(_abc_44694_new_n2306_), .B(_abc_44694_new_n1400__bF_buf1), .Y(_abc_44694_new_n2307_));
OR2X2 OR2X2_5780 ( .A(alu__abc_42281_new_n2127_), .B(alu__abc_42281_new_n195_), .Y(alu__abc_42281_new_n2128_));
OR2X2 OR2X2_5781 ( .A(alu__abc_42281_new_n1452_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n2132_));
OR2X2 OR2X2_5782 ( .A(alu__abc_42281_new_n1812_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n2135_));
OR2X2 OR2X2_5783 ( .A(alu__abc_42281_new_n2136_), .B(alu_b_i_1_bF_buf6_), .Y(alu__abc_42281_new_n2137_));
OR2X2 OR2X2_5784 ( .A(alu__abc_42281_new_n2051_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n2138_));
OR2X2 OR2X2_5785 ( .A(alu__abc_42281_new_n2139_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n2140_));
OR2X2 OR2X2_5786 ( .A(alu__abc_42281_new_n1972_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n2141_));
OR2X2 OR2X2_5787 ( .A(alu__abc_42281_new_n2142_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n2143_));
OR2X2 OR2X2_5788 ( .A(alu__abc_42281_new_n2148_), .B(alu__abc_42281_new_n2149_), .Y(alu__abc_42281_new_n2150_));
OR2X2 OR2X2_5789 ( .A(alu__abc_42281_new_n2150_), .B(alu__abc_42281_new_n2147_), .Y(alu__abc_42281_new_n2151_));
OR2X2 OR2X2_579 ( .A(_abc_44694_new_n2285_), .B(_abc_44694_new_n1399__bF_buf0), .Y(_abc_44694_new_n2308_));
OR2X2 OR2X2_5790 ( .A(alu__abc_42281_new_n2151_), .B(alu__abc_42281_new_n2146_), .Y(alu__abc_42281_new_n2152_));
OR2X2 OR2X2_5791 ( .A(alu__abc_42281_new_n2145_), .B(alu__abc_42281_new_n2152_), .Y(alu__abc_42281_new_n2153_));
OR2X2 OR2X2_5792 ( .A(alu__abc_42281_new_n2153_), .B(alu__abc_42281_new_n2134_), .Y(alu__abc_42281_new_n2154_));
OR2X2 OR2X2_5793 ( .A(alu__abc_42281_new_n2154_), .B(alu__abc_42281_new_n2133_), .Y(alu__abc_42281_new_n2155_));
OR2X2 OR2X2_5794 ( .A(alu__abc_42281_new_n2131_), .B(alu__abc_42281_new_n2155_), .Y(alu__abc_42281_new_n2156_));
OR2X2 OR2X2_5795 ( .A(alu__abc_42281_new_n2130_), .B(alu__abc_42281_new_n2156_), .Y(alu__abc_42281_new_n2157_));
OR2X2 OR2X2_5796 ( .A(alu__abc_42281_new_n2125_), .B(alu__abc_42281_new_n2157_), .Y(alu_p_o_24_));
OR2X2 OR2X2_5797 ( .A(alu__abc_42281_new_n2122_), .B(alu__abc_42281_new_n671_), .Y(alu__abc_42281_new_n2161_));
OR2X2 OR2X2_5798 ( .A(alu__abc_42281_new_n2165_), .B(alu__abc_42281_new_n188_), .Y(alu__abc_42281_new_n2166_));
OR2X2 OR2X2_5799 ( .A(alu__abc_42281_new_n2164_), .B(alu__abc_42281_new_n187_), .Y(alu__abc_42281_new_n2167_));
OR2X2 OR2X2_58 ( .A(_abc_44694_new_n673__bF_buf2), .B(_abc_44694_new_n801_), .Y(_abc_44694_new_n802_));
OR2X2 OR2X2_580 ( .A(_abc_44694_new_n2309_), .B(_abc_44694_new_n1278__bF_buf1), .Y(_abc_44694_new_n2310_));
OR2X2 OR2X2_5800 ( .A(alu__abc_42281_new_n1495_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n2171_));
OR2X2 OR2X2_5801 ( .A(alu__abc_42281_new_n2174_), .B(alu_b_i_1_bF_buf5_), .Y(alu__abc_42281_new_n2175_));
OR2X2 OR2X2_5802 ( .A(alu__abc_42281_new_n2092_), .B(alu__abc_42281_new_n281__bF_buf6), .Y(alu__abc_42281_new_n2176_));
OR2X2 OR2X2_5803 ( .A(alu__abc_42281_new_n2179_), .B(alu_b_i_3_bF_buf3_), .Y(alu__abc_42281_new_n2180_));
OR2X2 OR2X2_5804 ( .A(alu__abc_42281_new_n2180_), .B(alu__abc_42281_new_n2178_), .Y(alu__abc_42281_new_n2181_));
OR2X2 OR2X2_5805 ( .A(alu__abc_42281_new_n1863_), .B(alu__abc_42281_new_n299__bF_buf3), .Y(alu__abc_42281_new_n2182_));
OR2X2 OR2X2_5806 ( .A(alu__abc_42281_new_n2187_), .B(alu__abc_42281_new_n2188_), .Y(alu__abc_42281_new_n2189_));
OR2X2 OR2X2_5807 ( .A(alu__abc_42281_new_n2189_), .B(alu__abc_42281_new_n2186_), .Y(alu__abc_42281_new_n2190_));
OR2X2 OR2X2_5808 ( .A(alu__abc_42281_new_n2190_), .B(alu__abc_42281_new_n2185_), .Y(alu__abc_42281_new_n2191_));
OR2X2 OR2X2_5809 ( .A(alu__abc_42281_new_n2184_), .B(alu__abc_42281_new_n2191_), .Y(alu__abc_42281_new_n2192_));
OR2X2 OR2X2_581 ( .A(_abc_44694_new_n2311_), .B(_abc_44694_new_n2312_), .Y(_abc_44694_new_n2313_));
OR2X2 OR2X2_5810 ( .A(alu__abc_42281_new_n2192_), .B(alu__abc_42281_new_n2173_), .Y(alu__abc_42281_new_n2193_));
OR2X2 OR2X2_5811 ( .A(alu__abc_42281_new_n2172_), .B(alu__abc_42281_new_n2193_), .Y(alu__abc_42281_new_n2194_));
OR2X2 OR2X2_5812 ( .A(alu__abc_42281_new_n2170_), .B(alu__abc_42281_new_n2194_), .Y(alu__abc_42281_new_n2195_));
OR2X2 OR2X2_5813 ( .A(alu__abc_42281_new_n2169_), .B(alu__abc_42281_new_n2195_), .Y(alu__abc_42281_new_n2196_));
OR2X2 OR2X2_5814 ( .A(alu__abc_42281_new_n2163_), .B(alu__abc_42281_new_n2196_), .Y(alu_p_o_25_));
OR2X2 OR2X2_5815 ( .A(alu__abc_42281_new_n2159_), .B(alu__abc_42281_new_n815_), .Y(alu__abc_42281_new_n2198_));
OR2X2 OR2X2_5816 ( .A(alu__abc_42281_new_n2205_), .B(alu__abc_42281_new_n485_), .Y(alu__abc_42281_new_n2206_));
OR2X2 OR2X2_5817 ( .A(alu__abc_42281_new_n2206_), .B(alu__abc_42281_new_n204_), .Y(alu__abc_42281_new_n2207_));
OR2X2 OR2X2_5818 ( .A(alu__abc_42281_new_n2208_), .B(alu__abc_42281_new_n205_), .Y(alu__abc_42281_new_n2209_));
OR2X2 OR2X2_5819 ( .A(alu__abc_42281_new_n1541_), .B(alu_b_i_4_bF_buf5_), .Y(alu__abc_42281_new_n2213_));
OR2X2 OR2X2_582 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n2313_), .Y(_abc_44694_new_n2314_));
OR2X2 OR2X2_5820 ( .A(alu__abc_42281_new_n2215_), .B(alu_b_i_1_bF_buf4_), .Y(alu__abc_42281_new_n2216_));
OR2X2 OR2X2_5821 ( .A(alu__abc_42281_new_n2136_), .B(alu__abc_42281_new_n281__bF_buf5), .Y(alu__abc_42281_new_n2217_));
OR2X2 OR2X2_5822 ( .A(alu__abc_42281_new_n2220_), .B(alu_b_i_3_bF_buf2_), .Y(alu__abc_42281_new_n2221_));
OR2X2 OR2X2_5823 ( .A(alu__abc_42281_new_n2221_), .B(alu__abc_42281_new_n2219_), .Y(alu__abc_42281_new_n2222_));
OR2X2 OR2X2_5824 ( .A(alu__abc_42281_new_n1897_), .B(alu__abc_42281_new_n299__bF_buf2), .Y(alu__abc_42281_new_n2223_));
OR2X2 OR2X2_5825 ( .A(alu__abc_42281_new_n2230_), .B(alu__abc_42281_new_n2229_), .Y(alu__abc_42281_new_n2231_));
OR2X2 OR2X2_5826 ( .A(alu__abc_42281_new_n2231_), .B(alu__abc_42281_new_n2228_), .Y(alu__abc_42281_new_n2232_));
OR2X2 OR2X2_5827 ( .A(alu__abc_42281_new_n2232_), .B(alu__abc_42281_new_n2227_), .Y(alu__abc_42281_new_n2233_));
OR2X2 OR2X2_5828 ( .A(alu__abc_42281_new_n2226_), .B(alu__abc_42281_new_n2233_), .Y(alu__abc_42281_new_n2234_));
OR2X2 OR2X2_5829 ( .A(alu__abc_42281_new_n2234_), .B(alu__abc_42281_new_n2225_), .Y(alu__abc_42281_new_n2235_));
OR2X2 OR2X2_583 ( .A(_abc_44694_new_n2316_), .B(_abc_44694_new_n2287_), .Y(_abc_44694_new_n2317_));
OR2X2 OR2X2_5830 ( .A(alu__abc_42281_new_n2235_), .B(alu__abc_42281_new_n2214_), .Y(alu__abc_42281_new_n2236_));
OR2X2 OR2X2_5831 ( .A(alu__abc_42281_new_n2212_), .B(alu__abc_42281_new_n2236_), .Y(alu__abc_42281_new_n2237_));
OR2X2 OR2X2_5832 ( .A(alu__abc_42281_new_n2211_), .B(alu__abc_42281_new_n2237_), .Y(alu__abc_42281_new_n2238_));
OR2X2 OR2X2_5833 ( .A(alu__abc_42281_new_n2204_), .B(alu__abc_42281_new_n2238_), .Y(alu_p_o_26_));
OR2X2 OR2X2_5834 ( .A(alu__abc_42281_new_n2240_), .B(alu__abc_42281_new_n646_), .Y(alu__abc_42281_new_n2241_));
OR2X2 OR2X2_5835 ( .A(alu__abc_42281_new_n2249_), .B(alu__abc_42281_new_n213_), .Y(alu__abc_42281_new_n2250_));
OR2X2 OR2X2_5836 ( .A(alu__abc_42281_new_n2248_), .B(alu__abc_42281_new_n212_), .Y(alu__abc_42281_new_n2251_));
OR2X2 OR2X2_5837 ( .A(alu__abc_42281_new_n1583_), .B(alu_b_i_4_bF_buf4_), .Y(alu__abc_42281_new_n2254_));
OR2X2 OR2X2_5838 ( .A(alu__abc_42281_new_n2259_), .B(alu__abc_42281_new_n2258_), .Y(alu__abc_42281_new_n2260_));
OR2X2 OR2X2_5839 ( .A(alu__abc_42281_new_n2260_), .B(alu__abc_42281_new_n2261_), .Y(alu__abc_42281_new_n2262_));
OR2X2 OR2X2_584 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(epc_q_25_), .Y(_abc_44694_new_n2318_));
OR2X2 OR2X2_5840 ( .A(alu__abc_42281_new_n2262_), .B(alu__abc_42281_new_n2257_), .Y(alu__abc_42281_new_n2263_));
OR2X2 OR2X2_5841 ( .A(alu__abc_42281_new_n1935_), .B(alu__abc_42281_new_n299__bF_buf1), .Y(alu__abc_42281_new_n2264_));
OR2X2 OR2X2_5842 ( .A(alu__abc_42281_new_n2265_), .B(alu_b_i_1_bF_buf3_), .Y(alu__abc_42281_new_n2266_));
OR2X2 OR2X2_5843 ( .A(alu__abc_42281_new_n2174_), .B(alu__abc_42281_new_n281__bF_buf4), .Y(alu__abc_42281_new_n2267_));
OR2X2 OR2X2_5844 ( .A(alu__abc_42281_new_n2270_), .B(alu_b_i_3_bF_buf1_), .Y(alu__abc_42281_new_n2271_));
OR2X2 OR2X2_5845 ( .A(alu__abc_42281_new_n2271_), .B(alu__abc_42281_new_n2269_), .Y(alu__abc_42281_new_n2272_));
OR2X2 OR2X2_5846 ( .A(alu__abc_42281_new_n2274_), .B(alu__abc_42281_new_n2263_), .Y(alu__abc_42281_new_n2275_));
OR2X2 OR2X2_5847 ( .A(alu__abc_42281_new_n2275_), .B(alu__abc_42281_new_n2256_), .Y(alu__abc_42281_new_n2276_));
OR2X2 OR2X2_5848 ( .A(alu__abc_42281_new_n2276_), .B(alu__abc_42281_new_n2255_), .Y(alu__abc_42281_new_n2277_));
OR2X2 OR2X2_5849 ( .A(alu__abc_42281_new_n2253_), .B(alu__abc_42281_new_n2277_), .Y(alu__abc_42281_new_n2278_));
OR2X2 OR2X2_585 ( .A(_abc_44694_new_n2283_), .B(pc_q_26_), .Y(_abc_44694_new_n2321_));
OR2X2 OR2X2_5850 ( .A(alu__abc_42281_new_n2278_), .B(alu__abc_42281_new_n2246_), .Y(alu__abc_42281_new_n2279_));
OR2X2 OR2X2_5851 ( .A(alu__abc_42281_new_n2279_), .B(alu__abc_42281_new_n2245_), .Y(alu_p_o_27_));
OR2X2 OR2X2_5852 ( .A(alu__abc_42281_new_n2242_), .B(alu__abc_42281_new_n639_), .Y(alu__abc_42281_new_n2281_));
OR2X2 OR2X2_5853 ( .A(alu__abc_42281_new_n495_), .B(alu__abc_42281_new_n223_), .Y(alu__abc_42281_new_n2286_));
OR2X2 OR2X2_5854 ( .A(alu__abc_42281_new_n1632_), .B(alu_b_i_4_bF_buf3_), .Y(alu__abc_42281_new_n2292_));
OR2X2 OR2X2_5855 ( .A(alu__abc_42281_new_n1975_), .B(alu__abc_42281_new_n299__bF_buf0), .Y(alu__abc_42281_new_n2294_));
OR2X2 OR2X2_5856 ( .A(alu__abc_42281_new_n2297_), .B(alu_b_i_2_bF_buf4_), .Y(alu__abc_42281_new_n2298_));
OR2X2 OR2X2_5857 ( .A(alu__abc_42281_new_n2298_), .B(alu__abc_42281_new_n2296_), .Y(alu__abc_42281_new_n2299_));
OR2X2 OR2X2_5858 ( .A(alu__abc_42281_new_n2139_), .B(alu__abc_42281_new_n294__bF_buf3), .Y(alu__abc_42281_new_n2300_));
OR2X2 OR2X2_5859 ( .A(alu__abc_42281_new_n2301_), .B(alu_b_i_3_bF_buf0_), .Y(alu__abc_42281_new_n2302_));
OR2X2 OR2X2_586 ( .A(_abc_44694_new_n2325_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n2326_));
OR2X2 OR2X2_5860 ( .A(alu__abc_42281_new_n2308_), .B(alu__abc_42281_new_n2309_), .Y(alu__abc_42281_new_n2310_));
OR2X2 OR2X2_5861 ( .A(alu__abc_42281_new_n2310_), .B(alu__abc_42281_new_n2307_), .Y(alu__abc_42281_new_n2311_));
OR2X2 OR2X2_5862 ( .A(alu__abc_42281_new_n2311_), .B(alu__abc_42281_new_n2306_), .Y(alu__abc_42281_new_n2312_));
OR2X2 OR2X2_5863 ( .A(alu__abc_42281_new_n2305_), .B(alu__abc_42281_new_n2312_), .Y(alu__abc_42281_new_n2313_));
OR2X2 OR2X2_5864 ( .A(alu__abc_42281_new_n2313_), .B(alu__abc_42281_new_n2304_), .Y(alu__abc_42281_new_n2314_));
OR2X2 OR2X2_5865 ( .A(alu__abc_42281_new_n2314_), .B(alu__abc_42281_new_n2293_), .Y(alu__abc_42281_new_n2315_));
OR2X2 OR2X2_5866 ( .A(alu__abc_42281_new_n2291_), .B(alu__abc_42281_new_n2315_), .Y(alu__abc_42281_new_n2316_));
OR2X2 OR2X2_5867 ( .A(alu__abc_42281_new_n2290_), .B(alu__abc_42281_new_n2316_), .Y(alu__abc_42281_new_n2317_));
OR2X2 OR2X2_5868 ( .A(alu__abc_42281_new_n2285_), .B(alu__abc_42281_new_n2317_), .Y(alu_p_o_28_));
OR2X2 OR2X2_5869 ( .A(alu__abc_42281_new_n2319_), .B(alu__abc_42281_new_n637_), .Y(alu__abc_42281_new_n2320_));
OR2X2 OR2X2_587 ( .A(_abc_44694_new_n2295_), .B(_abc_44694_new_n2328_), .Y(_abc_44694_new_n2329_));
OR2X2 OR2X2_5870 ( .A(alu__abc_42281_new_n2325_), .B(alu__abc_42281_new_n230_), .Y(alu__abc_42281_new_n2326_));
OR2X2 OR2X2_5871 ( .A(alu__abc_42281_new_n2327_), .B(alu__abc_42281_new_n231_), .Y(alu__abc_42281_new_n2328_));
OR2X2 OR2X2_5872 ( .A(alu__abc_42281_new_n1672_), .B(alu_b_i_4_bF_buf2_), .Y(alu__abc_42281_new_n2332_));
OR2X2 OR2X2_5873 ( .A(alu_a_i_29_), .B(alu_b_i_0_bF_buf1_), .Y(alu__abc_42281_new_n2335_));
OR2X2 OR2X2_5874 ( .A(alu__abc_42281_new_n2336_), .B(alu_b_i_1_bF_buf1_), .Y(alu__abc_42281_new_n2337_));
OR2X2 OR2X2_5875 ( .A(alu__abc_42281_new_n2265_), .B(alu__abc_42281_new_n281__bF_buf2), .Y(alu__abc_42281_new_n2338_));
OR2X2 OR2X2_5876 ( .A(alu__abc_42281_new_n2339_), .B(alu_b_i_2_bF_buf3_), .Y(alu__abc_42281_new_n2340_));
OR2X2 OR2X2_5877 ( .A(alu__abc_42281_new_n2177_), .B(alu__abc_42281_new_n294__bF_buf2), .Y(alu__abc_42281_new_n2341_));
OR2X2 OR2X2_5878 ( .A(alu__abc_42281_new_n2342_), .B(alu_b_i_3_bF_buf6_), .Y(alu__abc_42281_new_n2343_));
OR2X2 OR2X2_5879 ( .A(alu__abc_42281_new_n2018_), .B(alu__abc_42281_new_n299__bF_buf6), .Y(alu__abc_42281_new_n2344_));
OR2X2 OR2X2_588 ( .A(opcode_q_24_), .B(pc_q_26_), .Y(_abc_44694_new_n2330_));
OR2X2 OR2X2_5880 ( .A(alu__abc_42281_new_n2349_), .B(alu__abc_42281_new_n2350_), .Y(alu__abc_42281_new_n2351_));
OR2X2 OR2X2_5881 ( .A(alu__abc_42281_new_n2351_), .B(alu__abc_42281_new_n2348_), .Y(alu__abc_42281_new_n2352_));
OR2X2 OR2X2_5882 ( .A(alu__abc_42281_new_n2352_), .B(alu__abc_42281_new_n2347_), .Y(alu__abc_42281_new_n2353_));
OR2X2 OR2X2_5883 ( .A(alu__abc_42281_new_n2346_), .B(alu__abc_42281_new_n2353_), .Y(alu__abc_42281_new_n2354_));
OR2X2 OR2X2_5884 ( .A(alu__abc_42281_new_n2354_), .B(alu__abc_42281_new_n2334_), .Y(alu__abc_42281_new_n2355_));
OR2X2 OR2X2_5885 ( .A(alu__abc_42281_new_n2333_), .B(alu__abc_42281_new_n2355_), .Y(alu__abc_42281_new_n2356_));
OR2X2 OR2X2_5886 ( .A(alu__abc_42281_new_n2331_), .B(alu__abc_42281_new_n2356_), .Y(alu__abc_42281_new_n2357_));
OR2X2 OR2X2_5887 ( .A(alu__abc_42281_new_n2330_), .B(alu__abc_42281_new_n2357_), .Y(alu__abc_42281_new_n2358_));
OR2X2 OR2X2_5888 ( .A(alu__abc_42281_new_n2324_), .B(alu__abc_42281_new_n2358_), .Y(alu_p_o_29_));
OR2X2 OR2X2_5889 ( .A(alu__abc_42281_new_n2321_), .B(alu__abc_42281_new_n630_), .Y(alu__abc_42281_new_n2362_));
OR2X2 OR2X2_589 ( .A(_abc_44694_new_n2329_), .B(_abc_44694_new_n2333_), .Y(_abc_44694_new_n2334_));
OR2X2 OR2X2_5890 ( .A(alu__abc_42281_new_n505_), .B(alu__abc_42281_new_n240_), .Y(alu__abc_42281_new_n2365_));
OR2X2 OR2X2_5891 ( .A(alu__abc_42281_new_n1718_), .B(alu_b_i_4_bF_buf1_), .Y(alu__abc_42281_new_n2370_));
OR2X2 OR2X2_5892 ( .A(alu__abc_42281_new_n2374_), .B(alu_b_i_2_bF_buf2_), .Y(alu__abc_42281_new_n2375_));
OR2X2 OR2X2_5893 ( .A(alu__abc_42281_new_n2375_), .B(alu__abc_42281_new_n2373_), .Y(alu__abc_42281_new_n2376_));
OR2X2 OR2X2_5894 ( .A(alu__abc_42281_new_n2218_), .B(alu__abc_42281_new_n294__bF_buf1), .Y(alu__abc_42281_new_n2377_));
OR2X2 OR2X2_5895 ( .A(alu__abc_42281_new_n2378_), .B(alu_b_i_3_bF_buf5_), .Y(alu__abc_42281_new_n2379_));
OR2X2 OR2X2_5896 ( .A(alu__abc_42281_new_n2057_), .B(alu__abc_42281_new_n299__bF_buf5), .Y(alu__abc_42281_new_n2380_));
OR2X2 OR2X2_5897 ( .A(alu__abc_42281_new_n2387_), .B(alu__abc_42281_new_n2386_), .Y(alu__abc_42281_new_n2388_));
OR2X2 OR2X2_5898 ( .A(alu__abc_42281_new_n2388_), .B(alu__abc_42281_new_n2385_), .Y(alu__abc_42281_new_n2389_));
OR2X2 OR2X2_5899 ( .A(alu__abc_42281_new_n2389_), .B(alu__abc_42281_new_n2384_), .Y(alu__abc_42281_new_n2390_));
OR2X2 OR2X2_59 ( .A(_abc_44694_new_n804_), .B(_abc_44694_new_n803_), .Y(_abc_44694_new_n805_));
OR2X2 OR2X2_590 ( .A(_abc_44694_new_n2338_), .B(_abc_44694_new_n2339_), .Y(_abc_44694_new_n2340_));
OR2X2 OR2X2_5900 ( .A(alu__abc_42281_new_n2383_), .B(alu__abc_42281_new_n2390_), .Y(alu__abc_42281_new_n2391_));
OR2X2 OR2X2_5901 ( .A(alu__abc_42281_new_n2391_), .B(alu__abc_42281_new_n2382_), .Y(alu__abc_42281_new_n2392_));
OR2X2 OR2X2_5902 ( .A(alu__abc_42281_new_n2392_), .B(alu__abc_42281_new_n2371_), .Y(alu__abc_42281_new_n2393_));
OR2X2 OR2X2_5903 ( .A(alu__abc_42281_new_n2369_), .B(alu__abc_42281_new_n2393_), .Y(alu__abc_42281_new_n2394_));
OR2X2 OR2X2_5904 ( .A(alu__abc_42281_new_n2368_), .B(alu__abc_42281_new_n2394_), .Y(alu__abc_42281_new_n2395_));
OR2X2 OR2X2_5905 ( .A(alu__abc_42281_new_n2364_), .B(alu__abc_42281_new_n2395_), .Y(alu_p_o_30_));
OR2X2 OR2X2_5906 ( .A(alu__abc_42281_new_n2360_), .B(alu__abc_42281_new_n628_), .Y(alu__abc_42281_new_n2397_));
OR2X2 OR2X2_5907 ( .A(alu__abc_42281_new_n509_), .B(alu__abc_42281_new_n512_), .Y(alu__abc_42281_new_n2402_));
OR2X2 OR2X2_5908 ( .A(alu__abc_42281_new_n508_), .B(alu__abc_42281_new_n245_), .Y(alu__abc_42281_new_n2403_));
OR2X2 OR2X2_5909 ( .A(alu__abc_42281_new_n1762_), .B(alu_b_i_4_bF_buf0_), .Y(alu__abc_42281_new_n2406_));
OR2X2 OR2X2_591 ( .A(_abc_44694_new_n2341_), .B(_abc_44694_new_n2342_), .Y(_abc_44694_new_n2343_));
OR2X2 OR2X2_5910 ( .A(alu__abc_42281_new_n963_), .B(alu__abc_42281_new_n966_), .Y(alu__abc_42281_new_n2408_));
OR2X2 OR2X2_5911 ( .A(alu__abc_42281_new_n2408_), .B(alu_b_i_1_bF_buf7_), .Y(alu__abc_42281_new_n2409_));
OR2X2 OR2X2_5912 ( .A(alu__abc_42281_new_n2336_), .B(alu__abc_42281_new_n281__bF_buf0), .Y(alu__abc_42281_new_n2410_));
OR2X2 OR2X2_5913 ( .A(alu__abc_42281_new_n2411_), .B(alu_b_i_2_bF_buf1_), .Y(alu__abc_42281_new_n2412_));
OR2X2 OR2X2_5914 ( .A(alu__abc_42281_new_n2268_), .B(alu__abc_42281_new_n294__bF_buf0), .Y(alu__abc_42281_new_n2413_));
OR2X2 OR2X2_5915 ( .A(alu__abc_42281_new_n2414_), .B(alu_b_i_3_bF_buf4_), .Y(alu__abc_42281_new_n2415_));
OR2X2 OR2X2_5916 ( .A(alu__abc_42281_new_n2098_), .B(alu__abc_42281_new_n299__bF_buf4), .Y(alu__abc_42281_new_n2416_));
OR2X2 OR2X2_5917 ( .A(alu__abc_42281_new_n2423_), .B(alu__abc_42281_new_n2422_), .Y(alu__abc_42281_new_n2424_));
OR2X2 OR2X2_5918 ( .A(alu__abc_42281_new_n2424_), .B(alu__abc_42281_new_n2421_), .Y(alu__abc_42281_new_n2425_));
OR2X2 OR2X2_5919 ( .A(alu__abc_42281_new_n2425_), .B(alu__abc_42281_new_n2420_), .Y(alu__abc_42281_new_n2426_));
OR2X2 OR2X2_592 ( .A(_abc_44694_new_n2343_), .B(_abc_44694_new_n1400__bF_buf0), .Y(_abc_44694_new_n2344_));
OR2X2 OR2X2_5920 ( .A(alu__abc_42281_new_n2419_), .B(alu__abc_42281_new_n2426_), .Y(alu__abc_42281_new_n2427_));
OR2X2 OR2X2_5921 ( .A(alu__abc_42281_new_n2427_), .B(alu__abc_42281_new_n2418_), .Y(alu__abc_42281_new_n2428_));
OR2X2 OR2X2_5922 ( .A(alu__abc_42281_new_n2428_), .B(alu__abc_42281_new_n2407_), .Y(alu__abc_42281_new_n2429_));
OR2X2 OR2X2_5923 ( .A(alu__abc_42281_new_n2405_), .B(alu__abc_42281_new_n2429_), .Y(alu__abc_42281_new_n2430_));
OR2X2 OR2X2_5924 ( .A(alu__abc_42281_new_n2430_), .B(alu__abc_42281_new_n2401_), .Y(alu__abc_42281_new_n2431_));
OR2X2 OR2X2_5925 ( .A(alu__abc_42281_new_n2400_), .B(alu__abc_42281_new_n2431_), .Y(alu_p_o_31_));
OR2X2 OR2X2_5926 ( .A(alu__abc_42281_new_n931_), .B(alu_a_i_1_), .Y(alu__abc_42281_new_n2436_));
OR2X2 OR2X2_5927 ( .A(alu__abc_42281_new_n2441_), .B(alu__abc_42281_new_n397_), .Y(alu__abc_42281_new_n2442_));
OR2X2 OR2X2_5928 ( .A(alu__abc_42281_new_n2439_), .B(alu__abc_42281_new_n2442_), .Y(alu__abc_42281_new_n2443_));
OR2X2 OR2X2_5929 ( .A(alu__abc_42281_new_n2446_), .B(alu__abc_42281_new_n389_), .Y(alu__abc_42281_new_n2447_));
OR2X2 OR2X2_593 ( .A(_abc_44694_new_n2324_), .B(_abc_44694_new_n1399__bF_buf4), .Y(_abc_44694_new_n2345_));
OR2X2 OR2X2_5930 ( .A(alu__abc_42281_new_n2449_), .B(alu__abc_42281_new_n393_), .Y(alu__abc_42281_new_n2450_));
OR2X2 OR2X2_5931 ( .A(alu__abc_42281_new_n2451_), .B(alu__abc_42281_new_n2447_), .Y(alu__abc_42281_new_n2452_));
OR2X2 OR2X2_5932 ( .A(alu__abc_42281_new_n2444_), .B(alu__abc_42281_new_n2452_), .Y(alu__abc_42281_new_n2453_));
OR2X2 OR2X2_5933 ( .A(alu__abc_42281_new_n2457_), .B(alu__abc_42281_new_n2455_), .Y(alu__abc_42281_new_n2458_));
OR2X2 OR2X2_5934 ( .A(alu__abc_42281_new_n419_), .B(alu__abc_42281_new_n2459_), .Y(alu__abc_42281_new_n2460_));
OR2X2 OR2X2_5935 ( .A(alu__abc_42281_new_n2458_), .B(alu__abc_42281_new_n2462_), .Y(alu__abc_42281_new_n2463_));
OR2X2 OR2X2_5936 ( .A(alu__abc_42281_new_n2467_), .B(alu__abc_42281_new_n2465_), .Y(alu__abc_42281_new_n2468_));
OR2X2 OR2X2_5937 ( .A(alu__abc_42281_new_n434_), .B(alu__abc_42281_new_n2469_), .Y(alu__abc_42281_new_n2470_));
OR2X2 OR2X2_5938 ( .A(alu__abc_42281_new_n2468_), .B(alu__abc_42281_new_n2472_), .Y(alu__abc_42281_new_n2473_));
OR2X2 OR2X2_5939 ( .A(alu__abc_42281_new_n2464_), .B(alu__abc_42281_new_n2473_), .Y(alu__abc_42281_new_n2474_));
OR2X2 OR2X2_594 ( .A(_abc_44694_new_n2346_), .B(_abc_44694_new_n1278__bF_buf0), .Y(_abc_44694_new_n2347_));
OR2X2 OR2X2_5940 ( .A(alu__abc_42281_new_n2454_), .B(alu__abc_42281_new_n2474_), .Y(alu__abc_42281_new_n2475_));
OR2X2 OR2X2_5941 ( .A(alu__abc_42281_new_n2479_), .B(alu__abc_42281_new_n2477_), .Y(alu__abc_42281_new_n2480_));
OR2X2 OR2X2_5942 ( .A(alu__abc_42281_new_n485_), .B(alu__abc_42281_new_n2481_), .Y(alu__abc_42281_new_n2482_));
OR2X2 OR2X2_5943 ( .A(alu__abc_42281_new_n2480_), .B(alu__abc_42281_new_n2484_), .Y(alu__abc_42281_new_n2485_));
OR2X2 OR2X2_5944 ( .A(alu__abc_42281_new_n2489_), .B(alu__abc_42281_new_n2487_), .Y(alu__abc_42281_new_n2490_));
OR2X2 OR2X2_5945 ( .A(alu__abc_42281_new_n497_), .B(alu__abc_42281_new_n2491_), .Y(alu__abc_42281_new_n2492_));
OR2X2 OR2X2_5946 ( .A(alu__abc_42281_new_n2494_), .B(alu__abc_42281_new_n2490_), .Y(alu__abc_42281_new_n2495_));
OR2X2 OR2X2_5947 ( .A(alu__abc_42281_new_n2486_), .B(alu__abc_42281_new_n2495_), .Y(alu__abc_42281_new_n2496_));
OR2X2 OR2X2_5948 ( .A(alu__abc_42281_new_n2499_), .B(alu__abc_42281_new_n2497_), .Y(alu__abc_42281_new_n2500_));
OR2X2 OR2X2_5949 ( .A(alu__abc_42281_new_n451_), .B(alu__abc_42281_new_n2501_), .Y(alu__abc_42281_new_n2502_));
OR2X2 OR2X2_595 ( .A(_abc_44694_new_n2348_), .B(_abc_44694_new_n2349_), .Y(_abc_44694_new_n2350_));
OR2X2 OR2X2_5950 ( .A(alu__abc_42281_new_n2500_), .B(alu__abc_42281_new_n2504_), .Y(alu__abc_42281_new_n2505_));
OR2X2 OR2X2_5951 ( .A(alu__abc_42281_new_n2509_), .B(alu__abc_42281_new_n2507_), .Y(alu__abc_42281_new_n2510_));
OR2X2 OR2X2_5952 ( .A(alu__abc_42281_new_n466_), .B(alu__abc_42281_new_n2511_), .Y(alu__abc_42281_new_n2512_));
OR2X2 OR2X2_5953 ( .A(alu__abc_42281_new_n2510_), .B(alu__abc_42281_new_n2514_), .Y(alu__abc_42281_new_n2515_));
OR2X2 OR2X2_5954 ( .A(alu__abc_42281_new_n2506_), .B(alu__abc_42281_new_n2515_), .Y(alu__abc_42281_new_n2516_));
OR2X2 OR2X2_5955 ( .A(alu__abc_42281_new_n2517_), .B(alu__abc_42281_new_n2496_), .Y(alu__abc_42281_new_n2518_));
OR2X2 OR2X2_5956 ( .A(alu__abc_42281_new_n2476_), .B(alu__abc_42281_new_n2518_), .Y(alu__abc_42281_new_n2519_));
OR2X2 OR2X2_596 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n2350_), .Y(_abc_44694_new_n2351_));
OR2X2 OR2X2_597 ( .A(_abc_44694_new_n2353_), .B(_abc_44694_new_n2326_), .Y(_abc_44694_new_n2354_));
OR2X2 OR2X2_598 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(epc_q_26_), .Y(_abc_44694_new_n2355_));
OR2X2 OR2X2_599 ( .A(_abc_44694_new_n2322_), .B(pc_q_27_), .Y(_abc_44694_new_n2358_));
OR2X2 OR2X2_6 ( .A(_abc_44694_new_n665_), .B(state_q_3_bF_buf5_), .Y(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_2_));
OR2X2 OR2X2_60 ( .A(_abc_44694_new_n805_), .B(_abc_44694_new_n644_), .Y(_abc_44694_new_n806_));
OR2X2 OR2X2_600 ( .A(_abc_44694_new_n2362_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n2363_));
OR2X2 OR2X2_601 ( .A(opcode_q_25_), .B(pc_q_27_), .Y(_abc_44694_new_n2364_));
OR2X2 OR2X2_602 ( .A(_abc_44694_new_n2367_), .B(_abc_44694_new_n2331_), .Y(_abc_44694_new_n2368_));
OR2X2 OR2X2_603 ( .A(_abc_44694_new_n2335_), .B(_abc_44694_new_n2368_), .Y(_abc_44694_new_n2369_));
OR2X2 OR2X2_604 ( .A(_abc_44694_new_n2377_), .B(_abc_44694_new_n2378_), .Y(_abc_44694_new_n2379_));
OR2X2 OR2X2_605 ( .A(_abc_44694_new_n2380_), .B(_abc_44694_new_n2381_), .Y(_abc_44694_new_n2382_));
OR2X2 OR2X2_606 ( .A(_abc_44694_new_n2382_), .B(_abc_44694_new_n1400__bF_buf4), .Y(_abc_44694_new_n2383_));
OR2X2 OR2X2_607 ( .A(_abc_44694_new_n2361_), .B(_abc_44694_new_n1399__bF_buf3), .Y(_abc_44694_new_n2384_));
OR2X2 OR2X2_608 ( .A(_abc_44694_new_n2385_), .B(_abc_44694_new_n1278__bF_buf5), .Y(_abc_44694_new_n2386_));
OR2X2 OR2X2_609 ( .A(_abc_44694_new_n2387_), .B(_abc_44694_new_n2388_), .Y(_abc_44694_new_n2389_));
OR2X2 OR2X2_61 ( .A(_abc_44694_new_n807_), .B(_abc_44694_new_n671_), .Y(_abc_44694_new_n808_));
OR2X2 OR2X2_610 ( .A(_abc_44694_new_n1334__bF_buf2), .B(_abc_44694_new_n2389_), .Y(_abc_44694_new_n2390_));
OR2X2 OR2X2_611 ( .A(_abc_44694_new_n2392_), .B(_abc_44694_new_n2363_), .Y(_abc_44694_new_n2393_));
OR2X2 OR2X2_612 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(epc_q_27_), .Y(_abc_44694_new_n2394_));
OR2X2 OR2X2_613 ( .A(_abc_44694_new_n2359_), .B(pc_q_28_), .Y(_abc_44694_new_n2397_));
OR2X2 OR2X2_614 ( .A(_abc_44694_new_n2401_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n2402_));
OR2X2 OR2X2_615 ( .A(_abc_44694_new_n2371_), .B(_abc_44694_new_n2404_), .Y(_abc_44694_new_n2405_));
OR2X2 OR2X2_616 ( .A(opcode_q_25_), .B(pc_q_28_), .Y(_abc_44694_new_n2406_));
OR2X2 OR2X2_617 ( .A(_abc_44694_new_n2405_), .B(_abc_44694_new_n2409_), .Y(_abc_44694_new_n2410_));
OR2X2 OR2X2_618 ( .A(_abc_44694_new_n2414_), .B(_abc_44694_new_n2415_), .Y(_abc_44694_new_n2416_));
OR2X2 OR2X2_619 ( .A(_abc_44694_new_n2417_), .B(_abc_44694_new_n2418_), .Y(_abc_44694_new_n2419_));
OR2X2 OR2X2_62 ( .A(state_q_1_bF_buf4_), .B(alu_p_o_7_), .Y(_abc_44694_new_n809_));
OR2X2 OR2X2_620 ( .A(_abc_44694_new_n2419_), .B(_abc_44694_new_n1400__bF_buf3), .Y(_abc_44694_new_n2420_));
OR2X2 OR2X2_621 ( .A(_abc_44694_new_n2400_), .B(_abc_44694_new_n1399__bF_buf2), .Y(_abc_44694_new_n2421_));
OR2X2 OR2X2_622 ( .A(_abc_44694_new_n2422_), .B(_abc_44694_new_n1278__bF_buf4), .Y(_abc_44694_new_n2423_));
OR2X2 OR2X2_623 ( .A(_abc_44694_new_n2424_), .B(_abc_44694_new_n2425_), .Y(_abc_44694_new_n2426_));
OR2X2 OR2X2_624 ( .A(_abc_44694_new_n1334__bF_buf1), .B(_abc_44694_new_n2426_), .Y(_abc_44694_new_n2427_));
OR2X2 OR2X2_625 ( .A(_abc_44694_new_n2429_), .B(_abc_44694_new_n2402_), .Y(_abc_44694_new_n2430_));
OR2X2 OR2X2_626 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(epc_q_28_), .Y(_abc_44694_new_n2431_));
OR2X2 OR2X2_627 ( .A(_abc_44694_new_n2398_), .B(pc_q_29_), .Y(_abc_44694_new_n2434_));
OR2X2 OR2X2_628 ( .A(_abc_44694_new_n2438_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n2439_));
OR2X2 OR2X2_629 ( .A(opcode_q_25_), .B(pc_q_29_), .Y(_abc_44694_new_n2442_));
OR2X2 OR2X2_63 ( .A(state_q_1_bF_buf3_), .B(alu_p_o_8_), .Y(_abc_44694_new_n811_));
OR2X2 OR2X2_630 ( .A(_abc_44694_new_n2441_), .B(_abc_44694_new_n2445_), .Y(_abc_44694_new_n2446_));
OR2X2 OR2X2_631 ( .A(_abc_44694_new_n2440_), .B(_abc_44694_new_n2447_), .Y(_abc_44694_new_n2448_));
OR2X2 OR2X2_632 ( .A(_abc_44694_new_n1337__bF_buf3), .B(_abc_44694_new_n2451_), .Y(_abc_44694_new_n2452_));
OR2X2 OR2X2_633 ( .A(_abc_44694_new_n2450_), .B(_abc_44694_new_n2452_), .Y(_abc_44694_new_n2453_));
OR2X2 OR2X2_634 ( .A(_abc_44694_new_n1340__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_44694_new_n2454_));
OR2X2 OR2X2_635 ( .A(_abc_44694_new_n2455_), .B(_abc_44694_new_n1400__bF_buf2), .Y(_abc_44694_new_n2456_));
OR2X2 OR2X2_636 ( .A(_abc_44694_new_n2437_), .B(_abc_44694_new_n1399__bF_buf1), .Y(_abc_44694_new_n2457_));
OR2X2 OR2X2_637 ( .A(_abc_44694_new_n2458_), .B(_abc_44694_new_n1278__bF_buf3), .Y(_abc_44694_new_n2459_));
OR2X2 OR2X2_638 ( .A(_abc_44694_new_n2460_), .B(_abc_44694_new_n2461_), .Y(_abc_44694_new_n2462_));
OR2X2 OR2X2_639 ( .A(_abc_44694_new_n1334__bF_buf0), .B(_abc_44694_new_n2462_), .Y(_abc_44694_new_n2463_));
OR2X2 OR2X2_64 ( .A(_abc_44694_new_n676_), .B(\mem_dat_i[8] ), .Y(_abc_44694_new_n812_));
OR2X2 OR2X2_640 ( .A(_abc_44694_new_n2465_), .B(_abc_44694_new_n2439_), .Y(_abc_44694_new_n2466_));
OR2X2 OR2X2_641 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(epc_q_29_), .Y(_abc_44694_new_n2467_));
OR2X2 OR2X2_642 ( .A(_abc_44694_new_n2435_), .B(pc_q_30_), .Y(_abc_44694_new_n2470_));
OR2X2 OR2X2_643 ( .A(_abc_44694_new_n2474_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n2475_));
OR2X2 OR2X2_644 ( .A(_abc_44694_new_n2476_), .B(_abc_44694_new_n2478_), .Y(_abc_44694_new_n2479_));
OR2X2 OR2X2_645 ( .A(_abc_44694_new_n2480_), .B(_abc_44694_new_n2486_), .Y(_abc_44694_new_n2487_));
OR2X2 OR2X2_646 ( .A(_abc_44694_new_n2479_), .B(_abc_44694_new_n2488_), .Y(_abc_44694_new_n2489_));
OR2X2 OR2X2_647 ( .A(_abc_44694_new_n2491_), .B(_abc_44694_new_n2492_), .Y(_abc_44694_new_n2493_));
OR2X2 OR2X2_648 ( .A(_abc_44694_new_n2494_), .B(_abc_44694_new_n2495_), .Y(_abc_44694_new_n2496_));
OR2X2 OR2X2_649 ( .A(_abc_44694_new_n2496_), .B(_abc_44694_new_n1400__bF_buf1), .Y(_abc_44694_new_n2497_));
OR2X2 OR2X2_65 ( .A(_abc_44694_new_n677__bF_buf2), .B(_abc_44694_new_n688_), .Y(_abc_44694_new_n813_));
OR2X2 OR2X2_650 ( .A(_abc_44694_new_n2473_), .B(_abc_44694_new_n1399__bF_buf0), .Y(_abc_44694_new_n2498_));
OR2X2 OR2X2_651 ( .A(_abc_44694_new_n2499_), .B(_abc_44694_new_n1278__bF_buf2), .Y(_abc_44694_new_n2500_));
OR2X2 OR2X2_652 ( .A(_abc_44694_new_n2501_), .B(_abc_44694_new_n2502_), .Y(_abc_44694_new_n2503_));
OR2X2 OR2X2_653 ( .A(_abc_44694_new_n1334__bF_buf4), .B(_abc_44694_new_n2503_), .Y(_abc_44694_new_n2504_));
OR2X2 OR2X2_654 ( .A(_abc_44694_new_n2506_), .B(_abc_44694_new_n2475_), .Y(_abc_44694_new_n2507_));
OR2X2 OR2X2_655 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(epc_q_30_), .Y(_abc_44694_new_n2508_));
OR2X2 OR2X2_656 ( .A(_abc_44694_new_n2471_), .B(pc_q_31_), .Y(_abc_44694_new_n2511_));
OR2X2 OR2X2_657 ( .A(_abc_44694_new_n2515_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n2516_));
OR2X2 OR2X2_658 ( .A(_abc_44694_new_n2479_), .B(_abc_44694_new_n2482_), .Y(_abc_44694_new_n2520_));
OR2X2 OR2X2_659 ( .A(_abc_44694_new_n2522_), .B(_abc_44694_new_n2517_), .Y(_abc_44694_new_n2523_));
OR2X2 OR2X2_66 ( .A(_abc_44694_new_n816_), .B(_abc_44694_new_n671_), .Y(_abc_44694_new_n817_));
OR2X2 OR2X2_660 ( .A(_abc_44694_new_n2521_), .B(pc_q_31_), .Y(_abc_44694_new_n2524_));
OR2X2 OR2X2_661 ( .A(_abc_44694_new_n1337__bF_buf1), .B(_abc_44694_new_n2527_), .Y(_abc_44694_new_n2528_));
OR2X2 OR2X2_662 ( .A(_abc_44694_new_n2526_), .B(_abc_44694_new_n2528_), .Y(_abc_44694_new_n2529_));
OR2X2 OR2X2_663 ( .A(_abc_44694_new_n1340__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_44694_new_n2530_));
OR2X2 OR2X2_664 ( .A(_abc_44694_new_n2531_), .B(_abc_44694_new_n1400__bF_buf0), .Y(_abc_44694_new_n2532_));
OR2X2 OR2X2_665 ( .A(_abc_44694_new_n2514_), .B(_abc_44694_new_n1399__bF_buf4), .Y(_abc_44694_new_n2533_));
OR2X2 OR2X2_666 ( .A(_abc_44694_new_n2534_), .B(_abc_44694_new_n1278__bF_buf1), .Y(_abc_44694_new_n2535_));
OR2X2 OR2X2_667 ( .A(_abc_44694_new_n2536_), .B(_abc_44694_new_n2537_), .Y(_abc_44694_new_n2538_));
OR2X2 OR2X2_668 ( .A(_abc_44694_new_n1334__bF_buf3), .B(_abc_44694_new_n2538_), .Y(_abc_44694_new_n2539_));
OR2X2 OR2X2_669 ( .A(_abc_44694_new_n2541_), .B(_abc_44694_new_n2516_), .Y(_abc_44694_new_n2542_));
OR2X2 OR2X2_67 ( .A(_abc_44694_new_n815_), .B(_abc_44694_new_n817__bF_buf3), .Y(_abc_44694_new_n818_));
OR2X2 OR2X2_670 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(epc_q_31_), .Y(_abc_44694_new_n2543_));
OR2X2 OR2X2_671 ( .A(_abc_44694_new_n2547_), .B(_abc_44694_new_n1210__bF_buf1), .Y(_abc_44694_new_n2548_));
OR2X2 OR2X2_672 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(next_pc_r_0_), .Y(_abc_44694_new_n2549_));
OR2X2 OR2X2_673 ( .A(_abc_44694_new_n2552_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n2553_));
OR2X2 OR2X2_674 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(next_pc_r_1_), .Y(_abc_44694_new_n2554_));
OR2X2 OR2X2_675 ( .A(_abc_44694_new_n2557_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n2558_));
OR2X2 OR2X2_676 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(pc_q_2_), .Y(_abc_44694_new_n2559_));
OR2X2 OR2X2_677 ( .A(_abc_44694_new_n2562_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n2563_));
OR2X2 OR2X2_678 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(pc_q_3_), .Y(_abc_44694_new_n2564_));
OR2X2 OR2X2_679 ( .A(_abc_44694_new_n2567_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n2568_));
OR2X2 OR2X2_68 ( .A(_abc_44694_new_n820_), .B(_abc_44694_new_n821_), .Y(_abc_44694_new_n822_));
OR2X2 OR2X2_680 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(pc_q_4_), .Y(_abc_44694_new_n2569_));
OR2X2 OR2X2_681 ( .A(_abc_44694_new_n2572_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n2573_));
OR2X2 OR2X2_682 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(pc_q_5_), .Y(_abc_44694_new_n2574_));
OR2X2 OR2X2_683 ( .A(_abc_44694_new_n2577_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n2578_));
OR2X2 OR2X2_684 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(pc_q_6_), .Y(_abc_44694_new_n2579_));
OR2X2 OR2X2_685 ( .A(_abc_44694_new_n2582_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n2583_));
OR2X2 OR2X2_686 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(pc_q_7_), .Y(_abc_44694_new_n2584_));
OR2X2 OR2X2_687 ( .A(_abc_44694_new_n1639_), .B(_abc_44694_new_n1334__bF_buf2), .Y(_abc_44694_new_n2587_));
OR2X2 OR2X2_688 ( .A(_abc_44694_new_n2589_), .B(_abc_44694_new_n657_), .Y(_abc_44694_new_n2590_));
OR2X2 OR2X2_689 ( .A(_abc_44694_new_n2588_), .B(_abc_44694_new_n2590_), .Y(_0pc_q_31_0__8_));
OR2X2 OR2X2_69 ( .A(_abc_44694_new_n823_), .B(_abc_44694_new_n817__bF_buf2), .Y(_abc_44694_new_n824_));
OR2X2 OR2X2_690 ( .A(_abc_44694_new_n1681_), .B(_abc_44694_new_n1334__bF_buf1), .Y(_abc_44694_new_n2592_));
OR2X2 OR2X2_691 ( .A(_abc_44694_new_n1203_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n2595_));
OR2X2 OR2X2_692 ( .A(_abc_44694_new_n2594_), .B(_abc_44694_new_n2595_), .Y(_abc_44694_new_n2596_));
OR2X2 OR2X2_693 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(pc_q_9_), .Y(_abc_44694_new_n2597_));
OR2X2 OR2X2_694 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(pc_q_10_), .Y(_abc_44694_new_n2600_));
OR2X2 OR2X2_695 ( .A(_abc_44694_new_n2601_), .B(_abc_44694_new_n1044_), .Y(_abc_44694_new_n2602_));
OR2X2 OR2X2_696 ( .A(_abc_44694_new_n2602_), .B(_abc_44694_new_n1049_), .Y(_abc_44694_new_n2603_));
OR2X2 OR2X2_697 ( .A(_abc_44694_new_n2604_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n2605_));
OR2X2 OR2X2_698 ( .A(_abc_44694_new_n2609_), .B(_abc_44694_new_n1205_), .Y(_abc_44694_new_n2610_));
OR2X2 OR2X2_699 ( .A(_abc_44694_new_n2611_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n2612_));
OR2X2 OR2X2_7 ( .A(_abc_44694_new_n668__bF_buf4), .B(_abc_44694_new_n669_), .Y(_abc_28031_auto_fsm_map_cc_170_map_fsm_2380_1_));
OR2X2 OR2X2_70 ( .A(state_q_1_bF_buf2_), .B(alu_p_o_9_), .Y(_abc_44694_new_n825_));
OR2X2 OR2X2_700 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(pc_q_11_), .Y(_abc_44694_new_n2613_));
OR2X2 OR2X2_701 ( .A(_abc_44694_new_n2616_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n2617_));
OR2X2 OR2X2_702 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(pc_q_12_), .Y(_abc_44694_new_n2618_));
OR2X2 OR2X2_703 ( .A(_abc_44694_new_n2621_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n2622_));
OR2X2 OR2X2_704 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(pc_q_13_), .Y(_abc_44694_new_n2623_));
OR2X2 OR2X2_705 ( .A(_abc_44694_new_n2626_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n2627_));
OR2X2 OR2X2_706 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(pc_q_14_), .Y(_abc_44694_new_n2628_));
OR2X2 OR2X2_707 ( .A(_abc_44694_new_n2631_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n2632_));
OR2X2 OR2X2_708 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(pc_q_15_), .Y(_abc_44694_new_n2633_));
OR2X2 OR2X2_709 ( .A(_abc_44694_new_n2636_), .B(_abc_44694_new_n1210__bF_buf1), .Y(_abc_44694_new_n2637_));
OR2X2 OR2X2_71 ( .A(_abc_44694_new_n827_), .B(_abc_44694_new_n828_), .Y(_abc_44694_new_n829_));
OR2X2 OR2X2_710 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(pc_q_16_), .Y(_abc_44694_new_n2638_));
OR2X2 OR2X2_711 ( .A(_abc_44694_new_n2641_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n2642_));
OR2X2 OR2X2_712 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(pc_q_17_), .Y(_abc_44694_new_n2643_));
OR2X2 OR2X2_713 ( .A(_abc_44694_new_n2646_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n2647_));
OR2X2 OR2X2_714 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(pc_q_18_), .Y(_abc_44694_new_n2648_));
OR2X2 OR2X2_715 ( .A(_abc_44694_new_n2651_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n2652_));
OR2X2 OR2X2_716 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(pc_q_19_), .Y(_abc_44694_new_n2653_));
OR2X2 OR2X2_717 ( .A(_abc_44694_new_n2656_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n2657_));
OR2X2 OR2X2_718 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(pc_q_20_), .Y(_abc_44694_new_n2658_));
OR2X2 OR2X2_719 ( .A(_abc_44694_new_n2661_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n2662_));
OR2X2 OR2X2_72 ( .A(_abc_44694_new_n830_), .B(_abc_44694_new_n817__bF_buf1), .Y(_abc_44694_new_n831_));
OR2X2 OR2X2_720 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(pc_q_21_), .Y(_abc_44694_new_n2663_));
OR2X2 OR2X2_721 ( .A(_abc_44694_new_n2666_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n2667_));
OR2X2 OR2X2_722 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(pc_q_22_), .Y(_abc_44694_new_n2668_));
OR2X2 OR2X2_723 ( .A(_abc_44694_new_n2671_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n2672_));
OR2X2 OR2X2_724 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(pc_q_23_), .Y(_abc_44694_new_n2673_));
OR2X2 OR2X2_725 ( .A(_abc_44694_new_n2676_), .B(_abc_44694_new_n1210__bF_buf1), .Y(_abc_44694_new_n2677_));
OR2X2 OR2X2_726 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf1), .B(pc_q_24_), .Y(_abc_44694_new_n2678_));
OR2X2 OR2X2_727 ( .A(_abc_44694_new_n2681_), .B(_abc_44694_new_n1210__bF_buf0), .Y(_abc_44694_new_n2682_));
OR2X2 OR2X2_728 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf0), .B(pc_q_25_), .Y(_abc_44694_new_n2683_));
OR2X2 OR2X2_729 ( .A(_abc_44694_new_n2686_), .B(_abc_44694_new_n1210__bF_buf7), .Y(_abc_44694_new_n2687_));
OR2X2 OR2X2_73 ( .A(state_q_1_bF_buf1_), .B(alu_p_o_10_), .Y(_abc_44694_new_n832_));
OR2X2 OR2X2_730 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf7), .B(pc_q_26_), .Y(_abc_44694_new_n2688_));
OR2X2 OR2X2_731 ( .A(_abc_44694_new_n2691_), .B(_abc_44694_new_n1210__bF_buf6), .Y(_abc_44694_new_n2692_));
OR2X2 OR2X2_732 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf6), .B(pc_q_27_), .Y(_abc_44694_new_n2693_));
OR2X2 OR2X2_733 ( .A(_abc_44694_new_n2696_), .B(_abc_44694_new_n1210__bF_buf5), .Y(_abc_44694_new_n2697_));
OR2X2 OR2X2_734 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf5), .B(pc_q_28_), .Y(_abc_44694_new_n2698_));
OR2X2 OR2X2_735 ( .A(_abc_44694_new_n2701_), .B(_abc_44694_new_n1210__bF_buf4), .Y(_abc_44694_new_n2702_));
OR2X2 OR2X2_736 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf4), .B(pc_q_29_), .Y(_abc_44694_new_n2703_));
OR2X2 OR2X2_737 ( .A(_abc_44694_new_n2706_), .B(_abc_44694_new_n1210__bF_buf3), .Y(_abc_44694_new_n2707_));
OR2X2 OR2X2_738 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf3), .B(pc_q_30_), .Y(_abc_44694_new_n2708_));
OR2X2 OR2X2_739 ( .A(_abc_44694_new_n2711_), .B(_abc_44694_new_n1210__bF_buf2), .Y(_abc_44694_new_n2712_));
OR2X2 OR2X2_74 ( .A(_abc_44694_new_n834_), .B(_abc_44694_new_n835_), .Y(_abc_44694_new_n836_));
OR2X2 OR2X2_740 ( .A(REGFILE_SIM_reg_bank_wr_i_bF_buf2), .B(pc_q_31_), .Y(_abc_44694_new_n2713_));
OR2X2 OR2X2_741 ( .A(_abc_44694_new_n2717_), .B(_abc_44694_new_n2718_), .Y(_abc_44694_new_n2719_));
OR2X2 OR2X2_742 ( .A(_abc_44694_new_n653_), .B(_abc_44694_new_n2723_), .Y(_abc_44694_new_n2724_));
OR2X2 OR2X2_743 ( .A(_abc_44694_new_n2716_), .B(_abc_44694_new_n2724_), .Y(_abc_44694_new_n2725_));
OR2X2 OR2X2_744 ( .A(_abc_44694_new_n2725_), .B(_abc_44694_new_n1162_), .Y(_abc_44694_new_n2726_));
OR2X2 OR2X2_745 ( .A(_abc_44694_new_n1080_), .B(_abc_44694_new_n1104_), .Y(_abc_44694_new_n2727_));
OR2X2 OR2X2_746 ( .A(_abc_44694_new_n1011_), .B(_abc_44694_new_n1037_), .Y(_abc_44694_new_n2728_));
OR2X2 OR2X2_747 ( .A(_abc_44694_new_n2728_), .B(_abc_44694_new_n1347__bF_buf3), .Y(_abc_44694_new_n2729_));
OR2X2 OR2X2_748 ( .A(_abc_44694_new_n2730_), .B(_abc_44694_new_n2727_), .Y(_abc_44694_new_n2731_));
OR2X2 OR2X2_749 ( .A(_abc_44694_new_n2731_), .B(_abc_44694_new_n2726_), .Y(_abc_44694_new_n2732_));
OR2X2 OR2X2_75 ( .A(_abc_44694_new_n837_), .B(_abc_44694_new_n817__bF_buf0), .Y(_abc_44694_new_n838_));
OR2X2 OR2X2_750 ( .A(_abc_44694_new_n2733_), .B(_abc_44694_new_n1178__bF_buf3), .Y(_0ex_rd_q_4_0__0_));
OR2X2 OR2X2_751 ( .A(_abc_44694_new_n2739_), .B(_abc_44694_new_n1178__bF_buf2), .Y(_0ex_rd_q_4_0__3_));
OR2X2 OR2X2_752 ( .A(_abc_44694_new_n2745_), .B(_abc_44694_new_n1187_), .Y(_abc_44694_new_n2746_));
OR2X2 OR2X2_753 ( .A(_abc_44694_new_n1144_), .B(_abc_44694_new_n2748_), .Y(_abc_44694_new_n2749_));
OR2X2 OR2X2_754 ( .A(_abc_44694_new_n2746_), .B(_abc_44694_new_n2749_), .Y(_abc_44694_new_n2750_));
OR2X2 OR2X2_755 ( .A(_abc_44694_new_n2750_), .B(_abc_44694_new_n2744_), .Y(_abc_44694_new_n2751_));
OR2X2 OR2X2_756 ( .A(_abc_44694_new_n2751_), .B(_abc_44694_new_n1146_), .Y(_abc_44694_new_n2752_));
OR2X2 OR2X2_757 ( .A(_abc_44694_new_n2727_), .B(_abc_44694_new_n1161_), .Y(_abc_44694_new_n2754_));
OR2X2 OR2X2_758 ( .A(_abc_44694_new_n2754_), .B(_abc_44694_new_n1086_), .Y(_abc_44694_new_n2755_));
OR2X2 OR2X2_759 ( .A(_abc_44694_new_n2756_), .B(_abc_44694_new_n2753_), .Y(alu_input_b_r_0_));
OR2X2 OR2X2_76 ( .A(state_q_1_bF_buf0_), .B(alu_p_o_11_), .Y(_abc_44694_new_n839_));
OR2X2 OR2X2_760 ( .A(_abc_44694_new_n2759_), .B(_abc_44694_new_n2758_), .Y(alu_input_b_r_1_));
OR2X2 OR2X2_761 ( .A(_abc_44694_new_n2762_), .B(_abc_44694_new_n2761_), .Y(alu_input_b_r_2_));
OR2X2 OR2X2_762 ( .A(_abc_44694_new_n2765_), .B(_abc_44694_new_n2764_), .Y(alu_input_b_r_3_));
OR2X2 OR2X2_763 ( .A(_abc_44694_new_n2768_), .B(_abc_44694_new_n2767_), .Y(alu_input_b_r_4_));
OR2X2 OR2X2_764 ( .A(_abc_44694_new_n2771_), .B(_abc_44694_new_n2770_), .Y(alu_input_b_r_5_));
OR2X2 OR2X2_765 ( .A(_abc_44694_new_n2774_), .B(_abc_44694_new_n1146_), .Y(_abc_44694_new_n2775_));
OR2X2 OR2X2_766 ( .A(_abc_44694_new_n2776_), .B(_abc_44694_new_n2777_), .Y(_abc_44694_new_n2778_));
OR2X2 OR2X2_767 ( .A(_abc_44694_new_n1080_), .B(_abc_44694_new_n1160_), .Y(_abc_44694_new_n2779_));
OR2X2 OR2X2_768 ( .A(_abc_44694_new_n2778_), .B(_abc_44694_new_n2780_), .Y(alu_input_b_r_6_));
OR2X2 OR2X2_769 ( .A(_abc_44694_new_n2782_), .B(_abc_44694_new_n2783_), .Y(_abc_44694_new_n2784_));
OR2X2 OR2X2_77 ( .A(state_q_1_bF_buf4_), .B(alu_p_o_12_), .Y(_abc_44694_new_n841_));
OR2X2 OR2X2_770 ( .A(_abc_44694_new_n2784_), .B(_abc_44694_new_n2785_), .Y(alu_input_b_r_7_));
OR2X2 OR2X2_771 ( .A(_abc_44694_new_n2787_), .B(_abc_44694_new_n2788_), .Y(_abc_44694_new_n2789_));
OR2X2 OR2X2_772 ( .A(_abc_44694_new_n2789_), .B(_abc_44694_new_n2790_), .Y(alu_input_b_r_8_));
OR2X2 OR2X2_773 ( .A(_abc_44694_new_n2792_), .B(_abc_44694_new_n2793_), .Y(_abc_44694_new_n2794_));
OR2X2 OR2X2_774 ( .A(_abc_44694_new_n2794_), .B(_abc_44694_new_n2795_), .Y(alu_input_b_r_9_));
OR2X2 OR2X2_775 ( .A(_abc_44694_new_n2797_), .B(_abc_44694_new_n2798_), .Y(_abc_44694_new_n2799_));
OR2X2 OR2X2_776 ( .A(_abc_44694_new_n2799_), .B(_abc_44694_new_n2800_), .Y(alu_input_b_r_10_));
OR2X2 OR2X2_777 ( .A(_abc_44694_new_n2802_), .B(_abc_44694_new_n2803_), .Y(_abc_44694_new_n2804_));
OR2X2 OR2X2_778 ( .A(_abc_44694_new_n2804_), .B(_abc_44694_new_n2805_), .Y(alu_input_b_r_11_));
OR2X2 OR2X2_779 ( .A(_abc_44694_new_n2807_), .B(_abc_44694_new_n2808_), .Y(_abc_44694_new_n2809_));
OR2X2 OR2X2_78 ( .A(_abc_44694_new_n676_), .B(\mem_dat_i[12] ), .Y(_abc_44694_new_n842_));
OR2X2 OR2X2_780 ( .A(_abc_44694_new_n2809_), .B(_abc_44694_new_n2810_), .Y(alu_input_b_r_12_));
OR2X2 OR2X2_781 ( .A(_abc_44694_new_n2812_), .B(_abc_44694_new_n2813_), .Y(_abc_44694_new_n2814_));
OR2X2 OR2X2_782 ( .A(_abc_44694_new_n2814_), .B(_abc_44694_new_n2815_), .Y(alu_input_b_r_13_));
OR2X2 OR2X2_783 ( .A(_abc_44694_new_n2817_), .B(_abc_44694_new_n2818_), .Y(_abc_44694_new_n2819_));
OR2X2 OR2X2_784 ( .A(_abc_44694_new_n2819_), .B(_abc_44694_new_n2820_), .Y(alu_input_b_r_14_));
OR2X2 OR2X2_785 ( .A(_abc_44694_new_n1087__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_15_), .Y(_abc_44694_new_n2822_));
OR2X2 OR2X2_786 ( .A(_abc_44694_new_n2773_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf3_), .Y(_abc_44694_new_n2824_));
OR2X2 OR2X2_787 ( .A(_abc_44694_new_n2825_), .B(_abc_44694_new_n1086_), .Y(_abc_44694_new_n2826_));
OR2X2 OR2X2_788 ( .A(_abc_44694_new_n2774_), .B(_abc_44694_new_n2826__bF_buf3), .Y(_abc_44694_new_n2827_));
OR2X2 OR2X2_789 ( .A(_abc_44694_new_n2823_), .B(_abc_44694_new_n2828_), .Y(_abc_44694_new_n2829_));
OR2X2 OR2X2_79 ( .A(_abc_44694_new_n677__bF_buf1), .B(_abc_44694_new_n754_), .Y(_abc_44694_new_n843_));
OR2X2 OR2X2_790 ( .A(_abc_44694_new_n2831_), .B(REGFILE_SIM_reg_bank_rb_i_4_bF_buf1_), .Y(_abc_44694_new_n2832_));
OR2X2 OR2X2_791 ( .A(_abc_44694_new_n1087__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_16_), .Y(_abc_44694_new_n2836_));
OR2X2 OR2X2_792 ( .A(_abc_44694_new_n2837_), .B(_abc_44694_new_n1084__bF_buf1), .Y(_abc_44694_new_n2838_));
OR2X2 OR2X2_793 ( .A(_abc_44694_new_n2839_), .B(_abc_44694_new_n1181__bF_buf1), .Y(_abc_44694_new_n2840_));
OR2X2 OR2X2_794 ( .A(_abc_44694_new_n2841_), .B(_abc_44694_new_n2842_), .Y(alu_input_b_r_16_));
OR2X2 OR2X2_795 ( .A(_abc_44694_new_n1087__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_17_), .Y(_abc_44694_new_n2844_));
OR2X2 OR2X2_796 ( .A(_abc_44694_new_n2845_), .B(_abc_44694_new_n1084__bF_buf0), .Y(_abc_44694_new_n2846_));
OR2X2 OR2X2_797 ( .A(_abc_44694_new_n2847_), .B(_abc_44694_new_n1181__bF_buf0), .Y(_abc_44694_new_n2848_));
OR2X2 OR2X2_798 ( .A(_abc_44694_new_n2849_), .B(_abc_44694_new_n2850_), .Y(alu_input_b_r_17_));
OR2X2 OR2X2_799 ( .A(_abc_44694_new_n1087__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_18_), .Y(_abc_44694_new_n2852_));
OR2X2 OR2X2_8 ( .A(_abc_44694_new_n677__bF_buf3), .B(_abc_44694_new_n675_), .Y(_abc_44694_new_n678_));
OR2X2 OR2X2_80 ( .A(_abc_44694_new_n845_), .B(_abc_44694_new_n817__bF_buf3), .Y(_abc_44694_new_n846_));
OR2X2 OR2X2_800 ( .A(_abc_44694_new_n2853_), .B(_abc_44694_new_n1084__bF_buf3), .Y(_abc_44694_new_n2854_));
OR2X2 OR2X2_801 ( .A(_abc_44694_new_n2855_), .B(_abc_44694_new_n1181__bF_buf3), .Y(_abc_44694_new_n2856_));
OR2X2 OR2X2_802 ( .A(_abc_44694_new_n2857_), .B(_abc_44694_new_n2858_), .Y(alu_input_b_r_18_));
OR2X2 OR2X2_803 ( .A(_abc_44694_new_n1087__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_19_), .Y(_abc_44694_new_n2860_));
OR2X2 OR2X2_804 ( .A(_abc_44694_new_n2861_), .B(_abc_44694_new_n1084__bF_buf2), .Y(_abc_44694_new_n2862_));
OR2X2 OR2X2_805 ( .A(_abc_44694_new_n2863_), .B(_abc_44694_new_n1181__bF_buf2), .Y(_abc_44694_new_n2864_));
OR2X2 OR2X2_806 ( .A(_abc_44694_new_n2865_), .B(_abc_44694_new_n2866_), .Y(alu_input_b_r_19_));
OR2X2 OR2X2_807 ( .A(_abc_44694_new_n1087__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_20_), .Y(_abc_44694_new_n2868_));
OR2X2 OR2X2_808 ( .A(_abc_44694_new_n2869_), .B(_abc_44694_new_n1084__bF_buf1), .Y(_abc_44694_new_n2870_));
OR2X2 OR2X2_809 ( .A(_abc_44694_new_n2871_), .B(_abc_44694_new_n1181__bF_buf1), .Y(_abc_44694_new_n2872_));
OR2X2 OR2X2_81 ( .A(state_q_1_bF_buf3_), .B(alu_p_o_13_), .Y(_abc_44694_new_n848_));
OR2X2 OR2X2_810 ( .A(_abc_44694_new_n2873_), .B(_abc_44694_new_n2874_), .Y(alu_input_b_r_20_));
OR2X2 OR2X2_811 ( .A(_abc_44694_new_n1087__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_21_), .Y(_abc_44694_new_n2876_));
OR2X2 OR2X2_812 ( .A(_abc_44694_new_n2877_), .B(_abc_44694_new_n1084__bF_buf0), .Y(_abc_44694_new_n2878_));
OR2X2 OR2X2_813 ( .A(_abc_44694_new_n2879_), .B(_abc_44694_new_n1181__bF_buf0), .Y(_abc_44694_new_n2880_));
OR2X2 OR2X2_814 ( .A(_abc_44694_new_n2881_), .B(_abc_44694_new_n2882_), .Y(alu_input_b_r_21_));
OR2X2 OR2X2_815 ( .A(_abc_44694_new_n1087__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_22_), .Y(_abc_44694_new_n2884_));
OR2X2 OR2X2_816 ( .A(_abc_44694_new_n2885_), .B(_abc_44694_new_n1084__bF_buf3), .Y(_abc_44694_new_n2886_));
OR2X2 OR2X2_817 ( .A(_abc_44694_new_n2887_), .B(_abc_44694_new_n1181__bF_buf3), .Y(_abc_44694_new_n2888_));
OR2X2 OR2X2_818 ( .A(_abc_44694_new_n2889_), .B(_abc_44694_new_n2890_), .Y(alu_input_b_r_22_));
OR2X2 OR2X2_819 ( .A(_abc_44694_new_n1087__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_23_), .Y(_abc_44694_new_n2892_));
OR2X2 OR2X2_82 ( .A(_abc_44694_new_n676_), .B(\mem_dat_i[13] ), .Y(_abc_44694_new_n849_));
OR2X2 OR2X2_820 ( .A(_abc_44694_new_n2893_), .B(_abc_44694_new_n1084__bF_buf2), .Y(_abc_44694_new_n2894_));
OR2X2 OR2X2_821 ( .A(_abc_44694_new_n2895_), .B(_abc_44694_new_n1181__bF_buf2), .Y(_abc_44694_new_n2896_));
OR2X2 OR2X2_822 ( .A(_abc_44694_new_n2897_), .B(_abc_44694_new_n2898_), .Y(alu_input_b_r_23_));
OR2X2 OR2X2_823 ( .A(_abc_44694_new_n1087__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_24_), .Y(_abc_44694_new_n2900_));
OR2X2 OR2X2_824 ( .A(_abc_44694_new_n2901_), .B(_abc_44694_new_n1084__bF_buf1), .Y(_abc_44694_new_n2902_));
OR2X2 OR2X2_825 ( .A(_abc_44694_new_n2903_), .B(_abc_44694_new_n1181__bF_buf1), .Y(_abc_44694_new_n2904_));
OR2X2 OR2X2_826 ( .A(_abc_44694_new_n2905_), .B(_abc_44694_new_n2906_), .Y(alu_input_b_r_24_));
OR2X2 OR2X2_827 ( .A(_abc_44694_new_n1087__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_25_), .Y(_abc_44694_new_n2908_));
OR2X2 OR2X2_828 ( .A(_abc_44694_new_n2909_), .B(_abc_44694_new_n1084__bF_buf0), .Y(_abc_44694_new_n2910_));
OR2X2 OR2X2_829 ( .A(_abc_44694_new_n2911_), .B(_abc_44694_new_n1181__bF_buf0), .Y(_abc_44694_new_n2912_));
OR2X2 OR2X2_83 ( .A(_abc_44694_new_n677__bF_buf0), .B(_abc_44694_new_n770_), .Y(_abc_44694_new_n850_));
OR2X2 OR2X2_830 ( .A(_abc_44694_new_n2913_), .B(_abc_44694_new_n2914_), .Y(alu_input_b_r_25_));
OR2X2 OR2X2_831 ( .A(_abc_44694_new_n1087__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_26_), .Y(_abc_44694_new_n2916_));
OR2X2 OR2X2_832 ( .A(_abc_44694_new_n2917_), .B(_abc_44694_new_n1084__bF_buf3), .Y(_abc_44694_new_n2918_));
OR2X2 OR2X2_833 ( .A(_abc_44694_new_n2919_), .B(_abc_44694_new_n1181__bF_buf3), .Y(_abc_44694_new_n2920_));
OR2X2 OR2X2_834 ( .A(_abc_44694_new_n2921_), .B(_abc_44694_new_n2922_), .Y(alu_input_b_r_26_));
OR2X2 OR2X2_835 ( .A(_abc_44694_new_n1087__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_27_), .Y(_abc_44694_new_n2924_));
OR2X2 OR2X2_836 ( .A(_abc_44694_new_n2925_), .B(_abc_44694_new_n1084__bF_buf2), .Y(_abc_44694_new_n2926_));
OR2X2 OR2X2_837 ( .A(_abc_44694_new_n2927_), .B(_abc_44694_new_n1181__bF_buf2), .Y(_abc_44694_new_n2928_));
OR2X2 OR2X2_838 ( .A(_abc_44694_new_n2929_), .B(_abc_44694_new_n2930_), .Y(alu_input_b_r_27_));
OR2X2 OR2X2_839 ( .A(_abc_44694_new_n1087__bF_buf1), .B(REGFILE_SIM_reg_bank_reg_rb_o_28_), .Y(_abc_44694_new_n2932_));
OR2X2 OR2X2_84 ( .A(_abc_44694_new_n852_), .B(_abc_44694_new_n817__bF_buf2), .Y(_abc_44694_new_n853_));
OR2X2 OR2X2_840 ( .A(_abc_44694_new_n2933_), .B(_abc_44694_new_n1084__bF_buf1), .Y(_abc_44694_new_n2934_));
OR2X2 OR2X2_841 ( .A(_abc_44694_new_n2935_), .B(_abc_44694_new_n1181__bF_buf1), .Y(_abc_44694_new_n2936_));
OR2X2 OR2X2_842 ( .A(_abc_44694_new_n2937_), .B(_abc_44694_new_n2938_), .Y(alu_input_b_r_28_));
OR2X2 OR2X2_843 ( .A(_abc_44694_new_n1087__bF_buf0), .B(REGFILE_SIM_reg_bank_reg_rb_o_29_), .Y(_abc_44694_new_n2940_));
OR2X2 OR2X2_844 ( .A(_abc_44694_new_n2941_), .B(_abc_44694_new_n1084__bF_buf0), .Y(_abc_44694_new_n2942_));
OR2X2 OR2X2_845 ( .A(_abc_44694_new_n2943_), .B(_abc_44694_new_n1181__bF_buf0), .Y(_abc_44694_new_n2944_));
OR2X2 OR2X2_846 ( .A(_abc_44694_new_n2945_), .B(_abc_44694_new_n2946_), .Y(alu_input_b_r_29_));
OR2X2 OR2X2_847 ( .A(_abc_44694_new_n1087__bF_buf3), .B(REGFILE_SIM_reg_bank_reg_rb_o_30_), .Y(_abc_44694_new_n2948_));
OR2X2 OR2X2_848 ( .A(_abc_44694_new_n2949_), .B(_abc_44694_new_n1084__bF_buf3), .Y(_abc_44694_new_n2950_));
OR2X2 OR2X2_849 ( .A(_abc_44694_new_n2951_), .B(_abc_44694_new_n1181__bF_buf3), .Y(_abc_44694_new_n2952_));
OR2X2 OR2X2_85 ( .A(_abc_44694_new_n855_), .B(_abc_44694_new_n856_), .Y(_abc_44694_new_n857_));
OR2X2 OR2X2_850 ( .A(_abc_44694_new_n2953_), .B(_abc_44694_new_n2954_), .Y(alu_input_b_r_30_));
OR2X2 OR2X2_851 ( .A(_abc_44694_new_n1087__bF_buf2), .B(REGFILE_SIM_reg_bank_reg_rb_o_31_), .Y(_abc_44694_new_n2956_));
OR2X2 OR2X2_852 ( .A(_abc_44694_new_n2957_), .B(_abc_44694_new_n1084__bF_buf2), .Y(_abc_44694_new_n2958_));
OR2X2 OR2X2_853 ( .A(_abc_44694_new_n2959_), .B(_abc_44694_new_n1181__bF_buf2), .Y(_abc_44694_new_n2960_));
OR2X2 OR2X2_854 ( .A(_abc_44694_new_n2961_), .B(_abc_44694_new_n2962_), .Y(alu_input_b_r_31_));
OR2X2 OR2X2_855 ( .A(_abc_44694_new_n1089_), .B(_abc_44694_new_n1146_), .Y(_abc_44694_new_n2964_));
OR2X2 OR2X2_856 ( .A(_abc_44694_new_n2750_), .B(_abc_44694_new_n2964_), .Y(_abc_44694_new_n2965_));
OR2X2 OR2X2_857 ( .A(_abc_44694_new_n2966_), .B(_abc_44694_new_n2968_), .Y(_abc_44694_new_n2969_));
OR2X2 OR2X2_858 ( .A(_abc_44694_new_n2969_), .B(_abc_44694_new_n2970_), .Y(_abc_44694_new_n2971_));
OR2X2 OR2X2_859 ( .A(_abc_44694_new_n2754_), .B(_abc_44694_new_n1183_), .Y(_abc_44694_new_n2972_));
OR2X2 OR2X2_86 ( .A(_abc_44694_new_n858_), .B(_abc_44694_new_n817__bF_buf1), .Y(_abc_44694_new_n859_));
OR2X2 OR2X2_860 ( .A(_abc_44694_new_n2973_), .B(_abc_44694_new_n2971_), .Y(alu_input_a_r_0_));
OR2X2 OR2X2_861 ( .A(_abc_44694_new_n2975_), .B(_abc_44694_new_n2977_), .Y(_abc_44694_new_n2978_));
OR2X2 OR2X2_862 ( .A(_abc_44694_new_n2978_), .B(_abc_44694_new_n2979_), .Y(_abc_44694_new_n2980_));
OR2X2 OR2X2_863 ( .A(_abc_44694_new_n2981_), .B(_abc_44694_new_n2980_), .Y(alu_input_a_r_1_));
OR2X2 OR2X2_864 ( .A(_abc_44694_new_n2984_), .B(_abc_44694_new_n2985_), .Y(_abc_44694_new_n2986_));
OR2X2 OR2X2_865 ( .A(_abc_44694_new_n2983_), .B(_abc_44694_new_n2986_), .Y(_abc_44694_new_n2987_));
OR2X2 OR2X2_866 ( .A(_abc_44694_new_n2989_), .B(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n2990_));
OR2X2 OR2X2_867 ( .A(_abc_44694_new_n2988_), .B(_abc_44694_new_n2990_), .Y(_abc_44694_new_n2991_));
OR2X2 OR2X2_868 ( .A(_abc_44694_new_n1179__bF_buf3), .B(_abc_44694_new_n1412_), .Y(_abc_44694_new_n2992_));
OR2X2 OR2X2_869 ( .A(_abc_44694_new_n2993_), .B(_abc_44694_new_n2994_), .Y(alu_input_a_r_2_));
OR2X2 OR2X2_87 ( .A(state_q_1_bF_buf2_), .B(alu_p_o_14_), .Y(_abc_44694_new_n860_));
OR2X2 OR2X2_870 ( .A(_abc_44694_new_n2996_), .B(_abc_44694_new_n2998_), .Y(_abc_44694_new_n2999_));
OR2X2 OR2X2_871 ( .A(_abc_44694_new_n2999_), .B(_abc_44694_new_n3000_), .Y(_abc_44694_new_n3001_));
OR2X2 OR2X2_872 ( .A(_abc_44694_new_n3002_), .B(_abc_44694_new_n3001_), .Y(alu_input_a_r_3_));
OR2X2 OR2X2_873 ( .A(_abc_44694_new_n3005_), .B(_abc_44694_new_n3007_), .Y(_abc_44694_new_n3008_));
OR2X2 OR2X2_874 ( .A(_abc_44694_new_n3008_), .B(_abc_44694_new_n3009_), .Y(_abc_44694_new_n3010_));
OR2X2 OR2X2_875 ( .A(_abc_44694_new_n3011_), .B(_abc_44694_new_n3010_), .Y(alu_input_a_r_4_));
OR2X2 OR2X2_876 ( .A(_abc_44694_new_n3013_), .B(_abc_44694_new_n3015_), .Y(_abc_44694_new_n3016_));
OR2X2 OR2X2_877 ( .A(_abc_44694_new_n3016_), .B(_abc_44694_new_n3017_), .Y(_abc_44694_new_n3018_));
OR2X2 OR2X2_878 ( .A(_abc_44694_new_n3019_), .B(_abc_44694_new_n3018_), .Y(alu_input_a_r_5_));
OR2X2 OR2X2_879 ( .A(_abc_44694_new_n3022_), .B(_abc_44694_new_n3024_), .Y(_abc_44694_new_n3025_));
OR2X2 OR2X2_88 ( .A(state_q_1_bF_buf1_), .B(alu_p_o_15_), .Y(_abc_44694_new_n862_));
OR2X2 OR2X2_880 ( .A(_abc_44694_new_n3025_), .B(_abc_44694_new_n3026_), .Y(_abc_44694_new_n3027_));
OR2X2 OR2X2_881 ( .A(_abc_44694_new_n3028_), .B(_abc_44694_new_n3027_), .Y(alu_input_a_r_6_));
OR2X2 OR2X2_882 ( .A(_abc_44694_new_n3030_), .B(_abc_44694_new_n3032_), .Y(_abc_44694_new_n3033_));
OR2X2 OR2X2_883 ( .A(_abc_44694_new_n3033_), .B(_abc_44694_new_n3034_), .Y(_abc_44694_new_n3035_));
OR2X2 OR2X2_884 ( .A(_abc_44694_new_n3036_), .B(_abc_44694_new_n3035_), .Y(alu_input_a_r_7_));
OR2X2 OR2X2_885 ( .A(_abc_44694_new_n3039_), .B(_abc_44694_new_n3041_), .Y(_abc_44694_new_n3042_));
OR2X2 OR2X2_886 ( .A(_abc_44694_new_n3042_), .B(_abc_44694_new_n3043_), .Y(_abc_44694_new_n3044_));
OR2X2 OR2X2_887 ( .A(_abc_44694_new_n3045_), .B(_abc_44694_new_n3044_), .Y(alu_input_a_r_8_));
OR2X2 OR2X2_888 ( .A(_abc_44694_new_n3048_), .B(_abc_44694_new_n1115_), .Y(_abc_44694_new_n3049_));
OR2X2 OR2X2_889 ( .A(_abc_44694_new_n3049_), .B(_abc_44694_new_n3047_), .Y(_abc_44694_new_n3050_));
OR2X2 OR2X2_89 ( .A(_abc_44694_new_n676_), .B(\mem_dat_i[15] ), .Y(_abc_44694_new_n863_));
OR2X2 OR2X2_890 ( .A(_abc_44694_new_n3051_), .B(_abc_44694_new_n3050_), .Y(_abc_44694_new_n3052_));
OR2X2 OR2X2_891 ( .A(_abc_44694_new_n3053_), .B(_abc_44694_new_n1114__bF_buf3), .Y(_abc_44694_new_n3054_));
OR2X2 OR2X2_892 ( .A(_abc_44694_new_n3055_), .B(_abc_44694_new_n3056_), .Y(_abc_44694_new_n3057_));
OR2X2 OR2X2_893 ( .A(_abc_44694_new_n3057_), .B(_abc_44694_new_n3058_), .Y(alu_input_a_r_9_));
OR2X2 OR2X2_894 ( .A(_abc_44694_new_n3061_), .B(_abc_44694_new_n3062_), .Y(_abc_44694_new_n3063_));
OR2X2 OR2X2_895 ( .A(_abc_44694_new_n3064_), .B(_abc_44694_new_n3063_), .Y(_abc_44694_new_n3065_));
OR2X2 OR2X2_896 ( .A(_abc_44694_new_n3066_), .B(_abc_44694_new_n3060_), .Y(_abc_44694_new_n3067_));
OR2X2 OR2X2_897 ( .A(_abc_44694_new_n3067_), .B(_abc_44694_new_n3068_), .Y(_abc_44694_new_n3069_));
OR2X2 OR2X2_898 ( .A(_abc_44694_new_n3069_), .B(_abc_44694_new_n3070_), .Y(alu_input_a_r_10_));
OR2X2 OR2X2_899 ( .A(_abc_44694_new_n3072_), .B(_abc_44694_new_n1115_), .Y(_abc_44694_new_n3073_));
OR2X2 OR2X2_9 ( .A(_abc_44694_new_n679_), .B(_abc_44694_new_n683_), .Y(_abc_44694_new_n684_));
OR2X2 OR2X2_90 ( .A(_abc_44694_new_n677__bF_buf3), .B(_abc_44694_new_n797_), .Y(_abc_44694_new_n864_));
OR2X2 OR2X2_900 ( .A(_abc_44694_new_n3074_), .B(_abc_44694_new_n1114__bF_buf1), .Y(_abc_44694_new_n3075_));
OR2X2 OR2X2_901 ( .A(_abc_44694_new_n3076_), .B(_abc_44694_new_n1178__bF_buf0), .Y(_abc_44694_new_n3077_));
OR2X2 OR2X2_902 ( .A(_abc_44694_new_n1734_), .B(_abc_44694_new_n1179__bF_buf2), .Y(_abc_44694_new_n3078_));
OR2X2 OR2X2_903 ( .A(_abc_44694_new_n3079_), .B(_abc_44694_new_n3080_), .Y(alu_input_a_r_11_));
OR2X2 OR2X2_904 ( .A(_abc_44694_new_n3082_), .B(_abc_44694_new_n3084_), .Y(_abc_44694_new_n3085_));
OR2X2 OR2X2_905 ( .A(_abc_44694_new_n3086_), .B(_abc_44694_new_n3085_), .Y(_abc_44694_new_n3087_));
OR2X2 OR2X2_906 ( .A(_abc_44694_new_n3087_), .B(_abc_44694_new_n3088_), .Y(alu_input_a_r_12_));
OR2X2 OR2X2_907 ( .A(_abc_44694_new_n3090_), .B(_abc_44694_new_n3092_), .Y(_abc_44694_new_n3093_));
OR2X2 OR2X2_908 ( .A(_abc_44694_new_n3094_), .B(_abc_44694_new_n3093_), .Y(_abc_44694_new_n3095_));
OR2X2 OR2X2_909 ( .A(_abc_44694_new_n3095_), .B(_abc_44694_new_n3096_), .Y(alu_input_a_r_13_));
OR2X2 OR2X2_91 ( .A(_abc_44694_new_n866_), .B(_abc_44694_new_n817__bF_buf0), .Y(_abc_44694_new_n867_));
OR2X2 OR2X2_910 ( .A(_abc_44694_new_n3098_), .B(_abc_44694_new_n3100_), .Y(_abc_44694_new_n3101_));
OR2X2 OR2X2_911 ( .A(_abc_44694_new_n3102_), .B(_abc_44694_new_n3101_), .Y(_abc_44694_new_n3103_));
OR2X2 OR2X2_912 ( .A(_abc_44694_new_n3103_), .B(_abc_44694_new_n3104_), .Y(alu_input_a_r_14_));
OR2X2 OR2X2_913 ( .A(_abc_44694_new_n3106_), .B(_abc_44694_new_n3108_), .Y(_abc_44694_new_n3109_));
OR2X2 OR2X2_914 ( .A(_abc_44694_new_n3110_), .B(_abc_44694_new_n3109_), .Y(_abc_44694_new_n3111_));
OR2X2 OR2X2_915 ( .A(_abc_44694_new_n3111_), .B(_abc_44694_new_n3112_), .Y(alu_input_a_r_15_));
OR2X2 OR2X2_916 ( .A(_abc_44694_new_n1924_), .B(_abc_44694_new_n1179__bF_buf1), .Y(_abc_44694_new_n3114_));
OR2X2 OR2X2_917 ( .A(_abc_44694_new_n3116_), .B(_abc_44694_new_n3117_), .Y(_abc_44694_new_n3118_));
OR2X2 OR2X2_918 ( .A(_abc_44694_new_n3120_), .B(_abc_44694_new_n1178__bF_buf0), .Y(_abc_44694_new_n3121_));
OR2X2 OR2X2_919 ( .A(_abc_44694_new_n3118_), .B(_abc_44694_new_n3121_), .Y(_abc_44694_new_n3122_));
OR2X2 OR2X2_92 ( .A(_abc_44694_new_n872_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n873_));
OR2X2 OR2X2_920 ( .A(_abc_44694_new_n3123_), .B(_abc_44694_new_n3124_), .Y(alu_input_a_r_16_));
OR2X2 OR2X2_921 ( .A(_abc_44694_new_n1970_), .B(_abc_44694_new_n1179__bF_buf0), .Y(_abc_44694_new_n3126_));
OR2X2 OR2X2_922 ( .A(_abc_44694_new_n3128_), .B(_abc_44694_new_n3129_), .Y(_abc_44694_new_n3130_));
OR2X2 OR2X2_923 ( .A(_abc_44694_new_n3132_), .B(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n3133_));
OR2X2 OR2X2_924 ( .A(_abc_44694_new_n3130_), .B(_abc_44694_new_n3133_), .Y(_abc_44694_new_n3134_));
OR2X2 OR2X2_925 ( .A(_abc_44694_new_n3135_), .B(_abc_44694_new_n3136_), .Y(alu_input_a_r_17_));
OR2X2 OR2X2_926 ( .A(_abc_44694_new_n2006_), .B(_abc_44694_new_n1179__bF_buf3), .Y(_abc_44694_new_n3138_));
OR2X2 OR2X2_927 ( .A(_abc_44694_new_n3140_), .B(_abc_44694_new_n3141_), .Y(_abc_44694_new_n3142_));
OR2X2 OR2X2_928 ( .A(_abc_44694_new_n3144_), .B(_abc_44694_new_n1178__bF_buf3), .Y(_abc_44694_new_n3145_));
OR2X2 OR2X2_929 ( .A(_abc_44694_new_n3142_), .B(_abc_44694_new_n3145_), .Y(_abc_44694_new_n3146_));
OR2X2 OR2X2_93 ( .A(_abc_44694_new_n874_), .B(_abc_44694_new_n817__bF_buf3), .Y(_abc_44694_new_n875_));
OR2X2 OR2X2_930 ( .A(_abc_44694_new_n3147_), .B(_abc_44694_new_n3148_), .Y(alu_input_a_r_18_));
OR2X2 OR2X2_931 ( .A(_abc_44694_new_n2042_), .B(_abc_44694_new_n1179__bF_buf2), .Y(_abc_44694_new_n3150_));
OR2X2 OR2X2_932 ( .A(_abc_44694_new_n3152_), .B(_abc_44694_new_n3153_), .Y(_abc_44694_new_n3154_));
OR2X2 OR2X2_933 ( .A(_abc_44694_new_n3156_), .B(_abc_44694_new_n1178__bF_buf2), .Y(_abc_44694_new_n3157_));
OR2X2 OR2X2_934 ( .A(_abc_44694_new_n3154_), .B(_abc_44694_new_n3157_), .Y(_abc_44694_new_n3158_));
OR2X2 OR2X2_935 ( .A(_abc_44694_new_n3159_), .B(_abc_44694_new_n3160_), .Y(alu_input_a_r_19_));
OR2X2 OR2X2_936 ( .A(_abc_44694_new_n2078_), .B(_abc_44694_new_n1179__bF_buf1), .Y(_abc_44694_new_n3162_));
OR2X2 OR2X2_937 ( .A(_abc_44694_new_n3164_), .B(_abc_44694_new_n3165_), .Y(_abc_44694_new_n3166_));
OR2X2 OR2X2_938 ( .A(_abc_44694_new_n3168_), .B(_abc_44694_new_n1178__bF_buf1), .Y(_abc_44694_new_n3169_));
OR2X2 OR2X2_939 ( .A(_abc_44694_new_n3166_), .B(_abc_44694_new_n3169_), .Y(_abc_44694_new_n3170_));
OR2X2 OR2X2_94 ( .A(state_q_1_bF_buf0_), .B(alu_p_o_16_), .Y(_abc_44694_new_n876_));
OR2X2 OR2X2_940 ( .A(_abc_44694_new_n3171_), .B(_abc_44694_new_n3172_), .Y(alu_input_a_r_20_));
OR2X2 OR2X2_941 ( .A(_abc_44694_new_n2127_), .B(_abc_44694_new_n1179__bF_buf0), .Y(_abc_44694_new_n3174_));
OR2X2 OR2X2_942 ( .A(_abc_44694_new_n3176_), .B(_abc_44694_new_n3177_), .Y(_abc_44694_new_n3178_));
OR2X2 OR2X2_943 ( .A(_abc_44694_new_n3180_), .B(_abc_44694_new_n1178__bF_buf0), .Y(_abc_44694_new_n3181_));
OR2X2 OR2X2_944 ( .A(_abc_44694_new_n3178_), .B(_abc_44694_new_n3181_), .Y(_abc_44694_new_n3182_));
OR2X2 OR2X2_945 ( .A(_abc_44694_new_n3183_), .B(_abc_44694_new_n3184_), .Y(alu_input_a_r_21_));
OR2X2 OR2X2_946 ( .A(_abc_44694_new_n2166_), .B(_abc_44694_new_n1179__bF_buf3), .Y(_abc_44694_new_n3186_));
OR2X2 OR2X2_947 ( .A(_abc_44694_new_n3188_), .B(_abc_44694_new_n3189_), .Y(_abc_44694_new_n3190_));
OR2X2 OR2X2_948 ( .A(_abc_44694_new_n3192_), .B(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n3193_));
OR2X2 OR2X2_949 ( .A(_abc_44694_new_n3190_), .B(_abc_44694_new_n3193_), .Y(_abc_44694_new_n3194_));
OR2X2 OR2X2_95 ( .A(_abc_44694_new_n878_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n879_));
OR2X2 OR2X2_950 ( .A(_abc_44694_new_n3195_), .B(_abc_44694_new_n3196_), .Y(alu_input_a_r_22_));
OR2X2 OR2X2_951 ( .A(_abc_44694_new_n2203_), .B(_abc_44694_new_n1179__bF_buf2), .Y(_abc_44694_new_n3198_));
OR2X2 OR2X2_952 ( .A(_abc_44694_new_n3200_), .B(_abc_44694_new_n3201_), .Y(_abc_44694_new_n3202_));
OR2X2 OR2X2_953 ( .A(_abc_44694_new_n3204_), .B(_abc_44694_new_n1178__bF_buf3), .Y(_abc_44694_new_n3205_));
OR2X2 OR2X2_954 ( .A(_abc_44694_new_n3202_), .B(_abc_44694_new_n3205_), .Y(_abc_44694_new_n3206_));
OR2X2 OR2X2_955 ( .A(_abc_44694_new_n3207_), .B(_abc_44694_new_n3208_), .Y(alu_input_a_r_23_));
OR2X2 OR2X2_956 ( .A(_abc_44694_new_n2239_), .B(_abc_44694_new_n1179__bF_buf1), .Y(_abc_44694_new_n3210_));
OR2X2 OR2X2_957 ( .A(_abc_44694_new_n3212_), .B(_abc_44694_new_n3213_), .Y(_abc_44694_new_n3214_));
OR2X2 OR2X2_958 ( .A(_abc_44694_new_n3216_), .B(_abc_44694_new_n1178__bF_buf2), .Y(_abc_44694_new_n3217_));
OR2X2 OR2X2_959 ( .A(_abc_44694_new_n3214_), .B(_abc_44694_new_n3217_), .Y(_abc_44694_new_n3218_));
OR2X2 OR2X2_96 ( .A(_abc_44694_new_n880_), .B(_abc_44694_new_n817__bF_buf2), .Y(_abc_44694_new_n881_));
OR2X2 OR2X2_960 ( .A(_abc_44694_new_n3219_), .B(_abc_44694_new_n3220_), .Y(alu_input_a_r_24_));
OR2X2 OR2X2_961 ( .A(_abc_44694_new_n2285_), .B(_abc_44694_new_n1179__bF_buf0), .Y(_abc_44694_new_n3222_));
OR2X2 OR2X2_962 ( .A(_abc_44694_new_n3224_), .B(_abc_44694_new_n3225_), .Y(_abc_44694_new_n3226_));
OR2X2 OR2X2_963 ( .A(_abc_44694_new_n3228_), .B(_abc_44694_new_n1178__bF_buf1), .Y(_abc_44694_new_n3229_));
OR2X2 OR2X2_964 ( .A(_abc_44694_new_n3226_), .B(_abc_44694_new_n3229_), .Y(_abc_44694_new_n3230_));
OR2X2 OR2X2_965 ( .A(_abc_44694_new_n3231_), .B(_abc_44694_new_n3232_), .Y(alu_input_a_r_25_));
OR2X2 OR2X2_966 ( .A(_abc_44694_new_n2324_), .B(_abc_44694_new_n1179__bF_buf3), .Y(_abc_44694_new_n3234_));
OR2X2 OR2X2_967 ( .A(_abc_44694_new_n3236_), .B(_abc_44694_new_n3237_), .Y(_abc_44694_new_n3238_));
OR2X2 OR2X2_968 ( .A(_abc_44694_new_n3240_), .B(_abc_44694_new_n1178__bF_buf0), .Y(_abc_44694_new_n3241_));
OR2X2 OR2X2_969 ( .A(_abc_44694_new_n3238_), .B(_abc_44694_new_n3241_), .Y(_abc_44694_new_n3242_));
OR2X2 OR2X2_97 ( .A(state_q_1_bF_buf4_), .B(alu_p_o_17_), .Y(_abc_44694_new_n882_));
OR2X2 OR2X2_970 ( .A(_abc_44694_new_n3243_), .B(_abc_44694_new_n3244_), .Y(alu_input_a_r_26_));
OR2X2 OR2X2_971 ( .A(_abc_44694_new_n2361_), .B(_abc_44694_new_n1179__bF_buf2), .Y(_abc_44694_new_n3246_));
OR2X2 OR2X2_972 ( .A(_abc_44694_new_n3248_), .B(_abc_44694_new_n3249_), .Y(_abc_44694_new_n3250_));
OR2X2 OR2X2_973 ( .A(_abc_44694_new_n3252_), .B(_abc_44694_new_n1178__bF_buf4), .Y(_abc_44694_new_n3253_));
OR2X2 OR2X2_974 ( .A(_abc_44694_new_n3250_), .B(_abc_44694_new_n3253_), .Y(_abc_44694_new_n3254_));
OR2X2 OR2X2_975 ( .A(_abc_44694_new_n3255_), .B(_abc_44694_new_n3256_), .Y(alu_input_a_r_27_));
OR2X2 OR2X2_976 ( .A(_abc_44694_new_n2400_), .B(_abc_44694_new_n1179__bF_buf1), .Y(_abc_44694_new_n3258_));
OR2X2 OR2X2_977 ( .A(_abc_44694_new_n3260_), .B(_abc_44694_new_n3261_), .Y(_abc_44694_new_n3262_));
OR2X2 OR2X2_978 ( .A(_abc_44694_new_n3264_), .B(_abc_44694_new_n1178__bF_buf3), .Y(_abc_44694_new_n3265_));
OR2X2 OR2X2_979 ( .A(_abc_44694_new_n3262_), .B(_abc_44694_new_n3265_), .Y(_abc_44694_new_n3266_));
OR2X2 OR2X2_98 ( .A(_abc_44694_new_n884_), .B(_abc_44694_new_n871_), .Y(_abc_44694_new_n885_));
OR2X2 OR2X2_980 ( .A(_abc_44694_new_n3267_), .B(_abc_44694_new_n3268_), .Y(alu_input_a_r_28_));
OR2X2 OR2X2_981 ( .A(_abc_44694_new_n2437_), .B(_abc_44694_new_n1179__bF_buf0), .Y(_abc_44694_new_n3270_));
OR2X2 OR2X2_982 ( .A(_abc_44694_new_n3272_), .B(_abc_44694_new_n3273_), .Y(_abc_44694_new_n3274_));
OR2X2 OR2X2_983 ( .A(_abc_44694_new_n3276_), .B(_abc_44694_new_n1178__bF_buf2), .Y(_abc_44694_new_n3277_));
OR2X2 OR2X2_984 ( .A(_abc_44694_new_n3274_), .B(_abc_44694_new_n3277_), .Y(_abc_44694_new_n3278_));
OR2X2 OR2X2_985 ( .A(_abc_44694_new_n3279_), .B(_abc_44694_new_n3280_), .Y(alu_input_a_r_29_));
OR2X2 OR2X2_986 ( .A(_abc_44694_new_n2473_), .B(_abc_44694_new_n1179__bF_buf3), .Y(_abc_44694_new_n3282_));
OR2X2 OR2X2_987 ( .A(_abc_44694_new_n3284_), .B(_abc_44694_new_n3285_), .Y(_abc_44694_new_n3286_));
OR2X2 OR2X2_988 ( .A(_abc_44694_new_n3288_), .B(_abc_44694_new_n1178__bF_buf1), .Y(_abc_44694_new_n3289_));
OR2X2 OR2X2_989 ( .A(_abc_44694_new_n3286_), .B(_abc_44694_new_n3289_), .Y(_abc_44694_new_n3290_));
OR2X2 OR2X2_99 ( .A(_abc_44694_new_n886_), .B(_abc_44694_new_n817__bF_buf1), .Y(_abc_44694_new_n887_));
OR2X2 OR2X2_990 ( .A(_abc_44694_new_n3291_), .B(_abc_44694_new_n3292_), .Y(alu_input_a_r_30_));
OR2X2 OR2X2_991 ( .A(_abc_44694_new_n2514_), .B(_abc_44694_new_n1179__bF_buf2), .Y(_abc_44694_new_n3294_));
OR2X2 OR2X2_992 ( .A(_abc_44694_new_n3296_), .B(_abc_44694_new_n3297_), .Y(_abc_44694_new_n3298_));
OR2X2 OR2X2_993 ( .A(_abc_44694_new_n3300_), .B(_abc_44694_new_n1178__bF_buf0), .Y(_abc_44694_new_n3301_));
OR2X2 OR2X2_994 ( .A(_abc_44694_new_n3298_), .B(_abc_44694_new_n3301_), .Y(_abc_44694_new_n3302_));
OR2X2 OR2X2_995 ( .A(_abc_44694_new_n3303_), .B(_abc_44694_new_n3304_), .Y(alu_input_a_r_31_));
OR2X2 OR2X2_996 ( .A(_abc_44694_new_n1155_), .B(_abc_44694_new_n1182_), .Y(_abc_44694_new_n3306_));
OR2X2 OR2X2_997 ( .A(_abc_44694_new_n3306_), .B(_abc_44694_new_n1078_), .Y(_abc_44694_new_n3307_));
OR2X2 OR2X2_998 ( .A(_abc_44694_new_n1148_), .B(_abc_44694_new_n1104_), .Y(_abc_44694_new_n3309_));
OR2X2 OR2X2_999 ( .A(_abc_44694_new_n3309_), .B(_abc_44694_new_n3308_), .Y(_abc_44694_new_n3310_));


endmodule