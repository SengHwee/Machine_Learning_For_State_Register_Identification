module aes_core(\bus_in[0] , \bus_in[1] , \bus_in[2] , \bus_in[3] , \bus_in[4] , \bus_in[5] , \bus_in[6] , \bus_in[7] , \bus_in[8] , \bus_in[9] , \bus_in[10] , \bus_in[11] , \bus_in[12] , \bus_in[13] , \bus_in[14] , \bus_in[15] , \bus_in[16] , \bus_in[17] , \bus_in[18] , \bus_in[19] , \bus_in[20] , \bus_in[21] , \bus_in[22] , \bus_in[23] , \bus_in[24] , \bus_in[25] , \bus_in[26] , \bus_in[27] , \bus_in[28] , \bus_in[29] , \bus_in[30] , \bus_in[31] , \iv_en[0] , \iv_en[1] , \iv_en[2] , \iv_en[3] , \iv_sel_rd[0] , \iv_sel_rd[1] , \iv_sel_rd[2] , \iv_sel_rd[3] , \key_en[0] , \key_en[1] , \key_en[2] , \key_en[3] , \key_sel_rd[0] , \key_sel_rd[1] , \data_type[0] , \data_type[1] , \addr[0] , \addr[1] , \op_mode[0] , \op_mode[1] , \aes_mode[0] , \aes_mode[1] , start, disable_core, write_en, read_en, first_block, rst_n, clk, \col_out[0] , \col_out[1] , \col_out[2] , \col_out[3] , \col_out[4] , \col_out[5] , \col_out[6] , \col_out[7] , \col_out[8] , \col_out[9] , \col_out[10] , \col_out[11] , \col_out[12] , \col_out[13] , \col_out[14] , \col_out[15] , \col_out[16] , \col_out[17] , \col_out[18] , \col_out[19] , \col_out[20] , \col_out[21] , \col_out[22] , \col_out[23] , \col_out[24] , \col_out[25] , \col_out[26] , \col_out[27] , \col_out[28] , \col_out[29] , \col_out[30] , \col_out[31] , \key_out[0] , \key_out[1] , \key_out[2] , \key_out[3] , \key_out[4] , \key_out[5] , \key_out[6] , \key_out[7] , \key_out[8] , \key_out[9] , \key_out[10] , \key_out[11] , \key_out[12] , \key_out[13] , \key_out[14] , \key_out[15] , \key_out[16] , \key_out[17] , \key_out[18] , \key_out[19] , \key_out[20] , \key_out[21] , \key_out[22] , \key_out[23] , \key_out[24] , \key_out[25] , \key_out[26] , \key_out[27] , \key_out[28] , \key_out[29] , \key_out[30] , \key_out[31] , \iv_out[0] , \iv_out[1] , \iv_out[2] , \iv_out[3] , \iv_out[4] , \iv_out[5] , \iv_out[6] , \iv_out[7] , \iv_out[8] , \iv_out[9] , \iv_out[10] , \iv_out[11] , \iv_out[12] , \iv_out[13] , \iv_out[14] , \iv_out[15] , \iv_out[16] , \iv_out[17] , \iv_out[18] , \iv_out[19] , \iv_out[20] , \iv_out[21] , \iv_out[22] , \iv_out[23] , \iv_out[24] , \iv_out[25] , \iv_out[26] , \iv_out[27] , \iv_out[28] , \iv_out[29] , \iv_out[30] , \iv_out[31] , end_aes);

wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__0_; 
wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__1_; 
wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__2_; 
wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__3_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1817; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1856; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1897; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1928; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_0_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_10_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_12_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_13_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_14_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_1_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_2_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_4_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_5_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_6_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_8_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_9_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n100_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n102_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n103_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n104_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n105_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n107_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n108_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n109_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n111_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n112_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n114_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n115_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n116_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n117_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n119_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n121_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n122_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n123_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n124_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n126_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n127_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n128_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n129_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n130_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n132_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n133_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n135_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n136_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n139_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n141_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n143_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n145_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n146_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n147_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n148_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n150_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n151_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n152_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n154_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n155_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n157_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n158_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n160_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n161_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n162_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n163_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n164_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n167_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n168_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n169_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n171_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n172_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n173_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n174_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n176_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n178_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n179_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n180_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n182_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n183_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n184_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n185_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n186_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n187_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n188_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n190_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n195_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n196_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n199_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n201_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n202_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n204_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n208_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n210_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n212_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n73_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n75_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n76_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n77_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n78_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n79_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n80_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n82_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n83_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n85_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n86_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n87_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n88_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n89_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n90_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n91_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n92_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n93_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n95_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n96_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n97_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n98_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n99_; 
wire AES_CORE_CONTROL_UNIT_bypass_key_en; 
wire AES_CORE_CONTROL_UNIT_bypass_rk; 
wire AES_CORE_CONTROL_UNIT_col_en_0_; 
wire AES_CORE_CONTROL_UNIT_col_en_1_; 
wire AES_CORE_CONTROL_UNIT_col_en_2_; 
wire AES_CORE_CONTROL_UNIT_col_en_3_; 
wire AES_CORE_CONTROL_UNIT_col_sel_0_; 
wire AES_CORE_CONTROL_UNIT_col_sel_1_; 
wire AES_CORE_CONTROL_UNIT_encrypt_decrypt; 
wire AES_CORE_CONTROL_UNIT_iv_cnt_en; 
wire AES_CORE_CONTROL_UNIT_key_derivation_en; 
wire AES_CORE_CONTROL_UNIT_key_en_0_; 
wire AES_CORE_CONTROL_UNIT_key_en_1_; 
wire AES_CORE_CONTROL_UNIT_key_en_2_; 
wire AES_CORE_CONTROL_UNIT_key_en_3_; 
wire AES_CORE_CONTROL_UNIT_key_gen; 
wire AES_CORE_CONTROL_UNIT_key_out_sel_0_; 
wire AES_CORE_CONTROL_UNIT_key_out_sel_1_; 
wire AES_CORE_CONTROL_UNIT_key_sel; 
wire AES_CORE_CONTROL_UNIT_last_round; 
wire AES_CORE_CONTROL_UNIT_mode_cbc; 
wire AES_CORE_CONTROL_UNIT_mode_ctr; 
wire AES_CORE_CONTROL_UNIT_rd_count_0_; 
wire AES_CORE_CONTROL_UNIT_rd_count_1_; 
wire AES_CORE_CONTROL_UNIT_rd_count_2_; 
wire AES_CORE_CONTROL_UNIT_rd_count_3_; 
wire AES_CORE_CONTROL_UNIT_rk_sel_0_; 
wire AES_CORE_CONTROL_UNIT_rk_sel_1_; 
wire AES_CORE_CONTROL_UNIT_sbox_sel_0_; 
wire AES_CORE_CONTROL_UNIT_sbox_sel_1_; 
wire AES_CORE_CONTROL_UNIT_sbox_sel_2_; 
wire AES_CORE_CONTROL_UNIT_state_0_; 
wire AES_CORE_CONTROL_UNIT_state_11_; 
wire AES_CORE_CONTROL_UNIT_state_12_; 
wire AES_CORE_CONTROL_UNIT_state_13_; 
wire AES_CORE_CONTROL_UNIT_state_14_; 
wire AES_CORE_CONTROL_UNIT_state_15_; 
wire AES_CORE_CONTROL_UNIT_state_1_; 
wire AES_CORE_CONTROL_UNIT_state_2_; 
wire AES_CORE_CONTROL_UNIT_state_3_; 
wire AES_CORE_CONTROL_UNIT_state_4_; 
wire AES_CORE_CONTROL_UNIT_state_6_; 
wire AES_CORE_CONTROL_UNIT_state_7_; 
wire AES_CORE_CONTROL_UNIT_state_8_; 
wire AES_CORE_CONTROL_UNIT_state_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n327_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n328_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n330_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n331_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n333_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n334_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n336_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n337_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n339_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n340_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n342_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n343_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n345_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n346_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n348_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n349_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n351_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n352_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n354_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n355_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n357_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n358_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n360_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n361_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n363_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n364_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n366_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n367_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n369_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n370_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n372_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n373_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n375_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n376_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n378_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n379_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n381_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n382_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n384_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n385_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n387_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n388_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n390_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n391_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n393_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n394_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n396_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n397_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n399_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n400_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n401_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n402_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n404_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n406_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n407_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n408_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n409_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n411_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n412_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n413_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n414_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n415_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n416_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n417_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n418_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n419_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n420_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n421_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n422_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n423_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n426_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n427_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n428_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n429_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n431_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n432_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n433_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n434_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n435_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n436_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n437_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n438_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n439_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n441_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n442_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n443_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n444_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n445_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n446_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n447_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n448_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n449_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n450_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n451_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n452_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n453_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n454_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n456_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n457_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n458_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n460_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n461_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n462_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n463_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n464_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n465_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n466_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n467_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n468_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n469_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n470_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n471_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n472_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n473_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n475_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n476_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n477_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n478_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n479_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n480_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n481_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n482_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n483_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n484_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n485_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n486_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n487_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n488_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n489_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n490_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n491_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n493_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n494_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n495_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n496_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n497_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n498_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n499_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n500_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n501_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n502_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n503_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n504_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n505_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n506_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n508_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n509_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n510_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n511_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n512_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n513_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n514_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n515_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n516_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n518_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n519_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n520_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n521_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n522_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n523_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n524_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n525_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n528_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n529_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n532_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n533_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n536_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n537_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n540_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n541_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n544_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n545_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n548_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n549_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n552_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n553_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n556_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n557_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n560_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n561_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n564_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n565_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n568_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n569_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n572_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n573_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n576_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n577_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n580_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n581_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n584_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n585_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n588_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n589_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n592_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n593_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n596_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n597_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n600_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n601_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n604_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n605_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n608_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n609_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n612_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n613_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n616_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n617_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n620_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n621_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n624_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n625_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n628_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n629_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n632_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n633_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n636_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n637_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n640_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n641_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n644_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n645_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n648_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n649_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n652_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n653_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n680_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n682_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n683_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n684_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n688_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n689_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n690_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n692_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n694_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_3_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n101_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n102_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n104_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n105_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n106_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n107_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n108_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n109_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n110_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n111_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n113_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n114_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n115_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n116_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n117_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n119_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n120_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n122_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n123_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n124_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n125_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n127_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n128_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n129_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n130_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n131_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n132_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n133_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n134_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n135_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n136_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n137_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n138_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n139_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n140_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n141_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n142_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n143_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n144_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n145_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n146_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n147_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n148_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n149_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n150_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n151_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n152_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n153_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n154_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n155_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n156_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n157_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n159_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n160_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n163_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n164_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n165_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n166_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n167_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n168_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n169_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n171_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n172_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n173_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n174_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n176_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n177_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n178_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n179_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n180_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n182_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n183_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n184_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n185_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n186_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n187_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n188_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n189_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n190_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n191_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n192_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n193_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n194_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n196_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n197_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n198_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n199_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n201_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n202_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n203_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n204_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n205_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n206_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n207_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n208_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n209_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n210_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n211_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n212_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n213_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n214_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n215_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n216_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n217_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n218_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n219_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n220_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n221_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n222_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n223_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n224_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n225_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n226_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n227_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n228_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n229_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n230_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n231_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n233_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n234_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n235_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n236_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n238_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n239_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n240_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n241_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n242_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n243_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n244_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n245_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n246_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n247_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n248_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n249_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n250_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n251_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n252_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n253_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n254_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n255_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n256_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n257_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n258_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n259_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n260_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n261_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n262_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n263_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n264_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n265_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n266_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n267_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n268_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n269_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n270_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n271_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n272_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n273_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n274_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n275_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n276_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n277_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n278_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n279_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n280_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n281_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n282_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n283_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n284_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n285_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n286_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n287_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n288_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n290_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n291_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n292_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n294_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n295_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n296_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n297_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n298_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n299_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n300_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n301_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n302_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n303_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n304_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n305_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n306_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n307_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n308_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n309_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n310_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n311_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n312_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n313_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n314_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n315_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n316_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n317_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n318_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n319_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n320_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n322_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n323_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n324_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n326_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n328_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n329_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n330_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n331_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n332_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n333_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n334_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n335_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n336_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n337_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n338_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n339_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n340_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n342_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n343_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n345_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n346_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n347_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n348_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n349_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n350_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n351_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n354_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n356_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n358_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n359_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n360_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n361_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n363_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n364_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n365_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n366_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n367_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n368_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n369_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n371_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n372_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n374_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n375_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n376_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n377_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n378_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n380_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n381_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n382_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n383_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n384_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n386_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n387_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n388_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n389_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n390_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n391_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n393_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n394_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n395_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n397_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n398_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n399_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n400_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n401_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n402_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n403_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n404_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n405_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n407_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n408_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n409_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n411_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n412_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n413_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n414_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n415_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n416_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n417_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n419_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n420_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n421_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n423_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n424_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n425_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n426_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n427_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n428_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n429_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n431_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n433_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n435_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n437_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n438_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n441_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n442_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n443_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n445_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n446_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n447_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n449_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n452_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n453_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n454_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n456_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n457_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n458_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n460_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n461_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n462_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n464_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n465_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n466_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n468_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n469_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n471_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n472_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n474_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n475_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n476_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n478_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n479_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n481_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n482_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n485_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n488_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n489_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n490_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n492_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n493_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n494_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n496_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n499_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n500_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n501_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n502_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n504_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n505_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n507_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n508_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n510_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n511_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n512_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n514_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n515_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n516_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n518_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n519_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n521_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n523_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n524_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n525_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n527_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n97_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n99_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__7_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__7_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__7_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__7_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n101_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n116_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n127_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n137_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n141_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n155_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n301_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n322_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n336_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n377_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n388_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n403_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n413_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n415_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n419_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n428_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n431_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n434_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n437_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n441_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n484_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n77_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n101_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n116_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n127_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n137_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n141_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n155_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n301_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n322_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n336_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n377_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n388_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n403_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n413_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n415_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n419_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n428_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n431_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n434_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n437_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n441_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n484_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n77_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n101_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n116_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n127_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n137_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n141_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n155_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n301_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n322_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n336_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n377_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n388_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n403_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n413_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n415_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n419_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n428_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n431_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n434_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n437_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n441_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n484_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n77_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n101_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n116_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n127_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n137_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n141_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n155_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n301_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n322_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n336_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n377_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n388_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n403_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n413_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n415_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n419_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n428_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n431_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n434_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n437_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n441_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n484_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n77_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n100_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n101_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n103_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n104_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n105_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n107_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n108_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n109_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n111_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n112_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n113_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n115_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n116_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n117_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n119_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n120_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n121_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n123_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n124_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n125_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n127_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n128_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n129_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n131_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n132_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n133_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n135_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n136_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n137_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n139_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n140_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n141_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n143_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n144_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n145_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n147_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n148_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n149_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n151_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n152_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n153_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n155_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n156_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n157_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n159_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n160_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n161_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n163_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n164_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n165_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n167_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n168_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n169_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n171_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n172_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n173_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n175_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n176_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n177_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n179_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n180_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n181_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n183_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n184_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n185_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n187_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n188_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n189_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n191_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n192_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n193_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n195_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n196_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n197_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n68_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n70_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n73_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n75_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n76_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n77_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n79_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n80_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n81_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n83_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n84_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n85_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n87_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n88_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n89_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n91_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n92_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n93_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n95_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n96_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n97_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n99_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_0_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_10_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_11_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_12_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_13_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_14_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_15_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_16_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_17_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_18_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_19_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_1_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_20_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_21_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_22_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_23_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_24_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_25_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_26_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_27_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_28_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_29_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_2_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_30_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_31_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_3_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_4_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_5_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_6_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_7_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_8_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_9_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n100_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n101_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n103_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n104_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n105_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n107_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n108_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n109_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n111_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n112_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n113_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n115_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n116_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n117_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n119_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n120_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n121_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n123_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n124_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n125_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n127_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n128_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n129_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n131_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n132_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n133_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n135_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n136_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n137_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n139_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n140_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n141_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n143_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n144_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n145_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n147_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n148_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n149_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n151_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n152_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n153_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n155_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n156_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n157_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n159_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n160_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n161_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n163_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n164_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n165_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n167_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n168_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n169_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n171_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n172_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n173_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n175_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n176_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n177_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n179_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n180_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n181_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n183_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n184_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n185_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n187_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n188_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n189_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n191_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n192_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n193_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n195_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n196_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n197_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n68_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n70_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n73_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n75_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n76_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n77_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n79_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n80_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n81_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n83_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n84_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n85_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n87_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n88_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n89_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n91_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n92_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n93_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n95_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n96_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n97_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n99_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__9_; 
wire AES_CORE_DATAPATH__0col_0__31_0__0_; 
wire AES_CORE_DATAPATH__0col_0__31_0__10_; 
wire AES_CORE_DATAPATH__0col_0__31_0__11_; 
wire AES_CORE_DATAPATH__0col_0__31_0__12_; 
wire AES_CORE_DATAPATH__0col_0__31_0__13_; 
wire AES_CORE_DATAPATH__0col_0__31_0__14_; 
wire AES_CORE_DATAPATH__0col_0__31_0__15_; 
wire AES_CORE_DATAPATH__0col_0__31_0__16_; 
wire AES_CORE_DATAPATH__0col_0__31_0__17_; 
wire AES_CORE_DATAPATH__0col_0__31_0__18_; 
wire AES_CORE_DATAPATH__0col_0__31_0__19_; 
wire AES_CORE_DATAPATH__0col_0__31_0__1_; 
wire AES_CORE_DATAPATH__0col_0__31_0__20_; 
wire AES_CORE_DATAPATH__0col_0__31_0__21_; 
wire AES_CORE_DATAPATH__0col_0__31_0__22_; 
wire AES_CORE_DATAPATH__0col_0__31_0__23_; 
wire AES_CORE_DATAPATH__0col_0__31_0__24_; 
wire AES_CORE_DATAPATH__0col_0__31_0__25_; 
wire AES_CORE_DATAPATH__0col_0__31_0__26_; 
wire AES_CORE_DATAPATH__0col_0__31_0__27_; 
wire AES_CORE_DATAPATH__0col_0__31_0__28_; 
wire AES_CORE_DATAPATH__0col_0__31_0__29_; 
wire AES_CORE_DATAPATH__0col_0__31_0__2_; 
wire AES_CORE_DATAPATH__0col_0__31_0__30_; 
wire AES_CORE_DATAPATH__0col_0__31_0__31_; 
wire AES_CORE_DATAPATH__0col_0__31_0__3_; 
wire AES_CORE_DATAPATH__0col_0__31_0__4_; 
wire AES_CORE_DATAPATH__0col_0__31_0__5_; 
wire AES_CORE_DATAPATH__0col_0__31_0__6_; 
wire AES_CORE_DATAPATH__0col_0__31_0__7_; 
wire AES_CORE_DATAPATH__0col_0__31_0__8_; 
wire AES_CORE_DATAPATH__0col_0__31_0__9_; 
wire AES_CORE_DATAPATH__0col_1__31_0__0_; 
wire AES_CORE_DATAPATH__0col_1__31_0__10_; 
wire AES_CORE_DATAPATH__0col_1__31_0__11_; 
wire AES_CORE_DATAPATH__0col_1__31_0__12_; 
wire AES_CORE_DATAPATH__0col_1__31_0__13_; 
wire AES_CORE_DATAPATH__0col_1__31_0__14_; 
wire AES_CORE_DATAPATH__0col_1__31_0__15_; 
wire AES_CORE_DATAPATH__0col_1__31_0__16_; 
wire AES_CORE_DATAPATH__0col_1__31_0__17_; 
wire AES_CORE_DATAPATH__0col_1__31_0__18_; 
wire AES_CORE_DATAPATH__0col_1__31_0__19_; 
wire AES_CORE_DATAPATH__0col_1__31_0__1_; 
wire AES_CORE_DATAPATH__0col_1__31_0__20_; 
wire AES_CORE_DATAPATH__0col_1__31_0__21_; 
wire AES_CORE_DATAPATH__0col_1__31_0__22_; 
wire AES_CORE_DATAPATH__0col_1__31_0__23_; 
wire AES_CORE_DATAPATH__0col_1__31_0__24_; 
wire AES_CORE_DATAPATH__0col_1__31_0__25_; 
wire AES_CORE_DATAPATH__0col_1__31_0__26_; 
wire AES_CORE_DATAPATH__0col_1__31_0__27_; 
wire AES_CORE_DATAPATH__0col_1__31_0__28_; 
wire AES_CORE_DATAPATH__0col_1__31_0__29_; 
wire AES_CORE_DATAPATH__0col_1__31_0__2_; 
wire AES_CORE_DATAPATH__0col_1__31_0__30_; 
wire AES_CORE_DATAPATH__0col_1__31_0__31_; 
wire AES_CORE_DATAPATH__0col_1__31_0__3_; 
wire AES_CORE_DATAPATH__0col_1__31_0__4_; 
wire AES_CORE_DATAPATH__0col_1__31_0__5_; 
wire AES_CORE_DATAPATH__0col_1__31_0__6_; 
wire AES_CORE_DATAPATH__0col_1__31_0__7_; 
wire AES_CORE_DATAPATH__0col_1__31_0__8_; 
wire AES_CORE_DATAPATH__0col_1__31_0__9_; 
wire AES_CORE_DATAPATH__0col_2__31_0__0_; 
wire AES_CORE_DATAPATH__0col_2__31_0__10_; 
wire AES_CORE_DATAPATH__0col_2__31_0__11_; 
wire AES_CORE_DATAPATH__0col_2__31_0__12_; 
wire AES_CORE_DATAPATH__0col_2__31_0__13_; 
wire AES_CORE_DATAPATH__0col_2__31_0__14_; 
wire AES_CORE_DATAPATH__0col_2__31_0__15_; 
wire AES_CORE_DATAPATH__0col_2__31_0__16_; 
wire AES_CORE_DATAPATH__0col_2__31_0__17_; 
wire AES_CORE_DATAPATH__0col_2__31_0__18_; 
wire AES_CORE_DATAPATH__0col_2__31_0__19_; 
wire AES_CORE_DATAPATH__0col_2__31_0__1_; 
wire AES_CORE_DATAPATH__0col_2__31_0__20_; 
wire AES_CORE_DATAPATH__0col_2__31_0__21_; 
wire AES_CORE_DATAPATH__0col_2__31_0__22_; 
wire AES_CORE_DATAPATH__0col_2__31_0__23_; 
wire AES_CORE_DATAPATH__0col_2__31_0__24_; 
wire AES_CORE_DATAPATH__0col_2__31_0__25_; 
wire AES_CORE_DATAPATH__0col_2__31_0__26_; 
wire AES_CORE_DATAPATH__0col_2__31_0__27_; 
wire AES_CORE_DATAPATH__0col_2__31_0__28_; 
wire AES_CORE_DATAPATH__0col_2__31_0__29_; 
wire AES_CORE_DATAPATH__0col_2__31_0__2_; 
wire AES_CORE_DATAPATH__0col_2__31_0__30_; 
wire AES_CORE_DATAPATH__0col_2__31_0__31_; 
wire AES_CORE_DATAPATH__0col_2__31_0__3_; 
wire AES_CORE_DATAPATH__0col_2__31_0__4_; 
wire AES_CORE_DATAPATH__0col_2__31_0__5_; 
wire AES_CORE_DATAPATH__0col_2__31_0__6_; 
wire AES_CORE_DATAPATH__0col_2__31_0__7_; 
wire AES_CORE_DATAPATH__0col_2__31_0__8_; 
wire AES_CORE_DATAPATH__0col_2__31_0__9_; 
wire AES_CORE_DATAPATH__0col_3__31_0__0_; 
wire AES_CORE_DATAPATH__0col_3__31_0__10_; 
wire AES_CORE_DATAPATH__0col_3__31_0__11_; 
wire AES_CORE_DATAPATH__0col_3__31_0__12_; 
wire AES_CORE_DATAPATH__0col_3__31_0__13_; 
wire AES_CORE_DATAPATH__0col_3__31_0__14_; 
wire AES_CORE_DATAPATH__0col_3__31_0__15_; 
wire AES_CORE_DATAPATH__0col_3__31_0__16_; 
wire AES_CORE_DATAPATH__0col_3__31_0__17_; 
wire AES_CORE_DATAPATH__0col_3__31_0__18_; 
wire AES_CORE_DATAPATH__0col_3__31_0__19_; 
wire AES_CORE_DATAPATH__0col_3__31_0__1_; 
wire AES_CORE_DATAPATH__0col_3__31_0__20_; 
wire AES_CORE_DATAPATH__0col_3__31_0__21_; 
wire AES_CORE_DATAPATH__0col_3__31_0__22_; 
wire AES_CORE_DATAPATH__0col_3__31_0__23_; 
wire AES_CORE_DATAPATH__0col_3__31_0__24_; 
wire AES_CORE_DATAPATH__0col_3__31_0__25_; 
wire AES_CORE_DATAPATH__0col_3__31_0__26_; 
wire AES_CORE_DATAPATH__0col_3__31_0__27_; 
wire AES_CORE_DATAPATH__0col_3__31_0__28_; 
wire AES_CORE_DATAPATH__0col_3__31_0__29_; 
wire AES_CORE_DATAPATH__0col_3__31_0__2_; 
wire AES_CORE_DATAPATH__0col_3__31_0__30_; 
wire AES_CORE_DATAPATH__0col_3__31_0__31_; 
wire AES_CORE_DATAPATH__0col_3__31_0__3_; 
wire AES_CORE_DATAPATH__0col_3__31_0__4_; 
wire AES_CORE_DATAPATH__0col_3__31_0__5_; 
wire AES_CORE_DATAPATH__0col_3__31_0__6_; 
wire AES_CORE_DATAPATH__0col_3__31_0__7_; 
wire AES_CORE_DATAPATH__0col_3__31_0__8_; 
wire AES_CORE_DATAPATH__0col_3__31_0__9_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__0_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__1_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__2_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__3_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__0_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__1_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__2_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__3_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__9_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__9_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__9_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__9_; 
wire AES_CORE_DATAPATH__0key_0__31_0__0_; 
wire AES_CORE_DATAPATH__0key_0__31_0__10_; 
wire AES_CORE_DATAPATH__0key_0__31_0__11_; 
wire AES_CORE_DATAPATH__0key_0__31_0__12_; 
wire AES_CORE_DATAPATH__0key_0__31_0__13_; 
wire AES_CORE_DATAPATH__0key_0__31_0__14_; 
wire AES_CORE_DATAPATH__0key_0__31_0__15_; 
wire AES_CORE_DATAPATH__0key_0__31_0__16_; 
wire AES_CORE_DATAPATH__0key_0__31_0__17_; 
wire AES_CORE_DATAPATH__0key_0__31_0__18_; 
wire AES_CORE_DATAPATH__0key_0__31_0__19_; 
wire AES_CORE_DATAPATH__0key_0__31_0__1_; 
wire AES_CORE_DATAPATH__0key_0__31_0__20_; 
wire AES_CORE_DATAPATH__0key_0__31_0__21_; 
wire AES_CORE_DATAPATH__0key_0__31_0__22_; 
wire AES_CORE_DATAPATH__0key_0__31_0__23_; 
wire AES_CORE_DATAPATH__0key_0__31_0__24_; 
wire AES_CORE_DATAPATH__0key_0__31_0__25_; 
wire AES_CORE_DATAPATH__0key_0__31_0__26_; 
wire AES_CORE_DATAPATH__0key_0__31_0__27_; 
wire AES_CORE_DATAPATH__0key_0__31_0__28_; 
wire AES_CORE_DATAPATH__0key_0__31_0__29_; 
wire AES_CORE_DATAPATH__0key_0__31_0__2_; 
wire AES_CORE_DATAPATH__0key_0__31_0__30_; 
wire AES_CORE_DATAPATH__0key_0__31_0__31_; 
wire AES_CORE_DATAPATH__0key_0__31_0__3_; 
wire AES_CORE_DATAPATH__0key_0__31_0__4_; 
wire AES_CORE_DATAPATH__0key_0__31_0__5_; 
wire AES_CORE_DATAPATH__0key_0__31_0__6_; 
wire AES_CORE_DATAPATH__0key_0__31_0__7_; 
wire AES_CORE_DATAPATH__0key_0__31_0__8_; 
wire AES_CORE_DATAPATH__0key_0__31_0__9_; 
wire AES_CORE_DATAPATH__0key_1__31_0__0_; 
wire AES_CORE_DATAPATH__0key_1__31_0__10_; 
wire AES_CORE_DATAPATH__0key_1__31_0__11_; 
wire AES_CORE_DATAPATH__0key_1__31_0__12_; 
wire AES_CORE_DATAPATH__0key_1__31_0__13_; 
wire AES_CORE_DATAPATH__0key_1__31_0__14_; 
wire AES_CORE_DATAPATH__0key_1__31_0__15_; 
wire AES_CORE_DATAPATH__0key_1__31_0__16_; 
wire AES_CORE_DATAPATH__0key_1__31_0__17_; 
wire AES_CORE_DATAPATH__0key_1__31_0__18_; 
wire AES_CORE_DATAPATH__0key_1__31_0__19_; 
wire AES_CORE_DATAPATH__0key_1__31_0__1_; 
wire AES_CORE_DATAPATH__0key_1__31_0__20_; 
wire AES_CORE_DATAPATH__0key_1__31_0__21_; 
wire AES_CORE_DATAPATH__0key_1__31_0__22_; 
wire AES_CORE_DATAPATH__0key_1__31_0__23_; 
wire AES_CORE_DATAPATH__0key_1__31_0__24_; 
wire AES_CORE_DATAPATH__0key_1__31_0__25_; 
wire AES_CORE_DATAPATH__0key_1__31_0__26_; 
wire AES_CORE_DATAPATH__0key_1__31_0__27_; 
wire AES_CORE_DATAPATH__0key_1__31_0__28_; 
wire AES_CORE_DATAPATH__0key_1__31_0__29_; 
wire AES_CORE_DATAPATH__0key_1__31_0__2_; 
wire AES_CORE_DATAPATH__0key_1__31_0__30_; 
wire AES_CORE_DATAPATH__0key_1__31_0__31_; 
wire AES_CORE_DATAPATH__0key_1__31_0__3_; 
wire AES_CORE_DATAPATH__0key_1__31_0__4_; 
wire AES_CORE_DATAPATH__0key_1__31_0__5_; 
wire AES_CORE_DATAPATH__0key_1__31_0__6_; 
wire AES_CORE_DATAPATH__0key_1__31_0__7_; 
wire AES_CORE_DATAPATH__0key_1__31_0__8_; 
wire AES_CORE_DATAPATH__0key_1__31_0__9_; 
wire AES_CORE_DATAPATH__0key_2__31_0__0_; 
wire AES_CORE_DATAPATH__0key_2__31_0__10_; 
wire AES_CORE_DATAPATH__0key_2__31_0__11_; 
wire AES_CORE_DATAPATH__0key_2__31_0__12_; 
wire AES_CORE_DATAPATH__0key_2__31_0__13_; 
wire AES_CORE_DATAPATH__0key_2__31_0__14_; 
wire AES_CORE_DATAPATH__0key_2__31_0__15_; 
wire AES_CORE_DATAPATH__0key_2__31_0__16_; 
wire AES_CORE_DATAPATH__0key_2__31_0__17_; 
wire AES_CORE_DATAPATH__0key_2__31_0__18_; 
wire AES_CORE_DATAPATH__0key_2__31_0__19_; 
wire AES_CORE_DATAPATH__0key_2__31_0__1_; 
wire AES_CORE_DATAPATH__0key_2__31_0__20_; 
wire AES_CORE_DATAPATH__0key_2__31_0__21_; 
wire AES_CORE_DATAPATH__0key_2__31_0__22_; 
wire AES_CORE_DATAPATH__0key_2__31_0__23_; 
wire AES_CORE_DATAPATH__0key_2__31_0__24_; 
wire AES_CORE_DATAPATH__0key_2__31_0__25_; 
wire AES_CORE_DATAPATH__0key_2__31_0__26_; 
wire AES_CORE_DATAPATH__0key_2__31_0__27_; 
wire AES_CORE_DATAPATH__0key_2__31_0__28_; 
wire AES_CORE_DATAPATH__0key_2__31_0__29_; 
wire AES_CORE_DATAPATH__0key_2__31_0__2_; 
wire AES_CORE_DATAPATH__0key_2__31_0__30_; 
wire AES_CORE_DATAPATH__0key_2__31_0__31_; 
wire AES_CORE_DATAPATH__0key_2__31_0__3_; 
wire AES_CORE_DATAPATH__0key_2__31_0__4_; 
wire AES_CORE_DATAPATH__0key_2__31_0__5_; 
wire AES_CORE_DATAPATH__0key_2__31_0__6_; 
wire AES_CORE_DATAPATH__0key_2__31_0__7_; 
wire AES_CORE_DATAPATH__0key_2__31_0__8_; 
wire AES_CORE_DATAPATH__0key_2__31_0__9_; 
wire AES_CORE_DATAPATH__0key_3__31_0__0_; 
wire AES_CORE_DATAPATH__0key_3__31_0__10_; 
wire AES_CORE_DATAPATH__0key_3__31_0__11_; 
wire AES_CORE_DATAPATH__0key_3__31_0__12_; 
wire AES_CORE_DATAPATH__0key_3__31_0__13_; 
wire AES_CORE_DATAPATH__0key_3__31_0__14_; 
wire AES_CORE_DATAPATH__0key_3__31_0__15_; 
wire AES_CORE_DATAPATH__0key_3__31_0__16_; 
wire AES_CORE_DATAPATH__0key_3__31_0__17_; 
wire AES_CORE_DATAPATH__0key_3__31_0__18_; 
wire AES_CORE_DATAPATH__0key_3__31_0__19_; 
wire AES_CORE_DATAPATH__0key_3__31_0__1_; 
wire AES_CORE_DATAPATH__0key_3__31_0__20_; 
wire AES_CORE_DATAPATH__0key_3__31_0__21_; 
wire AES_CORE_DATAPATH__0key_3__31_0__22_; 
wire AES_CORE_DATAPATH__0key_3__31_0__23_; 
wire AES_CORE_DATAPATH__0key_3__31_0__24_; 
wire AES_CORE_DATAPATH__0key_3__31_0__25_; 
wire AES_CORE_DATAPATH__0key_3__31_0__26_; 
wire AES_CORE_DATAPATH__0key_3__31_0__27_; 
wire AES_CORE_DATAPATH__0key_3__31_0__28_; 
wire AES_CORE_DATAPATH__0key_3__31_0__29_; 
wire AES_CORE_DATAPATH__0key_3__31_0__2_; 
wire AES_CORE_DATAPATH__0key_3__31_0__30_; 
wire AES_CORE_DATAPATH__0key_3__31_0__31_; 
wire AES_CORE_DATAPATH__0key_3__31_0__3_; 
wire AES_CORE_DATAPATH__0key_3__31_0__4_; 
wire AES_CORE_DATAPATH__0key_3__31_0__5_; 
wire AES_CORE_DATAPATH__0key_3__31_0__6_; 
wire AES_CORE_DATAPATH__0key_3__31_0__7_; 
wire AES_CORE_DATAPATH__0key_3__31_0__8_; 
wire AES_CORE_DATAPATH__0key_3__31_0__9_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__0_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__1_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__2_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__3_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__9_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__9_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__9_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__9_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__0_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__10_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__11_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__12_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__13_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__14_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__15_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__16_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__17_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__18_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__19_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__1_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__20_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__21_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__22_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__23_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__24_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__25_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__26_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__27_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__28_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__29_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__2_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__30_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__31_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__3_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__4_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__5_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__6_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__7_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__8_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__9_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2457_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2458_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2459_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2460_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2461_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2462_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2463_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2464_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2465_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2466_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2467_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2468_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2469_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2470_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2471_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2472_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2473_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2474_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2475_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2476_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2477_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2478_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2479_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2480_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2481_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2482_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2483_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2484_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2486_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2487_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2488_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2489_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2490_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2491_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2492_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2494_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2495_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2496_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2497_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2498_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2500_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2501_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2502_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2503_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2504_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2505_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2506_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2508_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2509_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2510_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2511_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2512_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2514_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2515_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2516_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2517_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2518_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2520_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2521_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2522_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2523_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2524_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2525_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2526_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2528_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2529_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2530_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2531_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2532_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2533_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2534_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2536_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2537_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2538_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2539_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2540_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2541_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2542_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2544_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2545_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2546_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2547_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2548_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2549_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2550_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2552_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2553_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2554_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2555_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2556_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2557_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2558_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2560_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2561_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2562_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2563_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2564_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2565_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2566_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2568_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2569_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2570_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2571_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2572_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2574_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2575_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2576_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2577_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2578_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2579_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2580_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2582_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2583_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2584_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2585_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2586_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2588_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2589_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2590_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2591_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2592_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2593_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2594_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2596_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2597_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2598_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2599_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2600_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2602_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2603_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2604_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2605_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2606_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2607_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2608_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2610_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2611_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2612_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2613_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2614_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2615_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2616_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2618_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2619_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2620_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2621_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2622_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2623_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2624_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2626_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2627_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2628_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2629_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2630_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2632_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2633_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2634_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2635_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2636_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2637_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2638_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2640_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2641_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2642_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2643_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2644_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2646_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2647_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2648_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2649_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2650_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2651_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2652_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2654_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2655_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2656_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2657_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2658_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2660_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2661_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2662_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2663_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2664_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2665_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2666_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2668_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2669_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2670_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2671_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2672_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2673_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2674_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2676_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2677_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2678_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2679_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2680_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2682_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2683_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2684_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2685_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2686_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2687_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2688_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2690_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2691_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2692_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2693_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2694_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2696_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2697_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2698_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2699_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2700_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2702_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2703_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2704_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2705_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2706_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2707_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2708_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2710_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2711_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2712_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2713_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2714_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2715_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2716_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2717_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2718_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2719_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2720_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2721_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2722_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2723_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2724_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2725_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2726_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2727_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2728_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2729_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2730_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2731_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2732_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2733_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2734_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2735_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2736_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2737_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2738_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2739_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2740_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2741_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2742_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2744_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2745_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2746_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2747_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2748_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2749_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2750_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2751_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2753_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2754_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2755_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2756_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2758_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2759_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2760_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2761_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2762_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2763_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2764_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2765_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2766_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2768_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2769_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2770_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2771_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2772_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2773_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2774_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2775_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2776_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2778_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2779_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2780_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2781_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2782_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2783_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2784_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2785_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2786_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2788_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2789_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2790_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2791_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2792_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2793_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2794_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2795_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2796_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2798_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2799_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2800_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2801_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2802_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2803_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2804_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2805_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2806_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2808_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2809_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2810_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2811_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2812_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2813_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2814_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2815_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2817_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2818_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2819_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2821_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2822_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2823_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2824_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2825_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2826_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2827_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2828_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2830_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2831_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2832_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2834_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2835_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2836_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2837_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2838_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2839_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2840_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2841_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2842_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2844_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2845_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2846_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2847_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2848_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2849_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2850_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2851_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2852_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2854_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2855_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2856_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2857_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2858_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2859_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2860_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2861_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2862_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2864_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2865_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2866_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2867_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2868_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2869_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2870_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2871_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2872_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2874_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2875_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2876_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2877_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2878_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2879_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2880_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2881_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2882_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2884_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2885_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2886_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2887_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2888_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2889_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2890_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2891_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2892_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2894_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2895_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2896_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2897_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2898_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2899_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2900_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2901_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2902_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2904_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2905_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2906_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2907_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2908_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2909_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2910_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2911_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2912_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2914_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2915_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2916_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2917_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2918_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2919_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2920_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2921_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2922_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2924_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2925_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2926_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2927_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2928_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2929_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2930_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2931_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2932_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2934_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2935_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2936_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2937_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2938_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2939_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2940_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2941_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2942_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2944_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2945_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2946_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2947_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2948_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2949_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2950_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2951_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2953_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2954_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2955_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2957_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2958_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2959_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2960_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2961_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2962_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2963_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2964_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2965_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2967_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2968_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2969_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2970_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2971_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2972_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2973_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2974_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2975_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2977_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2978_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2979_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2980_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2981_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2982_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2983_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2984_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2986_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2987_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2988_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2990_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2991_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2992_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2993_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2994_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2995_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2996_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2997_; 
wire AES_CORE_DATAPATH__abc_15863_new_n2999_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3000_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3001_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3003_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3004_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3005_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3006_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3007_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3008_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3009_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3010_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3011_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3013_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3014_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3015_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3016_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3017_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3018_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3019_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3020_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3021_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3023_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3024_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3025_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3026_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3027_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3028_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3029_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3030_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3031_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3033_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3034_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3035_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3036_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3037_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3038_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3039_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3040_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3041_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3043_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3044_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3045_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3046_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3047_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3048_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3049_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3050_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3051_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3053_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3054_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3055_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3056_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3057_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3058_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3059_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3060_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3061_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3063_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3064_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3065_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3066_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3067_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3068_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3069_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3070_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3071_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3073_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3074_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3075_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3076_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3077_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3078_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3079_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3080_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3081_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3082_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3083_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3084_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3085_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3086_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3087_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3088_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3089_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3090_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3091_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3092_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3093_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3094_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3095_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3096_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3097_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3098_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3099_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3100_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3101_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3102_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3103_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3104_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3105_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3106_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3107_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3108_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3109_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3110_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3111_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3112_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3113_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3115_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3116_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3117_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3118_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3119_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3120_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3121_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3122_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3124_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3125_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3126_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3127_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3128_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3129_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3130_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3131_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3132_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3133_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3134_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3135_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3136_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3138_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3139_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3140_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3141_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3142_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3143_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3144_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3146_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3147_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3148_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3149_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3150_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3151_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3152_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3153_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3154_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3155_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3156_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3157_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3158_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3160_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3161_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3162_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3163_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3164_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3165_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3166_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3168_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3169_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3170_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3171_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3172_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3173_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3174_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3175_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3176_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3177_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3178_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3179_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3180_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3181_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3183_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3184_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3185_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3186_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3187_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3188_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3189_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3191_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3192_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3193_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3194_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3195_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3196_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3197_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3198_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3199_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3200_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3201_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3202_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3203_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3205_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3206_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3207_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3208_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3209_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3210_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3211_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3213_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3214_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3215_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3216_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3217_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3218_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3219_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3220_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3221_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3222_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3223_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3224_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3225_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3227_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3228_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3229_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3230_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3231_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3232_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3233_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3235_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3236_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3237_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3238_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3239_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3240_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3241_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3242_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3243_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3244_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3245_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3246_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3247_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3249_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3250_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3251_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3252_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3253_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3254_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3255_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3257_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3258_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3259_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3260_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3261_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3262_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3263_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3264_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3265_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3266_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3267_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3268_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3269_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3271_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3272_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3273_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3274_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3275_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3276_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3277_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3279_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3280_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3281_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3282_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3283_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3284_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3285_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3286_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3287_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3288_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3289_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3290_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3291_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3293_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3294_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3295_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3296_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3297_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3298_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3299_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3301_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3302_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3303_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3304_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3305_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3306_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3307_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3308_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3309_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3310_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3311_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3312_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3313_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3315_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3316_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3317_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3318_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3319_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3320_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3321_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3323_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3324_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3325_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3326_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3327_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3328_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3329_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3330_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3331_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3332_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3333_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3334_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3335_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3337_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3338_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3339_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3340_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3341_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3342_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3343_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3345_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3346_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3347_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3348_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3349_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3350_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3351_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3352_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3353_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3354_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3355_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3356_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3357_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3359_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3360_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3361_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3362_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3363_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3364_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3365_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3367_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3368_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3369_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3370_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3371_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3372_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3373_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3374_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3375_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3376_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3377_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3378_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3379_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3381_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3382_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3383_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3384_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3385_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3386_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3387_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3389_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3390_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3391_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3392_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3393_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3394_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3395_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3396_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3397_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3398_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3399_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3400_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3401_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3403_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3404_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3405_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3406_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3407_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3408_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3409_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3411_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3412_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3413_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3414_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3415_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3416_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3417_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3418_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3419_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3420_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3421_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3422_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3423_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3425_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3426_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3427_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3428_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3429_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3430_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3431_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3433_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3434_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3435_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3436_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3437_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3438_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3439_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3440_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3441_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3442_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3443_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3444_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3445_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3447_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3448_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3449_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3450_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3451_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3452_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3453_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3455_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3456_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3457_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3458_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3459_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3460_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3461_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3462_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3463_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3464_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3465_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3466_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3467_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3469_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3470_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3471_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3472_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3473_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3474_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3475_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3477_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3478_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3479_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3480_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3481_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3482_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3483_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3484_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3485_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3486_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3487_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3488_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3489_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3491_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3492_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3493_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3494_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3495_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3496_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3497_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3499_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3500_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3501_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3502_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3503_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3504_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3505_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3506_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3507_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3508_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3509_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3510_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3511_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3513_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3514_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3515_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3516_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3517_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3518_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3519_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3521_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3522_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3523_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3524_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3525_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3526_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3527_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3528_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3529_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3530_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3531_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3532_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3533_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3535_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3536_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3537_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3538_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3539_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3540_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3541_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3543_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3544_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3545_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3546_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3547_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3548_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3549_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3550_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3551_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3552_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3553_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3554_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3555_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3557_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3558_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3559_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3560_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3561_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3562_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3563_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3565_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3566_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3567_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3568_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3569_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3570_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3571_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3572_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3573_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3574_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3575_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3576_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3577_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3579_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3580_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3581_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3582_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3583_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3584_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3585_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3587_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3588_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3589_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3590_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3591_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3592_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3593_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3594_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3595_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3596_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3597_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3598_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3599_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3601_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3602_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3603_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3604_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3605_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3606_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3607_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3609_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3610_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3611_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3612_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3613_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3614_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3615_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3616_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3617_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3618_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3619_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3620_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3621_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3623_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3624_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3625_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3626_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3627_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3628_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3629_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3631_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3632_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3633_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3634_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3635_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3636_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3637_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3638_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3639_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3640_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3641_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3642_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3643_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3645_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3646_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3647_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3648_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3649_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3650_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3651_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3653_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3654_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3655_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3656_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3657_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3658_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3659_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3660_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3661_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3662_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3663_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3664_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3665_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3667_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3668_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3669_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3670_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3671_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3672_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3673_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3675_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3676_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3677_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3678_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3679_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3680_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3681_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3682_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3683_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3684_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3685_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3686_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3687_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3689_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3690_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3691_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3692_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3693_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3694_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3695_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3697_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3698_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3699_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3700_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3701_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3702_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3703_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3704_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3705_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3706_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3707_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3708_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3709_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3711_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3712_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3713_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3714_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3715_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3716_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3717_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3719_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3720_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3721_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3722_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3723_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3724_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3725_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3726_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3727_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3728_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3729_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3730_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3731_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3733_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3734_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3735_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3736_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3737_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3738_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3739_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3741_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3742_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3743_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3744_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3745_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3746_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3747_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3748_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3749_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3750_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3751_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3752_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3753_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3755_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3756_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3757_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3758_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3759_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3760_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3761_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3763_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3764_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3765_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3766_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3767_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3768_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3769_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3770_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3771_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3772_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3773_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3774_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3775_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3777_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3778_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3779_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3780_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3781_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3782_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3783_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3785_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3786_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3787_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3788_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3789_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3790_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3791_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3792_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3793_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3794_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3795_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3796_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3797_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3799_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3801_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3803_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3805_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3807_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3809_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3811_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3813_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3815_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3817_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3819_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3821_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3823_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3825_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3827_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3829_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3831_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3833_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3835_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3837_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3839_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3841_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3843_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3845_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3847_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3849_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3851_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3853_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3855_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3857_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3859_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3861_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3864_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3865_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3866_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3867_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3868_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3869_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3870_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3871_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3873_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3874_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3875_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3876_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3878_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3879_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3880_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3881_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3883_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3884_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3885_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3886_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3888_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3889_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3890_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3891_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3893_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3894_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3895_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3896_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3898_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3899_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3900_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3901_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3903_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3904_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3905_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3906_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3908_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3909_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3910_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3911_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3913_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3914_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3915_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3916_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3918_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3919_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3920_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3921_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3923_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3924_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3925_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3926_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3928_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3929_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3930_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3931_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3933_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3934_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3935_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3936_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3938_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3939_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3940_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3941_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3943_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3944_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3945_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3946_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3948_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3949_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3950_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3951_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3953_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3954_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3955_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3956_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3958_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3959_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3960_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3961_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3963_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3964_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3965_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3966_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3968_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3969_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3970_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3971_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3973_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3974_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3975_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3976_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3978_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3979_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3980_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3981_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3983_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3984_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3985_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3986_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3988_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3989_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3990_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3991_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3993_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3994_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3995_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3996_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3998_; 
wire AES_CORE_DATAPATH__abc_15863_new_n3999_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4000_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4001_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4003_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4004_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4005_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4006_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4008_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4009_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4010_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4011_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4013_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4014_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4015_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4016_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4018_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4019_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4020_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4021_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4023_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4024_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4025_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4026_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4027_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4028_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4030_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4031_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4032_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4033_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4034_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4035_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4036_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4037_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4038_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4040_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4041_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4042_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4043_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4045_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4046_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4047_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4048_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4050_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4051_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4052_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4053_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4055_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4056_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4057_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4058_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4060_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4061_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4062_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4063_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4065_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4066_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4067_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4068_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4070_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4071_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4072_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4073_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4075_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4076_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4077_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4078_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4080_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4081_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4082_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4083_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4085_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4086_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4087_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4088_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4090_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4091_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4092_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4093_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4095_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4096_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4097_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4098_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4100_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4101_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4102_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4103_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4105_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4106_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4107_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4108_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4110_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4111_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4112_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4113_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4115_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4116_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4117_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4118_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4120_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4121_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4122_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4123_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4125_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4126_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4127_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4128_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4130_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4131_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4132_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4133_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4135_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4136_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4137_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4138_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4140_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4141_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4142_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4143_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4145_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4146_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4147_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4148_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4150_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4151_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4152_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4153_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4155_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4156_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4157_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4158_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4160_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4161_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4162_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4163_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4165_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4166_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4167_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4168_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4170_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4171_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4172_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4173_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4175_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4176_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4177_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4178_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4180_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4181_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4182_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4183_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4185_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4186_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4187_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4188_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4190_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4191_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4192_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4193_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4194_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4196_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4198_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4230_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4231_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4232_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4233_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4235_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4236_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4237_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4238_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4240_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4241_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4242_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4243_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4245_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4246_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4247_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4248_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4250_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4251_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4252_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4253_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4255_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4256_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4257_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4258_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4260_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4261_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4263_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4264_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4266_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4267_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4269_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4270_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4272_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4273_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4275_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4276_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4278_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4279_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4280_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4281_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4283_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4284_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4285_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4286_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4288_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4289_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4290_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4291_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4293_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4294_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4295_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4296_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4298_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4299_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4300_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4301_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4303_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4304_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4305_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4306_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4308_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4309_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4310_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4311_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4313_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4314_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4315_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4316_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4318_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4319_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4320_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4321_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4323_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4324_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4325_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4326_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4328_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4329_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4330_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4331_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4333_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4334_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4335_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4336_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4338_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4339_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4340_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4341_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4343_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4344_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4345_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4346_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4348_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4349_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4350_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4351_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4353_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4354_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4355_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4356_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4358_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4359_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4360_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4361_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4363_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4364_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4365_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4366_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4368_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4369_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4370_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4371_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4373_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4374_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4376_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4378_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4380_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4382_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4384_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4386_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4388_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4390_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4392_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4394_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4396_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4398_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4400_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4402_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4404_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4406_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4408_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4410_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4412_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4414_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4416_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4418_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4420_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4422_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4424_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4426_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4428_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4430_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4432_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4434_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4436_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4438_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4440_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4441_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4442_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4443_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4444_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4445_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4447_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4448_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4449_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4451_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4452_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4453_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4455_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4456_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4457_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4459_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4460_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4461_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4463_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4464_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4465_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4467_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4468_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4469_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4471_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4472_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4473_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4475_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4476_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4477_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4479_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4480_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4481_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4483_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4484_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4485_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4487_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4488_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4489_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4491_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4492_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4493_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4495_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4496_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4497_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4499_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4500_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4501_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4503_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4504_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4505_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4507_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4508_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4509_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4511_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4512_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4513_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4515_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4516_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4517_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4519_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4520_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4521_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4523_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4524_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4525_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4527_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4528_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4529_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4531_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4532_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4533_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4535_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4536_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4537_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4539_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4540_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4541_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4543_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4544_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4545_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4547_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4548_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4549_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4551_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4552_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4553_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4555_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4556_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4557_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4559_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4560_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4561_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4563_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4564_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4565_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4567_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4568_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4569_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4571_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4572_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4573_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4574_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4575_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4576_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4577_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4578_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4579_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4580_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4581_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4582_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4583_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4584_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4585_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4586_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4587_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4588_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4589_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4590_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4591_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4592_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4593_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4594_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4595_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4596_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4597_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4598_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4599_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4600_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4601_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4602_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4603_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4604_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4605_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4606_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4607_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4608_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4609_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4610_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4611_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4612_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4613_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4614_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4615_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4616_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4617_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4618_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4619_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4620_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4621_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4622_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4623_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4624_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4625_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4626_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4627_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4628_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4629_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4630_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4631_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4633_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4634_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4635_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4636_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4637_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4638_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4639_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4640_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4641_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4642_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4643_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4644_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4645_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4646_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4647_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4648_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4649_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4650_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4651_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4652_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4653_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4654_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4655_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4656_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4657_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4658_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4659_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4660_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4661_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4662_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4663_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4664_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4665_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4666_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4667_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4668_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4669_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4670_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4672_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4673_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4674_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4675_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4676_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4677_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4678_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4679_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4680_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4681_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4682_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4683_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4684_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4685_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4686_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4687_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4688_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4689_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4690_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4691_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4692_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4693_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4694_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4695_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4696_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4697_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4698_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4699_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4700_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4701_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4702_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4703_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4704_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4705_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4706_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4707_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4708_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4709_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4711_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4712_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4713_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4714_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4715_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4716_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4717_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4718_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4719_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4720_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4721_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4722_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4723_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4724_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4725_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4726_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4727_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4728_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4729_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4730_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4731_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4732_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4733_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4734_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4735_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4736_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4737_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4738_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4739_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4740_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4741_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4742_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4743_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4744_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4745_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4746_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4747_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4748_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4749_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4751_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4752_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4753_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4754_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4755_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4756_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4757_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4758_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4759_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4760_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4761_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4762_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4763_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4764_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4765_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4766_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4767_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4768_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4769_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4770_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4771_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4772_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4773_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4774_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4775_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4776_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4777_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4778_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4779_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4780_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4781_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4782_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4783_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4784_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4785_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4787_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4788_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4789_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4790_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4791_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4792_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4793_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4794_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4795_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4796_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4797_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4798_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4799_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4800_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4801_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4802_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4803_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4804_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4805_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4806_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4807_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4808_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4809_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4810_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4811_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4812_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4813_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4814_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4815_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4816_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4817_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4818_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4819_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4820_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4821_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4822_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4823_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4824_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4826_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4827_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4828_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4829_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4830_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4831_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4832_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4833_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4834_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4835_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4836_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4837_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4838_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4839_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4840_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4841_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4842_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4843_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4844_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4845_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4846_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4847_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4848_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4849_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4850_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4851_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4852_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4853_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4854_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4855_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4856_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4857_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4858_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4859_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4861_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4862_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4863_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4864_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4865_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4866_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4867_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4868_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4869_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4870_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4871_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4872_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4873_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4874_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4875_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4876_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4877_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4878_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4879_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4880_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4881_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4882_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4883_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4884_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4885_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4886_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4887_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4888_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4889_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4890_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4891_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4892_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4893_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4894_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4895_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4896_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4897_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4898_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4900_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4901_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4902_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4903_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4904_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4905_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4906_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4907_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4908_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4909_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4910_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4911_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4912_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4913_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4914_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4915_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4916_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4917_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4918_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4919_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4920_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4921_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4922_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4923_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4924_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4925_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4926_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4927_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4928_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4929_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4930_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4931_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4932_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4933_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4935_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4936_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4937_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4938_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4939_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4940_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4941_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4942_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4943_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4944_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4945_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4946_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4947_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4948_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4949_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4950_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4951_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4952_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4953_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4954_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4955_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4956_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4957_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4958_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4959_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4960_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4961_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4962_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4963_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4964_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4965_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4966_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4967_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4968_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4969_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4970_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4971_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4972_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4974_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4975_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4976_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4977_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4978_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4979_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4980_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4981_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4982_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4983_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4984_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4985_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4986_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4987_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4988_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4989_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4990_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4991_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4992_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4993_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4994_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4995_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4996_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4997_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4998_; 
wire AES_CORE_DATAPATH__abc_15863_new_n4999_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5000_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5001_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5002_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5003_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5004_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5005_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5006_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5007_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5008_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5009_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5010_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5011_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5013_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5014_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5015_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5016_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5017_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5018_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5019_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5020_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5021_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5022_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5023_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5024_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5025_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5026_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5027_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5028_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5029_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5030_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5031_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5032_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5033_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5034_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5035_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5036_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5037_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5038_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5039_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5040_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5041_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5042_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5043_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5044_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5045_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5046_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5047_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5048_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5049_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5050_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5052_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5053_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5054_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5055_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5056_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5057_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5058_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5059_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5060_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5061_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5062_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5063_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5064_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5065_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5066_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5067_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5068_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5069_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5070_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5071_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5072_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5073_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5074_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5075_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5076_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5077_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5078_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5079_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5080_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5081_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5082_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5083_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5084_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5085_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5086_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5087_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5088_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5089_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5091_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5092_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5093_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5094_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5095_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5096_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5097_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5098_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5099_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5100_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5101_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5102_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5103_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5104_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5105_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5106_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5107_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5108_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5109_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5110_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5111_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5112_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5113_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5114_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5115_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5116_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5117_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5118_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5119_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5120_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5121_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5122_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5123_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5124_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5125_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5126_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5127_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5128_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5130_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5131_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5132_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5133_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5134_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5135_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5136_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5137_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5138_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5139_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5140_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5141_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5142_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5143_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5144_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5145_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5146_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5147_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5148_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5149_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5150_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5151_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5152_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5153_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5154_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5155_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5156_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5157_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5158_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5159_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5160_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5161_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5162_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5163_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5164_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5166_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5167_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5168_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5169_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5170_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5171_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5172_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5173_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5174_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5175_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5176_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5177_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5178_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5179_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5180_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5181_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5182_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5183_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5184_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5185_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5186_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5187_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5188_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5189_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5190_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5191_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5192_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5193_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5194_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5195_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5196_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5197_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5198_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5199_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5200_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5201_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5202_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5203_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5205_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5206_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5207_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5208_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5209_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5210_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5211_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5212_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5213_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5214_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5215_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5216_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5217_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5218_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5219_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5220_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5221_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5222_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5223_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5224_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5225_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5226_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5227_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5228_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5229_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5230_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5231_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5232_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5233_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5234_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5235_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5236_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5237_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5238_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5239_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5240_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5241_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5242_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5244_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5245_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5246_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5247_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5248_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5249_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5250_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5251_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5252_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5253_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5254_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5255_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5256_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5257_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5258_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5259_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5260_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5261_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5262_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5263_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5264_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5265_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5266_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5267_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5268_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5269_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5270_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5271_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5272_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5273_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5274_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5275_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5276_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5277_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5278_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5279_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5280_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5281_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5283_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5284_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5285_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5286_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5287_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5288_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5289_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5290_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5291_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5292_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5293_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5294_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5295_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5296_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5297_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5298_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5299_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5300_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5301_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5302_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5303_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5304_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5305_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5306_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5307_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5308_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5309_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5310_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5311_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5312_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5313_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5314_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5315_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5316_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5317_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5318_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5319_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5320_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5322_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5323_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5324_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5325_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5326_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5327_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5328_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5329_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5330_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5331_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5332_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5333_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5334_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5335_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5336_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5337_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5338_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5339_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5340_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5341_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5342_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5343_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5344_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5345_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5346_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5347_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5348_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5349_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5350_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5351_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5352_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5353_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5354_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5355_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5356_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5357_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5358_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5359_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5361_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5362_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5363_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5364_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5365_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5366_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5367_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5368_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5369_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5370_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5371_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5372_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5373_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5374_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5375_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5376_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5377_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5378_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5379_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5380_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5381_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5382_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5383_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5384_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5385_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5386_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5387_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5388_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5389_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5390_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5391_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5392_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5393_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5394_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5395_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5396_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5397_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5398_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5400_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5401_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5402_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5403_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5404_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5405_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5406_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5407_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5408_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5409_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5410_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5411_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5412_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5413_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5414_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5415_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5416_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5417_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5418_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5419_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5420_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5421_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5422_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5423_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5424_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5425_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5426_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5427_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5428_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5429_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5430_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5431_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5432_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5433_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5434_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5435_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5436_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5437_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5439_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5440_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5441_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5442_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5443_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5444_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5445_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5446_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5447_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5448_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5449_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5450_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5451_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5452_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5453_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5454_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5455_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5456_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5457_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5458_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5459_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5460_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5461_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5462_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5463_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5464_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5465_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5466_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5467_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5468_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5469_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5470_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5471_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5472_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5473_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5475_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5476_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5477_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5478_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5479_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5480_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5481_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5482_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5483_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5484_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5485_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5486_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5487_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5488_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5489_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5490_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5491_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5492_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5493_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5494_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5495_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5496_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5497_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5498_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5499_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5500_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5501_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5502_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5503_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5504_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5505_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5506_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5507_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5508_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5509_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5510_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5511_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5512_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5514_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5515_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5516_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5517_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5518_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5519_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5520_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5521_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5522_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5523_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5524_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5525_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5526_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5527_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5528_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5529_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5530_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5531_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5532_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5533_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5534_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5535_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5536_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5537_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5538_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5539_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5540_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5541_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5542_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5543_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5544_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5545_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5546_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5547_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5548_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5549_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5550_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5551_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5553_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5554_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5555_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5556_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5557_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5558_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5559_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5560_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5561_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5562_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5563_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5564_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5565_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5566_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5567_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5568_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5569_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5570_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5571_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5572_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5573_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5574_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5575_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5576_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5577_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5578_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5579_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5580_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5581_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5582_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5583_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5584_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5585_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5586_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5587_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5588_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5589_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5590_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5592_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5593_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5594_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5595_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5596_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5597_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5598_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5599_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5600_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5601_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5602_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5603_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5604_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5605_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5606_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5607_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5608_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5609_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5610_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5611_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5612_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5613_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5614_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5615_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5616_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5617_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5618_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5619_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5620_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5621_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5622_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5623_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5624_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5625_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5626_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5627_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5628_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5629_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5631_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5632_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5633_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5634_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5635_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5636_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5637_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5638_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5639_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5640_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5641_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5642_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5643_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5644_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5645_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5646_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5647_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5648_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5649_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5650_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5651_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5652_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5653_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5654_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5655_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5656_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5657_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5658_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5659_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5660_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5661_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5662_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5663_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5664_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5665_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5666_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5667_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5668_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5670_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5671_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5672_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5673_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5674_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5675_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5676_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5677_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5678_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5679_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5680_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5681_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5682_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5683_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5684_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5685_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5686_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5687_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5688_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5689_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5690_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5691_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5692_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5693_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5694_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5695_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5696_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5697_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5698_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5699_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5700_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5701_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5702_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5703_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5704_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5705_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5706_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5707_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5709_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5710_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5711_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5712_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5713_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5714_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5715_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5716_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5717_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5718_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5719_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5720_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5721_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5722_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5723_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5724_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5725_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5726_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5727_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5728_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5729_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5730_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5731_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5732_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5733_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5734_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5735_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5736_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5737_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5738_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5739_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5740_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5741_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5742_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5743_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5745_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5746_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5747_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5748_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5749_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5750_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5751_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5752_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5753_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5754_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5755_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5756_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5757_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5758_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5759_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5760_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5761_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5762_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5763_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5764_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5765_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5766_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5767_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5768_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5769_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5770_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5771_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5772_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5773_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5774_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5775_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5776_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5777_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5778_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5779_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5780_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5781_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5782_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5784_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5785_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5786_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5787_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5788_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5789_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5790_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5791_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5792_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5793_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5794_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5795_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5796_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5797_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5798_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5799_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5800_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5801_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5802_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5803_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5804_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5805_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5806_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5807_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5808_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5809_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5810_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5811_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5812_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5813_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5814_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5815_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5816_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5817_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5818_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5819_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5820_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5821_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5823_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5824_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5825_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5826_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5827_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5828_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5829_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5831_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5832_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5833_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5834_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5836_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5837_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5838_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5839_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5841_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5842_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5843_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5844_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5846_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5847_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5848_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5849_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5851_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5852_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5853_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5854_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5856_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5857_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5858_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5859_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5861_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5862_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5863_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5864_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5866_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5867_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5868_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5869_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5871_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5872_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5873_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5874_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5876_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5877_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5878_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5879_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5881_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5882_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5883_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5884_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5886_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5887_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5888_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5889_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5891_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5892_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5893_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5894_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5896_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5897_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5898_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5899_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5901_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5902_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5903_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5904_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5906_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5907_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5908_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5909_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5911_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5912_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5913_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5914_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5916_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5917_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5918_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5919_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5921_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5922_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5923_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5924_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5926_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5927_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5928_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5929_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5931_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5932_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5933_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5934_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5936_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5937_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5938_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5939_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5941_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5942_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5943_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5944_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5946_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5947_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5948_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5949_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5951_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5952_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5953_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5954_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5956_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5957_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5958_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5959_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5961_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5962_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5963_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5964_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5966_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5967_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5968_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5969_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5971_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5972_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5973_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5974_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5976_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5977_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5978_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5979_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5981_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5982_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5983_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5984_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5985_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5987_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5989_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5991_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5993_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5995_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5997_; 
wire AES_CORE_DATAPATH__abc_15863_new_n5999_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6001_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6003_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6005_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6007_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6009_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6011_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6013_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6015_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6017_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6019_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6021_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6023_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6025_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6027_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6029_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6031_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6033_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6035_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6037_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6039_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6041_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6043_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6045_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6047_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6049_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6051_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6052_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6053_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6054_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6055_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6056_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6058_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6059_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6060_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6061_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6062_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6063_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6065_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6066_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6067_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6068_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6069_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6070_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6072_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6073_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6074_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6075_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6076_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6077_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6079_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6080_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6081_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6082_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6083_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6084_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6086_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6087_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6088_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6089_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6090_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6091_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6093_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6094_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6095_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6096_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6097_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6098_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6100_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6101_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6102_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6103_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6104_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6105_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6107_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6108_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6109_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6110_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6111_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6112_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6114_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6115_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6116_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6117_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6118_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6119_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6121_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6122_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6123_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6124_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6125_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6126_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6128_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6129_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6130_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6131_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6132_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6133_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6135_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6136_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6137_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6138_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6139_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6140_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6142_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6143_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6144_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6145_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6146_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6147_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6149_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6150_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6151_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6152_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6153_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6154_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6156_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6157_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6158_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6159_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6160_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6161_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6163_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6164_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6165_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6166_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6167_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6168_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6170_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6171_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6172_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6173_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6174_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6175_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6177_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6178_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6179_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6180_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6181_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6182_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6184_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6185_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6186_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6187_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6188_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6189_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6191_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6192_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6193_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6194_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6195_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6196_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6198_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6199_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6200_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6201_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6202_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6203_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6205_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6206_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6207_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6208_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6209_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6210_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6212_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6213_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6214_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6215_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6216_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6217_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6219_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6220_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6221_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6222_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6223_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6224_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6226_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6227_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6228_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6229_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6230_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6231_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6233_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6234_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6235_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6236_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6237_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6238_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6240_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6241_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6242_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6243_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6244_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6245_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6247_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6248_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6249_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6250_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6251_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6252_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6254_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6255_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6256_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6257_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6258_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6259_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6261_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6262_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6263_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6264_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6265_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6266_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6268_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6269_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6270_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6271_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6272_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6273_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6275_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6276_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6277_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6278_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6279_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6280_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6282_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6283_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6284_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6285_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6286_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6287_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6289_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6290_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6291_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6292_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6293_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6294_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6296_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6297_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6298_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6299_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6300_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6301_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6303_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6304_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6305_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6306_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6307_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6308_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6310_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6311_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6312_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6313_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6314_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6315_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6317_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6318_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6319_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6320_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6321_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6322_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6324_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6325_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6326_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6327_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6328_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6329_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6331_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6332_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6333_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6334_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6335_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6336_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6338_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6339_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6340_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6341_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6342_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6343_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6345_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6346_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6347_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6348_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6349_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6350_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6352_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6353_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6354_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6355_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6356_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6357_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6359_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6360_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6361_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6362_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6363_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6364_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6366_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6367_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6368_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6369_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6370_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6371_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6373_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6374_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6375_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6376_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6377_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6378_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6380_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6381_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6382_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6383_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6384_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6385_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6387_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6388_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6389_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6390_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6391_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6392_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6394_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6395_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6396_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6397_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6398_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6399_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6401_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6402_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6403_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6404_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6405_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6406_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6408_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6409_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6410_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6411_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6412_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6413_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6415_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6416_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6417_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6418_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6419_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6420_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6422_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6423_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6424_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6425_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6426_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6427_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6429_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6430_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6431_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6432_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6433_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6434_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6436_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6437_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6438_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6439_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6440_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6441_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6443_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6444_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6445_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6446_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6447_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6448_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6450_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6451_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6452_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6453_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6454_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6455_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6457_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6458_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6459_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6460_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6461_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6462_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6464_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6465_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6466_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6467_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6468_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6469_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6471_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6472_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6473_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6474_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6475_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6476_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6478_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6479_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6480_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6481_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6482_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6483_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6485_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6486_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6487_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6488_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6489_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6490_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6492_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6493_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6494_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6495_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6496_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6497_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6499_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6500_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6501_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6502_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6503_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6504_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6505_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6507_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6508_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6509_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6510_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6511_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6513_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6514_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6515_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6516_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6517_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6518_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6520_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6521_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6522_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6523_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6524_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6526_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6527_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6528_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6529_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6530_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6531_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6533_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6534_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6535_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6536_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6537_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6538_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6540_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6541_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6542_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6543_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6544_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6545_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6547_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6548_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6549_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6550_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6551_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6553_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6554_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6555_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6556_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6557_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6558_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6560_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6561_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6562_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6563_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6564_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6566_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6567_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6568_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6569_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6570_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6571_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6573_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6574_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6575_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6576_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6577_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6579_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6580_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6581_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6582_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6583_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6584_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6586_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6587_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6588_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6589_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6590_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6592_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6593_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6594_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6595_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6596_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6597_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6599_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6600_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6601_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6602_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6603_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6605_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6606_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6607_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6608_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6609_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6610_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6612_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6613_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6614_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6615_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6616_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6618_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6619_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6620_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6621_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6622_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6624_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6625_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6626_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6627_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6628_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6630_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6631_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6632_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6633_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6634_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6635_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6637_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6638_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6639_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6640_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6641_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6643_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6644_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6645_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6646_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6647_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6648_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6650_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6651_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6652_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6653_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6654_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6656_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6657_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6658_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6659_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6660_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6661_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6663_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6664_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6665_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6666_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6667_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6669_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6670_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6671_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6672_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6673_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6675_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6676_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6677_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6678_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6679_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6680_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6682_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6683_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6684_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6685_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6686_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6688_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6689_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6690_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6691_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6692_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6693_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6695_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6696_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6697_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6698_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6699_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6700_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6702_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6703_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6704_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6705_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6706_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6708_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6709_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6710_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6711_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6712_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6713_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6714_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6716_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6718_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6720_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6722_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6724_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6726_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6728_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6730_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6732_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6734_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6736_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6738_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6740_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6742_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6744_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6746_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6748_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6750_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6752_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6754_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6756_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6758_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6760_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6762_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6764_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6766_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6768_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6770_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6772_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6774_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6776_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6778_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6779_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6780_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6781_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6782_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6783_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6785_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6786_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6787_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6788_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6789_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6791_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6792_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6793_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6794_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6795_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6797_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6798_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6799_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6800_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6801_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6803_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6804_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6805_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6806_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6807_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6808_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6810_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6811_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6812_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6813_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6814_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6816_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6817_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6818_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6819_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6820_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6821_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6823_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6824_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6825_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6826_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6827_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6829_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6830_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6831_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6832_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6833_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6834_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6836_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6837_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6838_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6839_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6840_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6842_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6843_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6844_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6845_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6846_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6848_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6849_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6850_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6851_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6852_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6854_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6855_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6856_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6857_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6858_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6860_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6861_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6862_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6863_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6864_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6866_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6867_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6868_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6869_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6870_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6871_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6873_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6874_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6875_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6876_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6877_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6879_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6880_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6881_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6882_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6883_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6885_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6886_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6887_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6888_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6889_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6891_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6892_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6893_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6894_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6895_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6897_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6898_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6899_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6900_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6901_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6903_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6904_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6905_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6906_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6907_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6909_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6910_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6911_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6912_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6913_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6915_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6916_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6917_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6918_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6919_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6920_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6922_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6923_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6924_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6925_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6926_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6928_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6929_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6930_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6931_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6932_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6934_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6935_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6936_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6937_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6938_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6940_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6941_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6942_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6943_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6944_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6946_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6947_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6948_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6949_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6950_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6952_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6953_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6954_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6955_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6956_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6958_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6959_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6960_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6961_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6962_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6963_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6965_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6966_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6967_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6968_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6969_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6971_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6972_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6973_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6974_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6975_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6977_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6978_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6979_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6980_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6981_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6982_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6983_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6985_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6986_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6987_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6988_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6989_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6990_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6991_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6993_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6994_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6995_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6996_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6997_; 
wire AES_CORE_DATAPATH__abc_15863_new_n6999_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7000_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7001_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7002_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7003_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7004_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7005_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7007_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7008_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7009_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7010_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7011_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7013_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7014_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7015_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7016_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7017_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7018_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7019_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7021_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7022_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7023_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7024_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7026_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7027_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7028_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7029_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7030_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7031_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7032_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7034_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7035_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7036_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7037_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7039_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7040_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7041_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7042_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7043_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7044_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7045_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7047_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7048_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7049_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7050_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7051_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7052_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7054_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7055_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7056_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7057_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7058_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7060_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7061_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7062_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7063_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7064_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7066_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7067_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7068_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7069_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7071_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7072_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7073_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7074_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7075_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7076_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7078_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7079_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7080_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7081_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7082_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7084_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7085_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7086_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7087_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7088_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7089_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7091_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7092_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7093_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7094_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7096_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7097_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7098_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7099_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7100_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7102_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7103_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7104_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7105_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7107_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7108_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7109_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7110_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7111_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7112_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7113_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7114_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7115_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7116_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7117_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7118_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7119_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7120_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7121_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7123_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7124_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7125_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7126_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7127_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7128_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7130_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7131_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7132_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7133_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7134_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7135_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7136_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7138_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7139_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7140_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7141_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7142_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7143_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7145_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7146_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7147_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7148_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7149_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7150_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7151_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7152_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7153_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7154_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7156_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7157_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7158_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7159_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7160_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7161_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7163_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7164_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7165_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7166_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7167_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7168_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7169_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7170_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7172_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7173_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7174_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7175_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7176_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7177_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7179_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7180_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7181_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7182_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7183_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7184_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7185_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7186_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7188_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7189_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7190_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7191_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7192_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7193_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7195_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7196_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7197_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7198_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7199_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7200_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7201_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7203_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7204_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7205_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7206_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7207_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7208_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7210_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7212_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7214_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7216_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7218_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7220_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7222_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7224_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7226_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7228_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7230_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7232_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7234_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7236_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7238_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7240_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7242_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7244_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7246_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7248_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7250_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7252_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7254_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7256_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7258_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7260_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7262_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7264_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7266_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7268_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7270_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7272_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7274_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7275_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7277_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7279_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7281_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7283_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7285_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7287_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7289_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7291_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7293_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7295_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7297_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7299_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7301_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7303_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7305_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7307_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7309_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7311_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7313_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7315_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7317_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7319_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7321_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7323_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7325_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7327_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7329_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7331_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7333_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7335_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7337_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7339_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7340_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7341_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7342_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7344_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7345_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7346_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7347_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7349_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7350_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7351_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7352_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7354_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7355_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7356_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7357_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7359_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7360_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7361_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7362_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7364_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7365_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7366_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7367_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7369_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7370_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7371_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7372_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7374_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7375_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7376_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7377_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7379_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7380_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7381_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7382_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7384_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7385_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7386_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7387_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7389_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7390_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7391_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7392_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7394_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7395_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7396_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7397_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7399_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7400_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7401_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7402_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7404_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7405_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7406_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7407_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7409_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7410_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7411_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7412_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7414_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7415_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7416_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7417_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7419_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7420_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7421_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7422_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7424_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7425_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7426_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7427_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7429_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7430_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7431_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7432_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7434_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7435_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7436_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7437_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7439_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7440_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7441_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7442_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7444_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7445_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7446_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7447_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7449_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7450_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7451_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7452_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7454_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7455_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7456_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7457_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7459_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7460_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7461_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7462_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7464_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7465_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7466_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7467_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7469_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7470_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7471_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7472_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7474_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7475_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7476_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7477_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7479_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7480_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7481_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7482_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7484_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7485_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7486_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7487_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7489_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7490_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7491_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7492_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7494_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7495_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7496_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7497_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7499_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7501_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7503_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7505_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7507_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7509_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7511_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7513_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7515_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7517_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7519_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7521_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7523_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7525_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7527_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7529_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7531_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7533_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7535_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7537_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7539_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7541_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7543_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7545_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7547_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7549_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7551_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7553_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7555_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7557_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7559_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7561_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7563_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7564_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7566_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7567_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7569_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7571_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7572_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7574_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7576_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7578_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7580_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7581_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7583_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7585_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7586_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7588_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7590_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7591_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7593_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7595_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7596_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7598_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7600_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7601_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7603_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7605_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7606_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7608_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7609_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7611_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7612_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7614_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7616_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7617_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7619_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7621_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7622_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7624_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7626_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7627_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7629_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7630_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7632_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7634_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7635_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7637_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7639_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7641_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7642_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7644_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7645_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7646_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7647_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7648_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7650_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7651_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7652_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7653_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7655_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7656_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7657_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7658_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7659_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7661_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7662_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7663_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7664_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7666_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7667_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7668_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7669_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7670_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7672_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7673_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7674_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7675_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7676_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7678_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7679_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7680_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7681_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7682_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7684_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7685_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7686_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7687_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7689_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7690_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7691_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7692_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7693_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7695_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7696_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7697_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7698_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7700_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7701_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7702_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7703_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7704_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7706_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7707_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7708_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7709_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7711_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7712_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7713_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7714_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7715_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7717_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7718_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7719_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7720_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7722_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7723_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7724_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7725_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7726_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7728_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7729_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7730_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7731_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7733_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7734_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7735_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7736_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7737_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7739_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7740_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7741_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7742_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7744_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7745_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7746_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7747_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7749_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7750_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7751_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7752_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7754_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7755_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7756_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7757_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7758_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7760_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7761_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7762_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7763_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7765_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7766_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7767_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7768_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7769_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7771_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7772_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7773_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7774_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7776_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7777_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7778_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7779_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7780_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7782_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7783_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7784_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7785_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7787_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7788_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7789_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7790_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7792_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7793_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7794_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7795_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7796_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7798_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7799_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7800_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7801_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7803_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7804_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7805_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7806_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7807_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7809_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7810_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7811_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7812_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7813_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7815_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7816_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7817_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7818_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7820_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7822_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7824_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7826_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7828_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7830_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7832_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7833_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7835_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7836_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7838_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7839_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7841_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7842_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7844_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7845_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7847_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7848_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7850_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7852_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7854_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7856_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7858_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7860_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7862_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7864_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7866_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7868_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7870_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7872_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7874_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7876_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7878_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7880_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7882_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7884_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7886_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7888_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7890_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7891_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7893_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7895_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7897_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7899_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7901_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7903_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7905_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7907_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7909_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7911_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7913_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7915_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7917_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7919_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7921_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7923_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7925_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7927_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7929_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7931_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7933_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7935_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7937_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7939_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7941_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7943_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7945_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7947_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7949_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7951_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7953_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7955_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7956_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7957_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7958_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7959_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7961_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7962_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7963_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7964_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7965_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7967_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7968_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7969_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7970_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7971_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7973_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7974_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7975_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7976_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7977_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7979_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7980_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7981_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7982_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7983_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7985_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7986_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7987_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7988_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7989_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7991_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7992_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7993_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7994_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7995_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7997_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7998_; 
wire AES_CORE_DATAPATH__abc_15863_new_n7999_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8000_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8001_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8003_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8004_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8005_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8006_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8007_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8009_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8010_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8011_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8012_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8013_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8015_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8016_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8017_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8018_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8019_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8021_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8022_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8023_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8024_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8025_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8027_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8028_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8029_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8030_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8031_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8033_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8034_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8035_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8036_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8037_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8039_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8040_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8041_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8042_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8043_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8045_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8046_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8047_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8048_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8049_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8051_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8052_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8053_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8054_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8055_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8057_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8058_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8059_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8060_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8061_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8063_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8064_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8065_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8066_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8067_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8069_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8070_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8071_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8072_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8073_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8075_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8076_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8077_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8078_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8079_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8081_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8082_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8083_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8084_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8085_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8087_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8088_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8089_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8090_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8091_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8093_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8094_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8095_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8096_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8097_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8099_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8100_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8101_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8102_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8103_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8105_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8106_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8107_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8108_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8109_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8111_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8112_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8113_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8114_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8115_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8117_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8118_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8119_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8120_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8121_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8123_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8124_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8125_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8126_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8127_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8129_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8130_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8131_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8132_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8133_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8135_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8136_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8137_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8138_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8139_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8141_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8142_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8143_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8144_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8145_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8147_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8148_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8150_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8151_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8153_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8154_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8156_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8157_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8159_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8161_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8162_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8164_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8165_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8167_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8168_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8170_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8172_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8174_; 
wire AES_CORE_DATAPATH__abc_15863_new_n8176_; 
wire AES_CORE_DATAPATH_bkp_0__0_; 
wire AES_CORE_DATAPATH_bkp_0__10_; 
wire AES_CORE_DATAPATH_bkp_0__11_; 
wire AES_CORE_DATAPATH_bkp_0__12_; 
wire AES_CORE_DATAPATH_bkp_0__13_; 
wire AES_CORE_DATAPATH_bkp_0__14_; 
wire AES_CORE_DATAPATH_bkp_0__15_; 
wire AES_CORE_DATAPATH_bkp_0__16_; 
wire AES_CORE_DATAPATH_bkp_0__17_; 
wire AES_CORE_DATAPATH_bkp_0__18_; 
wire AES_CORE_DATAPATH_bkp_0__19_; 
wire AES_CORE_DATAPATH_bkp_0__1_; 
wire AES_CORE_DATAPATH_bkp_0__20_; 
wire AES_CORE_DATAPATH_bkp_0__21_; 
wire AES_CORE_DATAPATH_bkp_0__22_; 
wire AES_CORE_DATAPATH_bkp_0__23_; 
wire AES_CORE_DATAPATH_bkp_0__24_; 
wire AES_CORE_DATAPATH_bkp_0__25_; 
wire AES_CORE_DATAPATH_bkp_0__26_; 
wire AES_CORE_DATAPATH_bkp_0__27_; 
wire AES_CORE_DATAPATH_bkp_0__28_; 
wire AES_CORE_DATAPATH_bkp_0__29_; 
wire AES_CORE_DATAPATH_bkp_0__2_; 
wire AES_CORE_DATAPATH_bkp_0__30_; 
wire AES_CORE_DATAPATH_bkp_0__31_; 
wire AES_CORE_DATAPATH_bkp_0__3_; 
wire AES_CORE_DATAPATH_bkp_0__4_; 
wire AES_CORE_DATAPATH_bkp_0__5_; 
wire AES_CORE_DATAPATH_bkp_0__6_; 
wire AES_CORE_DATAPATH_bkp_0__7_; 
wire AES_CORE_DATAPATH_bkp_0__8_; 
wire AES_CORE_DATAPATH_bkp_0__9_; 
wire AES_CORE_DATAPATH_bkp_1_0__0_; 
wire AES_CORE_DATAPATH_bkp_1_0__10_; 
wire AES_CORE_DATAPATH_bkp_1_0__11_; 
wire AES_CORE_DATAPATH_bkp_1_0__12_; 
wire AES_CORE_DATAPATH_bkp_1_0__13_; 
wire AES_CORE_DATAPATH_bkp_1_0__14_; 
wire AES_CORE_DATAPATH_bkp_1_0__15_; 
wire AES_CORE_DATAPATH_bkp_1_0__16_; 
wire AES_CORE_DATAPATH_bkp_1_0__17_; 
wire AES_CORE_DATAPATH_bkp_1_0__18_; 
wire AES_CORE_DATAPATH_bkp_1_0__19_; 
wire AES_CORE_DATAPATH_bkp_1_0__1_; 
wire AES_CORE_DATAPATH_bkp_1_0__20_; 
wire AES_CORE_DATAPATH_bkp_1_0__21_; 
wire AES_CORE_DATAPATH_bkp_1_0__22_; 
wire AES_CORE_DATAPATH_bkp_1_0__23_; 
wire AES_CORE_DATAPATH_bkp_1_0__24_; 
wire AES_CORE_DATAPATH_bkp_1_0__25_; 
wire AES_CORE_DATAPATH_bkp_1_0__26_; 
wire AES_CORE_DATAPATH_bkp_1_0__27_; 
wire AES_CORE_DATAPATH_bkp_1_0__28_; 
wire AES_CORE_DATAPATH_bkp_1_0__29_; 
wire AES_CORE_DATAPATH_bkp_1_0__2_; 
wire AES_CORE_DATAPATH_bkp_1_0__30_; 
wire AES_CORE_DATAPATH_bkp_1_0__31_; 
wire AES_CORE_DATAPATH_bkp_1_0__3_; 
wire AES_CORE_DATAPATH_bkp_1_0__4_; 
wire AES_CORE_DATAPATH_bkp_1_0__5_; 
wire AES_CORE_DATAPATH_bkp_1_0__6_; 
wire AES_CORE_DATAPATH_bkp_1_0__7_; 
wire AES_CORE_DATAPATH_bkp_1_0__8_; 
wire AES_CORE_DATAPATH_bkp_1_0__9_; 
wire AES_CORE_DATAPATH_bkp_1_1__0_; 
wire AES_CORE_DATAPATH_bkp_1_1__10_; 
wire AES_CORE_DATAPATH_bkp_1_1__11_; 
wire AES_CORE_DATAPATH_bkp_1_1__12_; 
wire AES_CORE_DATAPATH_bkp_1_1__13_; 
wire AES_CORE_DATAPATH_bkp_1_1__14_; 
wire AES_CORE_DATAPATH_bkp_1_1__15_; 
wire AES_CORE_DATAPATH_bkp_1_1__16_; 
wire AES_CORE_DATAPATH_bkp_1_1__17_; 
wire AES_CORE_DATAPATH_bkp_1_1__18_; 
wire AES_CORE_DATAPATH_bkp_1_1__19_; 
wire AES_CORE_DATAPATH_bkp_1_1__1_; 
wire AES_CORE_DATAPATH_bkp_1_1__20_; 
wire AES_CORE_DATAPATH_bkp_1_1__21_; 
wire AES_CORE_DATAPATH_bkp_1_1__22_; 
wire AES_CORE_DATAPATH_bkp_1_1__23_; 
wire AES_CORE_DATAPATH_bkp_1_1__24_; 
wire AES_CORE_DATAPATH_bkp_1_1__25_; 
wire AES_CORE_DATAPATH_bkp_1_1__26_; 
wire AES_CORE_DATAPATH_bkp_1_1__27_; 
wire AES_CORE_DATAPATH_bkp_1_1__28_; 
wire AES_CORE_DATAPATH_bkp_1_1__29_; 
wire AES_CORE_DATAPATH_bkp_1_1__2_; 
wire AES_CORE_DATAPATH_bkp_1_1__30_; 
wire AES_CORE_DATAPATH_bkp_1_1__31_; 
wire AES_CORE_DATAPATH_bkp_1_1__3_; 
wire AES_CORE_DATAPATH_bkp_1_1__4_; 
wire AES_CORE_DATAPATH_bkp_1_1__5_; 
wire AES_CORE_DATAPATH_bkp_1_1__6_; 
wire AES_CORE_DATAPATH_bkp_1_1__7_; 
wire AES_CORE_DATAPATH_bkp_1_1__8_; 
wire AES_CORE_DATAPATH_bkp_1_1__9_; 
wire AES_CORE_DATAPATH_bkp_1_2__0_; 
wire AES_CORE_DATAPATH_bkp_1_2__10_; 
wire AES_CORE_DATAPATH_bkp_1_2__11_; 
wire AES_CORE_DATAPATH_bkp_1_2__12_; 
wire AES_CORE_DATAPATH_bkp_1_2__13_; 
wire AES_CORE_DATAPATH_bkp_1_2__14_; 
wire AES_CORE_DATAPATH_bkp_1_2__15_; 
wire AES_CORE_DATAPATH_bkp_1_2__16_; 
wire AES_CORE_DATAPATH_bkp_1_2__17_; 
wire AES_CORE_DATAPATH_bkp_1_2__18_; 
wire AES_CORE_DATAPATH_bkp_1_2__19_; 
wire AES_CORE_DATAPATH_bkp_1_2__1_; 
wire AES_CORE_DATAPATH_bkp_1_2__20_; 
wire AES_CORE_DATAPATH_bkp_1_2__21_; 
wire AES_CORE_DATAPATH_bkp_1_2__22_; 
wire AES_CORE_DATAPATH_bkp_1_2__23_; 
wire AES_CORE_DATAPATH_bkp_1_2__24_; 
wire AES_CORE_DATAPATH_bkp_1_2__25_; 
wire AES_CORE_DATAPATH_bkp_1_2__26_; 
wire AES_CORE_DATAPATH_bkp_1_2__27_; 
wire AES_CORE_DATAPATH_bkp_1_2__28_; 
wire AES_CORE_DATAPATH_bkp_1_2__29_; 
wire AES_CORE_DATAPATH_bkp_1_2__2_; 
wire AES_CORE_DATAPATH_bkp_1_2__30_; 
wire AES_CORE_DATAPATH_bkp_1_2__31_; 
wire AES_CORE_DATAPATH_bkp_1_2__3_; 
wire AES_CORE_DATAPATH_bkp_1_2__4_; 
wire AES_CORE_DATAPATH_bkp_1_2__5_; 
wire AES_CORE_DATAPATH_bkp_1_2__6_; 
wire AES_CORE_DATAPATH_bkp_1_2__7_; 
wire AES_CORE_DATAPATH_bkp_1_2__8_; 
wire AES_CORE_DATAPATH_bkp_1_2__9_; 
wire AES_CORE_DATAPATH_bkp_1_3__0_; 
wire AES_CORE_DATAPATH_bkp_1_3__10_; 
wire AES_CORE_DATAPATH_bkp_1_3__11_; 
wire AES_CORE_DATAPATH_bkp_1_3__12_; 
wire AES_CORE_DATAPATH_bkp_1_3__13_; 
wire AES_CORE_DATAPATH_bkp_1_3__14_; 
wire AES_CORE_DATAPATH_bkp_1_3__15_; 
wire AES_CORE_DATAPATH_bkp_1_3__16_; 
wire AES_CORE_DATAPATH_bkp_1_3__17_; 
wire AES_CORE_DATAPATH_bkp_1_3__18_; 
wire AES_CORE_DATAPATH_bkp_1_3__19_; 
wire AES_CORE_DATAPATH_bkp_1_3__1_; 
wire AES_CORE_DATAPATH_bkp_1_3__20_; 
wire AES_CORE_DATAPATH_bkp_1_3__21_; 
wire AES_CORE_DATAPATH_bkp_1_3__22_; 
wire AES_CORE_DATAPATH_bkp_1_3__23_; 
wire AES_CORE_DATAPATH_bkp_1_3__24_; 
wire AES_CORE_DATAPATH_bkp_1_3__25_; 
wire AES_CORE_DATAPATH_bkp_1_3__26_; 
wire AES_CORE_DATAPATH_bkp_1_3__27_; 
wire AES_CORE_DATAPATH_bkp_1_3__28_; 
wire AES_CORE_DATAPATH_bkp_1_3__29_; 
wire AES_CORE_DATAPATH_bkp_1_3__2_; 
wire AES_CORE_DATAPATH_bkp_1_3__30_; 
wire AES_CORE_DATAPATH_bkp_1_3__31_; 
wire AES_CORE_DATAPATH_bkp_1_3__3_; 
wire AES_CORE_DATAPATH_bkp_1_3__4_; 
wire AES_CORE_DATAPATH_bkp_1_3__5_; 
wire AES_CORE_DATAPATH_bkp_1_3__6_; 
wire AES_CORE_DATAPATH_bkp_1_3__7_; 
wire AES_CORE_DATAPATH_bkp_1_3__8_; 
wire AES_CORE_DATAPATH_bkp_1_3__9_; 
wire AES_CORE_DATAPATH_bkp_1__0_; 
wire AES_CORE_DATAPATH_bkp_1__10_; 
wire AES_CORE_DATAPATH_bkp_1__11_; 
wire AES_CORE_DATAPATH_bkp_1__12_; 
wire AES_CORE_DATAPATH_bkp_1__13_; 
wire AES_CORE_DATAPATH_bkp_1__14_; 
wire AES_CORE_DATAPATH_bkp_1__15_; 
wire AES_CORE_DATAPATH_bkp_1__16_; 
wire AES_CORE_DATAPATH_bkp_1__17_; 
wire AES_CORE_DATAPATH_bkp_1__18_; 
wire AES_CORE_DATAPATH_bkp_1__19_; 
wire AES_CORE_DATAPATH_bkp_1__1_; 
wire AES_CORE_DATAPATH_bkp_1__20_; 
wire AES_CORE_DATAPATH_bkp_1__21_; 
wire AES_CORE_DATAPATH_bkp_1__22_; 
wire AES_CORE_DATAPATH_bkp_1__23_; 
wire AES_CORE_DATAPATH_bkp_1__24_; 
wire AES_CORE_DATAPATH_bkp_1__25_; 
wire AES_CORE_DATAPATH_bkp_1__26_; 
wire AES_CORE_DATAPATH_bkp_1__27_; 
wire AES_CORE_DATAPATH_bkp_1__28_; 
wire AES_CORE_DATAPATH_bkp_1__29_; 
wire AES_CORE_DATAPATH_bkp_1__2_; 
wire AES_CORE_DATAPATH_bkp_1__30_; 
wire AES_CORE_DATAPATH_bkp_1__31_; 
wire AES_CORE_DATAPATH_bkp_1__3_; 
wire AES_CORE_DATAPATH_bkp_1__4_; 
wire AES_CORE_DATAPATH_bkp_1__5_; 
wire AES_CORE_DATAPATH_bkp_1__6_; 
wire AES_CORE_DATAPATH_bkp_1__7_; 
wire AES_CORE_DATAPATH_bkp_1__8_; 
wire AES_CORE_DATAPATH_bkp_1__9_; 
wire AES_CORE_DATAPATH_bkp_2__0_; 
wire AES_CORE_DATAPATH_bkp_2__10_; 
wire AES_CORE_DATAPATH_bkp_2__11_; 
wire AES_CORE_DATAPATH_bkp_2__12_; 
wire AES_CORE_DATAPATH_bkp_2__13_; 
wire AES_CORE_DATAPATH_bkp_2__14_; 
wire AES_CORE_DATAPATH_bkp_2__15_; 
wire AES_CORE_DATAPATH_bkp_2__16_; 
wire AES_CORE_DATAPATH_bkp_2__17_; 
wire AES_CORE_DATAPATH_bkp_2__18_; 
wire AES_CORE_DATAPATH_bkp_2__19_; 
wire AES_CORE_DATAPATH_bkp_2__1_; 
wire AES_CORE_DATAPATH_bkp_2__20_; 
wire AES_CORE_DATAPATH_bkp_2__21_; 
wire AES_CORE_DATAPATH_bkp_2__22_; 
wire AES_CORE_DATAPATH_bkp_2__23_; 
wire AES_CORE_DATAPATH_bkp_2__24_; 
wire AES_CORE_DATAPATH_bkp_2__25_; 
wire AES_CORE_DATAPATH_bkp_2__26_; 
wire AES_CORE_DATAPATH_bkp_2__27_; 
wire AES_CORE_DATAPATH_bkp_2__28_; 
wire AES_CORE_DATAPATH_bkp_2__29_; 
wire AES_CORE_DATAPATH_bkp_2__2_; 
wire AES_CORE_DATAPATH_bkp_2__30_; 
wire AES_CORE_DATAPATH_bkp_2__31_; 
wire AES_CORE_DATAPATH_bkp_2__3_; 
wire AES_CORE_DATAPATH_bkp_2__4_; 
wire AES_CORE_DATAPATH_bkp_2__5_; 
wire AES_CORE_DATAPATH_bkp_2__6_; 
wire AES_CORE_DATAPATH_bkp_2__7_; 
wire AES_CORE_DATAPATH_bkp_2__8_; 
wire AES_CORE_DATAPATH_bkp_2__9_; 
wire AES_CORE_DATAPATH_bkp_3__0_; 
wire AES_CORE_DATAPATH_bkp_3__10_; 
wire AES_CORE_DATAPATH_bkp_3__11_; 
wire AES_CORE_DATAPATH_bkp_3__12_; 
wire AES_CORE_DATAPATH_bkp_3__13_; 
wire AES_CORE_DATAPATH_bkp_3__14_; 
wire AES_CORE_DATAPATH_bkp_3__15_; 
wire AES_CORE_DATAPATH_bkp_3__16_; 
wire AES_CORE_DATAPATH_bkp_3__17_; 
wire AES_CORE_DATAPATH_bkp_3__18_; 
wire AES_CORE_DATAPATH_bkp_3__19_; 
wire AES_CORE_DATAPATH_bkp_3__1_; 
wire AES_CORE_DATAPATH_bkp_3__20_; 
wire AES_CORE_DATAPATH_bkp_3__21_; 
wire AES_CORE_DATAPATH_bkp_3__22_; 
wire AES_CORE_DATAPATH_bkp_3__23_; 
wire AES_CORE_DATAPATH_bkp_3__24_; 
wire AES_CORE_DATAPATH_bkp_3__25_; 
wire AES_CORE_DATAPATH_bkp_3__26_; 
wire AES_CORE_DATAPATH_bkp_3__27_; 
wire AES_CORE_DATAPATH_bkp_3__28_; 
wire AES_CORE_DATAPATH_bkp_3__29_; 
wire AES_CORE_DATAPATH_bkp_3__2_; 
wire AES_CORE_DATAPATH_bkp_3__30_; 
wire AES_CORE_DATAPATH_bkp_3__31_; 
wire AES_CORE_DATAPATH_bkp_3__3_; 
wire AES_CORE_DATAPATH_bkp_3__4_; 
wire AES_CORE_DATAPATH_bkp_3__5_; 
wire AES_CORE_DATAPATH_bkp_3__6_; 
wire AES_CORE_DATAPATH_bkp_3__7_; 
wire AES_CORE_DATAPATH_bkp_3__8_; 
wire AES_CORE_DATAPATH_bkp_3__9_; 
wire AES_CORE_DATAPATH_col_0__0_; 
wire AES_CORE_DATAPATH_col_0__10_; 
wire AES_CORE_DATAPATH_col_0__11_; 
wire AES_CORE_DATAPATH_col_0__12_; 
wire AES_CORE_DATAPATH_col_0__13_; 
wire AES_CORE_DATAPATH_col_0__14_; 
wire AES_CORE_DATAPATH_col_0__15_; 
wire AES_CORE_DATAPATH_col_0__16_; 
wire AES_CORE_DATAPATH_col_0__17_; 
wire AES_CORE_DATAPATH_col_0__18_; 
wire AES_CORE_DATAPATH_col_0__19_; 
wire AES_CORE_DATAPATH_col_0__1_; 
wire AES_CORE_DATAPATH_col_0__20_; 
wire AES_CORE_DATAPATH_col_0__21_; 
wire AES_CORE_DATAPATH_col_0__22_; 
wire AES_CORE_DATAPATH_col_0__23_; 
wire AES_CORE_DATAPATH_col_0__24_; 
wire AES_CORE_DATAPATH_col_0__25_; 
wire AES_CORE_DATAPATH_col_0__26_; 
wire AES_CORE_DATAPATH_col_0__27_; 
wire AES_CORE_DATAPATH_col_0__28_; 
wire AES_CORE_DATAPATH_col_0__29_; 
wire AES_CORE_DATAPATH_col_0__2_; 
wire AES_CORE_DATAPATH_col_0__30_; 
wire AES_CORE_DATAPATH_col_0__31_; 
wire AES_CORE_DATAPATH_col_0__3_; 
wire AES_CORE_DATAPATH_col_0__4_; 
wire AES_CORE_DATAPATH_col_0__5_; 
wire AES_CORE_DATAPATH_col_0__6_; 
wire AES_CORE_DATAPATH_col_0__7_; 
wire AES_CORE_DATAPATH_col_0__8_; 
wire AES_CORE_DATAPATH_col_0__9_; 
wire AES_CORE_DATAPATH_col_3__0_; 
wire AES_CORE_DATAPATH_col_3__10_; 
wire AES_CORE_DATAPATH_col_3__11_; 
wire AES_CORE_DATAPATH_col_3__12_; 
wire AES_CORE_DATAPATH_col_3__13_; 
wire AES_CORE_DATAPATH_col_3__14_; 
wire AES_CORE_DATAPATH_col_3__15_; 
wire AES_CORE_DATAPATH_col_3__16_; 
wire AES_CORE_DATAPATH_col_3__17_; 
wire AES_CORE_DATAPATH_col_3__18_; 
wire AES_CORE_DATAPATH_col_3__19_; 
wire AES_CORE_DATAPATH_col_3__1_; 
wire AES_CORE_DATAPATH_col_3__20_; 
wire AES_CORE_DATAPATH_col_3__21_; 
wire AES_CORE_DATAPATH_col_3__22_; 
wire AES_CORE_DATAPATH_col_3__23_; 
wire AES_CORE_DATAPATH_col_3__24_; 
wire AES_CORE_DATAPATH_col_3__25_; 
wire AES_CORE_DATAPATH_col_3__26_; 
wire AES_CORE_DATAPATH_col_3__27_; 
wire AES_CORE_DATAPATH_col_3__28_; 
wire AES_CORE_DATAPATH_col_3__29_; 
wire AES_CORE_DATAPATH_col_3__2_; 
wire AES_CORE_DATAPATH_col_3__30_; 
wire AES_CORE_DATAPATH_col_3__31_; 
wire AES_CORE_DATAPATH_col_3__3_; 
wire AES_CORE_DATAPATH_col_3__4_; 
wire AES_CORE_DATAPATH_col_3__5_; 
wire AES_CORE_DATAPATH_col_3__6_; 
wire AES_CORE_DATAPATH_col_3__7_; 
wire AES_CORE_DATAPATH_col_3__8_; 
wire AES_CORE_DATAPATH_col_3__9_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_; 
wire AES_CORE_DATAPATH_col_en_host_0_; 
wire AES_CORE_DATAPATH_col_en_host_1_; 
wire AES_CORE_DATAPATH_col_en_host_2_; 
wire AES_CORE_DATAPATH_col_en_host_3_; 
wire AES_CORE_DATAPATH_col_sel_host_0_; 
wire AES_CORE_DATAPATH_col_sel_host_1_; 
wire AES_CORE_DATAPATH_col_sel_pp1_0_; 
wire AES_CORE_DATAPATH_col_sel_pp1_1_; 
wire AES_CORE_DATAPATH_col_sel_pp2_0_; 
wire AES_CORE_DATAPATH_col_sel_pp2_1_; 
wire AES_CORE_DATAPATH_iv_0__0_; 
wire AES_CORE_DATAPATH_iv_0__10_; 
wire AES_CORE_DATAPATH_iv_0__11_; 
wire AES_CORE_DATAPATH_iv_0__12_; 
wire AES_CORE_DATAPATH_iv_0__13_; 
wire AES_CORE_DATAPATH_iv_0__14_; 
wire AES_CORE_DATAPATH_iv_0__15_; 
wire AES_CORE_DATAPATH_iv_0__16_; 
wire AES_CORE_DATAPATH_iv_0__17_; 
wire AES_CORE_DATAPATH_iv_0__18_; 
wire AES_CORE_DATAPATH_iv_0__19_; 
wire AES_CORE_DATAPATH_iv_0__1_; 
wire AES_CORE_DATAPATH_iv_0__20_; 
wire AES_CORE_DATAPATH_iv_0__21_; 
wire AES_CORE_DATAPATH_iv_0__22_; 
wire AES_CORE_DATAPATH_iv_0__23_; 
wire AES_CORE_DATAPATH_iv_0__24_; 
wire AES_CORE_DATAPATH_iv_0__25_; 
wire AES_CORE_DATAPATH_iv_0__26_; 
wire AES_CORE_DATAPATH_iv_0__27_; 
wire AES_CORE_DATAPATH_iv_0__28_; 
wire AES_CORE_DATAPATH_iv_0__29_; 
wire AES_CORE_DATAPATH_iv_0__2_; 
wire AES_CORE_DATAPATH_iv_0__30_; 
wire AES_CORE_DATAPATH_iv_0__31_; 
wire AES_CORE_DATAPATH_iv_0__3_; 
wire AES_CORE_DATAPATH_iv_0__4_; 
wire AES_CORE_DATAPATH_iv_0__5_; 
wire AES_CORE_DATAPATH_iv_0__6_; 
wire AES_CORE_DATAPATH_iv_0__7_; 
wire AES_CORE_DATAPATH_iv_0__8_; 
wire AES_CORE_DATAPATH_iv_0__9_; 
wire AES_CORE_DATAPATH_iv_1__0_; 
wire AES_CORE_DATAPATH_iv_1__10_; 
wire AES_CORE_DATAPATH_iv_1__11_; 
wire AES_CORE_DATAPATH_iv_1__12_; 
wire AES_CORE_DATAPATH_iv_1__13_; 
wire AES_CORE_DATAPATH_iv_1__14_; 
wire AES_CORE_DATAPATH_iv_1__15_; 
wire AES_CORE_DATAPATH_iv_1__16_; 
wire AES_CORE_DATAPATH_iv_1__17_; 
wire AES_CORE_DATAPATH_iv_1__18_; 
wire AES_CORE_DATAPATH_iv_1__19_; 
wire AES_CORE_DATAPATH_iv_1__1_; 
wire AES_CORE_DATAPATH_iv_1__20_; 
wire AES_CORE_DATAPATH_iv_1__21_; 
wire AES_CORE_DATAPATH_iv_1__22_; 
wire AES_CORE_DATAPATH_iv_1__23_; 
wire AES_CORE_DATAPATH_iv_1__24_; 
wire AES_CORE_DATAPATH_iv_1__25_; 
wire AES_CORE_DATAPATH_iv_1__26_; 
wire AES_CORE_DATAPATH_iv_1__27_; 
wire AES_CORE_DATAPATH_iv_1__28_; 
wire AES_CORE_DATAPATH_iv_1__29_; 
wire AES_CORE_DATAPATH_iv_1__2_; 
wire AES_CORE_DATAPATH_iv_1__30_; 
wire AES_CORE_DATAPATH_iv_1__31_; 
wire AES_CORE_DATAPATH_iv_1__3_; 
wire AES_CORE_DATAPATH_iv_1__4_; 
wire AES_CORE_DATAPATH_iv_1__5_; 
wire AES_CORE_DATAPATH_iv_1__6_; 
wire AES_CORE_DATAPATH_iv_1__7_; 
wire AES_CORE_DATAPATH_iv_1__8_; 
wire AES_CORE_DATAPATH_iv_1__9_; 
wire AES_CORE_DATAPATH_iv_2__0_; 
wire AES_CORE_DATAPATH_iv_2__10_; 
wire AES_CORE_DATAPATH_iv_2__11_; 
wire AES_CORE_DATAPATH_iv_2__12_; 
wire AES_CORE_DATAPATH_iv_2__13_; 
wire AES_CORE_DATAPATH_iv_2__14_; 
wire AES_CORE_DATAPATH_iv_2__15_; 
wire AES_CORE_DATAPATH_iv_2__16_; 
wire AES_CORE_DATAPATH_iv_2__17_; 
wire AES_CORE_DATAPATH_iv_2__18_; 
wire AES_CORE_DATAPATH_iv_2__19_; 
wire AES_CORE_DATAPATH_iv_2__1_; 
wire AES_CORE_DATAPATH_iv_2__20_; 
wire AES_CORE_DATAPATH_iv_2__21_; 
wire AES_CORE_DATAPATH_iv_2__22_; 
wire AES_CORE_DATAPATH_iv_2__23_; 
wire AES_CORE_DATAPATH_iv_2__24_; 
wire AES_CORE_DATAPATH_iv_2__25_; 
wire AES_CORE_DATAPATH_iv_2__26_; 
wire AES_CORE_DATAPATH_iv_2__27_; 
wire AES_CORE_DATAPATH_iv_2__28_; 
wire AES_CORE_DATAPATH_iv_2__29_; 
wire AES_CORE_DATAPATH_iv_2__2_; 
wire AES_CORE_DATAPATH_iv_2__30_; 
wire AES_CORE_DATAPATH_iv_2__31_; 
wire AES_CORE_DATAPATH_iv_2__3_; 
wire AES_CORE_DATAPATH_iv_2__4_; 
wire AES_CORE_DATAPATH_iv_2__5_; 
wire AES_CORE_DATAPATH_iv_2__6_; 
wire AES_CORE_DATAPATH_iv_2__7_; 
wire AES_CORE_DATAPATH_iv_2__8_; 
wire AES_CORE_DATAPATH_iv_2__9_; 
wire AES_CORE_DATAPATH_iv_3__0_; 
wire AES_CORE_DATAPATH_iv_3__10_; 
wire AES_CORE_DATAPATH_iv_3__11_; 
wire AES_CORE_DATAPATH_iv_3__12_; 
wire AES_CORE_DATAPATH_iv_3__13_; 
wire AES_CORE_DATAPATH_iv_3__14_; 
wire AES_CORE_DATAPATH_iv_3__15_; 
wire AES_CORE_DATAPATH_iv_3__16_; 
wire AES_CORE_DATAPATH_iv_3__17_; 
wire AES_CORE_DATAPATH_iv_3__18_; 
wire AES_CORE_DATAPATH_iv_3__19_; 
wire AES_CORE_DATAPATH_iv_3__1_; 
wire AES_CORE_DATAPATH_iv_3__20_; 
wire AES_CORE_DATAPATH_iv_3__21_; 
wire AES_CORE_DATAPATH_iv_3__22_; 
wire AES_CORE_DATAPATH_iv_3__23_; 
wire AES_CORE_DATAPATH_iv_3__24_; 
wire AES_CORE_DATAPATH_iv_3__25_; 
wire AES_CORE_DATAPATH_iv_3__26_; 
wire AES_CORE_DATAPATH_iv_3__27_; 
wire AES_CORE_DATAPATH_iv_3__28_; 
wire AES_CORE_DATAPATH_iv_3__29_; 
wire AES_CORE_DATAPATH_iv_3__2_; 
wire AES_CORE_DATAPATH_iv_3__30_; 
wire AES_CORE_DATAPATH_iv_3__31_; 
wire AES_CORE_DATAPATH_iv_3__3_; 
wire AES_CORE_DATAPATH_iv_3__4_; 
wire AES_CORE_DATAPATH_iv_3__5_; 
wire AES_CORE_DATAPATH_iv_3__6_; 
wire AES_CORE_DATAPATH_iv_3__7_; 
wire AES_CORE_DATAPATH_iv_3__8_; 
wire AES_CORE_DATAPATH_iv_3__9_; 
wire AES_CORE_DATAPATH_key_en_pp1_0_; 
wire AES_CORE_DATAPATH_key_en_pp1_1_; 
wire AES_CORE_DATAPATH_key_en_pp1_2_; 
wire AES_CORE_DATAPATH_key_en_pp1_3_; 
wire AES_CORE_DATAPATH_key_host_0__0_; 
wire AES_CORE_DATAPATH_key_host_0__10_; 
wire AES_CORE_DATAPATH_key_host_0__11_; 
wire AES_CORE_DATAPATH_key_host_0__12_; 
wire AES_CORE_DATAPATH_key_host_0__13_; 
wire AES_CORE_DATAPATH_key_host_0__14_; 
wire AES_CORE_DATAPATH_key_host_0__15_; 
wire AES_CORE_DATAPATH_key_host_0__16_; 
wire AES_CORE_DATAPATH_key_host_0__17_; 
wire AES_CORE_DATAPATH_key_host_0__18_; 
wire AES_CORE_DATAPATH_key_host_0__19_; 
wire AES_CORE_DATAPATH_key_host_0__1_; 
wire AES_CORE_DATAPATH_key_host_0__20_; 
wire AES_CORE_DATAPATH_key_host_0__21_; 
wire AES_CORE_DATAPATH_key_host_0__22_; 
wire AES_CORE_DATAPATH_key_host_0__23_; 
wire AES_CORE_DATAPATH_key_host_0__24_; 
wire AES_CORE_DATAPATH_key_host_0__25_; 
wire AES_CORE_DATAPATH_key_host_0__26_; 
wire AES_CORE_DATAPATH_key_host_0__27_; 
wire AES_CORE_DATAPATH_key_host_0__28_; 
wire AES_CORE_DATAPATH_key_host_0__29_; 
wire AES_CORE_DATAPATH_key_host_0__2_; 
wire AES_CORE_DATAPATH_key_host_0__30_; 
wire AES_CORE_DATAPATH_key_host_0__31_; 
wire AES_CORE_DATAPATH_key_host_0__3_; 
wire AES_CORE_DATAPATH_key_host_0__4_; 
wire AES_CORE_DATAPATH_key_host_0__5_; 
wire AES_CORE_DATAPATH_key_host_0__6_; 
wire AES_CORE_DATAPATH_key_host_0__7_; 
wire AES_CORE_DATAPATH_key_host_0__8_; 
wire AES_CORE_DATAPATH_key_host_0__9_; 
wire AES_CORE_DATAPATH_key_host_1__0_; 
wire AES_CORE_DATAPATH_key_host_1__10_; 
wire AES_CORE_DATAPATH_key_host_1__11_; 
wire AES_CORE_DATAPATH_key_host_1__12_; 
wire AES_CORE_DATAPATH_key_host_1__13_; 
wire AES_CORE_DATAPATH_key_host_1__14_; 
wire AES_CORE_DATAPATH_key_host_1__15_; 
wire AES_CORE_DATAPATH_key_host_1__16_; 
wire AES_CORE_DATAPATH_key_host_1__17_; 
wire AES_CORE_DATAPATH_key_host_1__18_; 
wire AES_CORE_DATAPATH_key_host_1__19_; 
wire AES_CORE_DATAPATH_key_host_1__1_; 
wire AES_CORE_DATAPATH_key_host_1__20_; 
wire AES_CORE_DATAPATH_key_host_1__21_; 
wire AES_CORE_DATAPATH_key_host_1__22_; 
wire AES_CORE_DATAPATH_key_host_1__23_; 
wire AES_CORE_DATAPATH_key_host_1__24_; 
wire AES_CORE_DATAPATH_key_host_1__25_; 
wire AES_CORE_DATAPATH_key_host_1__26_; 
wire AES_CORE_DATAPATH_key_host_1__27_; 
wire AES_CORE_DATAPATH_key_host_1__28_; 
wire AES_CORE_DATAPATH_key_host_1__29_; 
wire AES_CORE_DATAPATH_key_host_1__2_; 
wire AES_CORE_DATAPATH_key_host_1__30_; 
wire AES_CORE_DATAPATH_key_host_1__31_; 
wire AES_CORE_DATAPATH_key_host_1__3_; 
wire AES_CORE_DATAPATH_key_host_1__4_; 
wire AES_CORE_DATAPATH_key_host_1__5_; 
wire AES_CORE_DATAPATH_key_host_1__6_; 
wire AES_CORE_DATAPATH_key_host_1__7_; 
wire AES_CORE_DATAPATH_key_host_1__8_; 
wire AES_CORE_DATAPATH_key_host_1__9_; 
wire AES_CORE_DATAPATH_key_host_2__0_; 
wire AES_CORE_DATAPATH_key_host_2__10_; 
wire AES_CORE_DATAPATH_key_host_2__11_; 
wire AES_CORE_DATAPATH_key_host_2__12_; 
wire AES_CORE_DATAPATH_key_host_2__13_; 
wire AES_CORE_DATAPATH_key_host_2__14_; 
wire AES_CORE_DATAPATH_key_host_2__15_; 
wire AES_CORE_DATAPATH_key_host_2__16_; 
wire AES_CORE_DATAPATH_key_host_2__17_; 
wire AES_CORE_DATAPATH_key_host_2__18_; 
wire AES_CORE_DATAPATH_key_host_2__19_; 
wire AES_CORE_DATAPATH_key_host_2__1_; 
wire AES_CORE_DATAPATH_key_host_2__20_; 
wire AES_CORE_DATAPATH_key_host_2__21_; 
wire AES_CORE_DATAPATH_key_host_2__22_; 
wire AES_CORE_DATAPATH_key_host_2__23_; 
wire AES_CORE_DATAPATH_key_host_2__24_; 
wire AES_CORE_DATAPATH_key_host_2__25_; 
wire AES_CORE_DATAPATH_key_host_2__26_; 
wire AES_CORE_DATAPATH_key_host_2__27_; 
wire AES_CORE_DATAPATH_key_host_2__28_; 
wire AES_CORE_DATAPATH_key_host_2__29_; 
wire AES_CORE_DATAPATH_key_host_2__2_; 
wire AES_CORE_DATAPATH_key_host_2__30_; 
wire AES_CORE_DATAPATH_key_host_2__31_; 
wire AES_CORE_DATAPATH_key_host_2__3_; 
wire AES_CORE_DATAPATH_key_host_2__4_; 
wire AES_CORE_DATAPATH_key_host_2__5_; 
wire AES_CORE_DATAPATH_key_host_2__6_; 
wire AES_CORE_DATAPATH_key_host_2__7_; 
wire AES_CORE_DATAPATH_key_host_2__8_; 
wire AES_CORE_DATAPATH_key_host_2__9_; 
wire AES_CORE_DATAPATH_key_host_3__0_; 
wire AES_CORE_DATAPATH_key_host_3__10_; 
wire AES_CORE_DATAPATH_key_host_3__11_; 
wire AES_CORE_DATAPATH_key_host_3__12_; 
wire AES_CORE_DATAPATH_key_host_3__13_; 
wire AES_CORE_DATAPATH_key_host_3__14_; 
wire AES_CORE_DATAPATH_key_host_3__15_; 
wire AES_CORE_DATAPATH_key_host_3__16_; 
wire AES_CORE_DATAPATH_key_host_3__17_; 
wire AES_CORE_DATAPATH_key_host_3__18_; 
wire AES_CORE_DATAPATH_key_host_3__19_; 
wire AES_CORE_DATAPATH_key_host_3__1_; 
wire AES_CORE_DATAPATH_key_host_3__20_; 
wire AES_CORE_DATAPATH_key_host_3__21_; 
wire AES_CORE_DATAPATH_key_host_3__22_; 
wire AES_CORE_DATAPATH_key_host_3__23_; 
wire AES_CORE_DATAPATH_key_host_3__24_; 
wire AES_CORE_DATAPATH_key_host_3__25_; 
wire AES_CORE_DATAPATH_key_host_3__26_; 
wire AES_CORE_DATAPATH_key_host_3__27_; 
wire AES_CORE_DATAPATH_key_host_3__28_; 
wire AES_CORE_DATAPATH_key_host_3__29_; 
wire AES_CORE_DATAPATH_key_host_3__2_; 
wire AES_CORE_DATAPATH_key_host_3__30_; 
wire AES_CORE_DATAPATH_key_host_3__31_; 
wire AES_CORE_DATAPATH_key_host_3__3_; 
wire AES_CORE_DATAPATH_key_host_3__4_; 
wire AES_CORE_DATAPATH_key_host_3__5_; 
wire AES_CORE_DATAPATH_key_host_3__6_; 
wire AES_CORE_DATAPATH_key_host_3__7_; 
wire AES_CORE_DATAPATH_key_host_3__8_; 
wire AES_CORE_DATAPATH_key_host_3__9_; 
wire AES_CORE_DATAPATH_key_out_sel_pp1_0_; 
wire AES_CORE_DATAPATH_key_out_sel_pp1_1_; 
wire AES_CORE_DATAPATH_key_out_sel_pp2_0_; 
wire AES_CORE_DATAPATH_key_out_sel_pp2_1_; 
wire AES_CORE_DATAPATH_key_sel_pp1; 
wire AES_CORE_DATAPATH_last_round_pp1; 
wire AES_CORE_DATAPATH_last_round_pp2; 
wire AES_CORE_DATAPATH_rk_out_sel; 
wire AES_CORE_DATAPATH_rk_out_sel_pp1; 
wire AES_CORE_DATAPATH_rk_out_sel_pp2; 
wire AES_CORE_DATAPATH_rk_sel_pp1_0_; 
wire AES_CORE_DATAPATH_rk_sel_pp1_1_; 
wire AES_CORE_DATAPATH_rk_sel_pp2_0_; 
wire AES_CORE_DATAPATH_rk_sel_pp2_1_; 
wire _abc_15574_new_n11_; 
wire _abc_15574_new_n13_; 
wire _abc_15574_new_n15_; 
wire _abc_15574_new_n17_; 
input \addr[0] ;
input \addr[1] ;
input \aes_mode[0] ;
input \aes_mode[1] ;
input \bus_in[0] ;
input \bus_in[10] ;
input \bus_in[11] ;
input \bus_in[12] ;
input \bus_in[13] ;
input \bus_in[14] ;
input \bus_in[15] ;
input \bus_in[16] ;
input \bus_in[17] ;
input \bus_in[18] ;
input \bus_in[19] ;
input \bus_in[1] ;
input \bus_in[20] ;
input \bus_in[21] ;
input \bus_in[22] ;
input \bus_in[23] ;
input \bus_in[24] ;
input \bus_in[25] ;
input \bus_in[26] ;
input \bus_in[27] ;
input \bus_in[28] ;
input \bus_in[29] ;
input \bus_in[2] ;
input \bus_in[30] ;
input \bus_in[31] ;
input \bus_in[3] ;
input \bus_in[4] ;
input \bus_in[5] ;
input \bus_in[6] ;
input \bus_in[7] ;
input \bus_in[8] ;
input \bus_in[9] ;
input clk;
output \col_out[0] ;
output \col_out[10] ;
output \col_out[11] ;
output \col_out[12] ;
output \col_out[13] ;
output \col_out[14] ;
output \col_out[15] ;
output \col_out[16] ;
output \col_out[17] ;
output \col_out[18] ;
output \col_out[19] ;
output \col_out[1] ;
output \col_out[20] ;
output \col_out[21] ;
output \col_out[22] ;
output \col_out[23] ;
output \col_out[24] ;
output \col_out[25] ;
output \col_out[26] ;
output \col_out[27] ;
output \col_out[28] ;
output \col_out[29] ;
output \col_out[2] ;
output \col_out[30] ;
output \col_out[31] ;
output \col_out[3] ;
output \col_out[4] ;
output \col_out[5] ;
output \col_out[6] ;
output \col_out[7] ;
output \col_out[8] ;
output \col_out[9] ;
input \data_type[0] ;
input \data_type[1] ;
input disable_core;
output end_aes;
input first_block;
input \iv_en[0] ;
input \iv_en[1] ;
input \iv_en[2] ;
input \iv_en[3] ;
output \iv_out[0] ;
output \iv_out[10] ;
output \iv_out[11] ;
output \iv_out[12] ;
output \iv_out[13] ;
output \iv_out[14] ;
output \iv_out[15] ;
output \iv_out[16] ;
output \iv_out[17] ;
output \iv_out[18] ;
output \iv_out[19] ;
output \iv_out[1] ;
output \iv_out[20] ;
output \iv_out[21] ;
output \iv_out[22] ;
output \iv_out[23] ;
output \iv_out[24] ;
output \iv_out[25] ;
output \iv_out[26] ;
output \iv_out[27] ;
output \iv_out[28] ;
output \iv_out[29] ;
output \iv_out[2] ;
output \iv_out[30] ;
output \iv_out[31] ;
output \iv_out[3] ;
output \iv_out[4] ;
output \iv_out[5] ;
output \iv_out[6] ;
output \iv_out[7] ;
output \iv_out[8] ;
output \iv_out[9] ;
input \iv_sel_rd[0] ;
input \iv_sel_rd[1] ;
input \iv_sel_rd[2] ;
input \iv_sel_rd[3] ;
input \key_en[0] ;
input \key_en[1] ;
input \key_en[2] ;
input \key_en[3] ;
output \key_out[0] ;
output \key_out[10] ;
output \key_out[11] ;
output \key_out[12] ;
output \key_out[13] ;
output \key_out[14] ;
output \key_out[15] ;
output \key_out[16] ;
output \key_out[17] ;
output \key_out[18] ;
output \key_out[19] ;
output \key_out[1] ;
output \key_out[20] ;
output \key_out[21] ;
output \key_out[22] ;
output \key_out[23] ;
output \key_out[24] ;
output \key_out[25] ;
output \key_out[26] ;
output \key_out[27] ;
output \key_out[28] ;
output \key_out[29] ;
output \key_out[2] ;
output \key_out[30] ;
output \key_out[31] ;
output \key_out[3] ;
output \key_out[4] ;
output \key_out[5] ;
output \key_out[6] ;
output \key_out[7] ;
output \key_out[8] ;
output \key_out[9] ;
input \key_sel_rd[0] ;
input \key_sel_rd[1] ;
input \op_mode[0] ;
input \op_mode[1] ;
input read_en;
input rst_n;
input start;
input write_en;
AND2X2 AND2X2_1 ( .A(\addr[0] ), .B(read_en), .Y(AES_CORE_DATAPATH_col_sel_host_0_));
AND2X2 AND2X2_10 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .B(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1817));
AND2X2 AND2X2_100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n138_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n214_));
AND2X2 AND2X2_101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n218_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n219_));
AND2X2 AND2X2_102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n209_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n211_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n226_));
AND2X2 AND2X2_103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n261_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n266_));
AND2X2 AND2X2_104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n398_));
AND2X2 AND2X2_105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_));
AND2X2 AND2X2_106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n415_));
AND2X2 AND2X2_107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n419_));
AND2X2 AND2X2_108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n52_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n57_));
AND2X2 AND2X2_109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n145_));
AND2X2 AND2X2_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2459_), .B(AES_CORE_DATAPATH__abc_15863_new_n2460_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2461_));
AND2X2 AND2X2_110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n138_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n214_));
AND2X2 AND2X2_111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n218_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n219_));
AND2X2 AND2X2_112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n209_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n211_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n226_));
AND2X2 AND2X2_113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n261_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n266_));
AND2X2 AND2X2_114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n398_));
AND2X2 AND2X2_115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_));
AND2X2 AND2X2_116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n415_));
AND2X2 AND2X2_117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n419_));
AND2X2 AND2X2_118 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_));
AND2X2 AND2X2_119 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_));
AND2X2 AND2X2_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2726_), .B(AES_CORE_DATAPATH__abc_15863_new_n2727_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2737_));
AND2X2 AND2X2_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3098_), .B(AES_CORE_DATAPATH__abc_15863_new_n3076_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3099_));
AND2X2 AND2X2_14 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3097_), .B(AES_CORE_DATAPATH__abc_15863_new_n3101_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3102_));
AND2X2 AND2X2_15 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3124_), .B(AES_CORE_DATAPATH__abc_15863_new_n3125_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3126_));
AND2X2 AND2X2_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3146_), .B(AES_CORE_DATAPATH__abc_15863_new_n3147_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3148_));
AND2X2 AND2X2_17 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3169_), .B(AES_CORE_DATAPATH__abc_15863_new_n3170_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3171_));
AND2X2 AND2X2_18 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3191_), .B(AES_CORE_DATAPATH__abc_15863_new_n3192_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3193_));
AND2X2 AND2X2_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3213_), .B(AES_CORE_DATAPATH__abc_15863_new_n3214_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3215_));
AND2X2 AND2X2_2 ( .A(\addr[1] ), .B(read_en), .Y(AES_CORE_DATAPATH_col_sel_host_1_));
AND2X2 AND2X2_20 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3235_), .B(AES_CORE_DATAPATH__abc_15863_new_n3236_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3237_));
AND2X2 AND2X2_21 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3257_), .B(AES_CORE_DATAPATH__abc_15863_new_n3258_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3259_));
AND2X2 AND2X2_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3279_), .B(AES_CORE_DATAPATH__abc_15863_new_n3280_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3281_));
AND2X2 AND2X2_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3301_), .B(AES_CORE_DATAPATH__abc_15863_new_n3302_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3303_));
AND2X2 AND2X2_24 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3323_), .B(AES_CORE_DATAPATH__abc_15863_new_n3324_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3325_));
AND2X2 AND2X2_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3345_), .B(AES_CORE_DATAPATH__abc_15863_new_n3346_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3347_));
AND2X2 AND2X2_26 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3367_), .B(AES_CORE_DATAPATH__abc_15863_new_n3368_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3369_));
AND2X2 AND2X2_27 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3389_), .B(AES_CORE_DATAPATH__abc_15863_new_n3390_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3391_));
AND2X2 AND2X2_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3411_), .B(AES_CORE_DATAPATH__abc_15863_new_n3412_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3413_));
AND2X2 AND2X2_29 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3433_), .B(AES_CORE_DATAPATH__abc_15863_new_n3434_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3435_));
AND2X2 AND2X2_3 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n78_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n79_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n80_));
AND2X2 AND2X2_30 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3455_), .B(AES_CORE_DATAPATH__abc_15863_new_n3456_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3457_));
AND2X2 AND2X2_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3477_), .B(AES_CORE_DATAPATH__abc_15863_new_n3478_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3479_));
AND2X2 AND2X2_32 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3499_), .B(AES_CORE_DATAPATH__abc_15863_new_n3500_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3503_));
AND2X2 AND2X2_33 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3521_), .B(AES_CORE_DATAPATH__abc_15863_new_n3522_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3523_));
AND2X2 AND2X2_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3543_), .B(AES_CORE_DATAPATH__abc_15863_new_n3544_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3545_));
AND2X2 AND2X2_35 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3565_), .B(AES_CORE_DATAPATH__abc_15863_new_n3566_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3567_));
AND2X2 AND2X2_36 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3587_), .B(AES_CORE_DATAPATH__abc_15863_new_n3588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3589_));
AND2X2 AND2X2_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3609_), .B(AES_CORE_DATAPATH__abc_15863_new_n3610_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3611_));
AND2X2 AND2X2_38 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3631_), .B(AES_CORE_DATAPATH__abc_15863_new_n3632_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3633_));
AND2X2 AND2X2_39 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3653_), .B(AES_CORE_DATAPATH__abc_15863_new_n3654_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3655_));
AND2X2 AND2X2_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n114_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n115_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n116_));
AND2X2 AND2X2_40 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3675_), .B(AES_CORE_DATAPATH__abc_15863_new_n3676_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3679_));
AND2X2 AND2X2_41 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3697_), .B(AES_CORE_DATAPATH__abc_15863_new_n3698_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3699_));
AND2X2 AND2X2_42 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3719_), .B(AES_CORE_DATAPATH__abc_15863_new_n3720_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3721_));
AND2X2 AND2X2_43 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3741_), .B(AES_CORE_DATAPATH__abc_15863_new_n3742_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3743_));
AND2X2 AND2X2_44 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3763_), .B(AES_CORE_DATAPATH__abc_15863_new_n3764_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3765_));
AND2X2 AND2X2_45 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3785_), .B(AES_CORE_DATAPATH__abc_15863_new_n3786_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3787_));
AND2X2 AND2X2_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3864_), .B(AES_CORE_DATAPATH__abc_15863_new_n3865_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3866_));
AND2X2 AND2X2_47 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4440_), .B(AES_CORE_DATAPATH__abc_15863_new_n4441_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4442_));
AND2X2 AND2X2_48 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5823_), .B(AES_CORE_DATAPATH__abc_15863_new_n5824_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5825_));
AND2X2 AND2X2_49 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6788_));
AND2X2 AND2X2_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n123_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n122_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n124_));
AND2X2 AND2X2_50 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6800_));
AND2X2 AND2X2_51 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6826_));
AND2X2 AND2X2_52 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6839_));
AND2X2 AND2X2_53 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6851_));
AND2X2 AND2X2_54 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6863_));
AND2X2 AND2X2_55 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6876_));
AND2X2 AND2X2_56 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6888_));
AND2X2 AND2X2_57 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6894_));
AND2X2 AND2X2_58 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6900_));
AND2X2 AND2X2_59 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6912_));
AND2X2 AND2X2_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n158_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__3_));
AND2X2 AND2X2_60 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6925_));
AND2X2 AND2X2_61 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6937_));
AND2X2 AND2X2_62 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6943_));
AND2X2 AND2X2_63 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6955_));
AND2X2 AND2X2_64 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6974_));
AND2X2 AND2X2_65 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7003_), .B(AES_CORE_DATAPATH__abc_15863_new_n7014_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7015_));
AND2X2 AND2X2_66 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7071_), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7072_));
AND2X2 AND2X2_67 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7072_), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7078_));
AND2X2 AND2X2_68 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7113_), .B(AES_CORE_DATAPATH__abc_15863_new_n7114_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7115_));
AND2X2 AND2X2_69 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7123_), .B(AES_CORE_DATAPATH__abc_15863_new_n2632_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7125_));
AND2X2 AND2X2_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n195_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n196_));
AND2X2 AND2X2_70 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7131_), .B(AES_CORE_DATAPATH__abc_15863_new_n2640_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7133_));
AND2X2 AND2X2_71 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7115_), .B(AES_CORE_DATAPATH__abc_15863_new_n7146_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7147_));
AND2X2 AND2X2_72 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7156_), .B(AES_CORE_DATAPATH__abc_15863_new_n2660_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7158_));
AND2X2 AND2X2_73 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7196_), .B(AES_CORE_DATAPATH__abc_15863_new_n2696_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7198_));
AND2X2 AND2X2_74 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n434_));
AND2X2 AND2X2_75 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n108_));
AND2X2 AND2X2_76 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n111_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n106_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_));
AND2X2 AND2X2_77 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n140_));
AND2X2 AND2X2_78 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n52_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n57_));
AND2X2 AND2X2_79 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n145_));
AND2X2 AND2X2_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1897));
AND2X2 AND2X2_80 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n138_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n214_));
AND2X2 AND2X2_81 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n218_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n219_));
AND2X2 AND2X2_82 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n209_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n211_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n226_));
AND2X2 AND2X2_83 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n261_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n266_));
AND2X2 AND2X2_84 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n398_));
AND2X2 AND2X2_85 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_));
AND2X2 AND2X2_86 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n415_));
AND2X2 AND2X2_87 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n419_));
AND2X2 AND2X2_88 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n52_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n57_));
AND2X2 AND2X2_89 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n145_));
AND2X2 AND2X2_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1928));
AND2X2 AND2X2_90 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n138_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n214_));
AND2X2 AND2X2_91 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n218_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n219_));
AND2X2 AND2X2_92 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n209_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n211_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n226_));
AND2X2 AND2X2_93 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n261_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n266_));
AND2X2 AND2X2_94 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n398_));
AND2X2 AND2X2_95 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_));
AND2X2 AND2X2_96 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n415_));
AND2X2 AND2X2_97 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n419_));
AND2X2 AND2X2_98 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n52_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n57_));
AND2X2 AND2X2_99 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n145_));
AOI21X1 AOI21X1_1 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n75_), .B(\aes_mode[1] ), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n77_));
AOI21X1 AOI21X1_10 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n172_), .B(AES_CORE_CONTROL_UNIT_state_6_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n179_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n180_));
AOI21X1 AOI21X1_100 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_1_), .C(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3865_));
AOI21X1 AOI21X1_101 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4238_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4235_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__1_));
AOI21X1 AOI21X1_102 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4243_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4240_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__2_));
AOI21X1 AOI21X1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4248_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4245_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__3_));
AOI21X1 AOI21X1_104 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4253_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4250_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__4_));
AOI21X1 AOI21X1_105 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4258_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4255_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__5_));
AOI21X1 AOI21X1_106 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4261_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4260_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__6_));
AOI21X1 AOI21X1_107 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4264_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4263_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__7_));
AOI21X1 AOI21X1_108 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4267_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4266_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__8_));
AOI21X1 AOI21X1_109 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4270_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4269_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__9_));
AOI21X1 AOI21X1_11 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n184_));
AOI21X1 AOI21X1_110 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4273_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4272_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__10_));
AOI21X1 AOI21X1_111 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4276_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4275_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__11_));
AOI21X1 AOI21X1_112 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4281_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4278_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__12_));
AOI21X1 AOI21X1_113 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4286_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4283_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__13_));
AOI21X1 AOI21X1_114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4291_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4288_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__14_));
AOI21X1 AOI21X1_115 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4296_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4293_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__15_));
AOI21X1 AOI21X1_116 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4301_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4298_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__16_));
AOI21X1 AOI21X1_117 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4306_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4303_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__17_));
AOI21X1 AOI21X1_118 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4311_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4308_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__18_));
AOI21X1 AOI21X1_119 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4316_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4313_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__19_));
AOI21X1 AOI21X1_12 ( .A(AES_CORE_CONTROL_UNIT_state_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n187_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n188_));
AOI21X1 AOI21X1_120 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4321_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4318_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__20_));
AOI21X1 AOI21X1_121 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4326_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4323_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__21_));
AOI21X1 AOI21X1_122 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4331_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4328_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__22_));
AOI21X1 AOI21X1_123 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4336_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4333_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__23_));
AOI21X1 AOI21X1_124 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4341_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4338_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__24_));
AOI21X1 AOI21X1_125 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4346_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4343_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__25_));
AOI21X1 AOI21X1_126 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4351_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4348_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__26_));
AOI21X1 AOI21X1_127 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4356_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4353_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__27_));
AOI21X1 AOI21X1_128 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4361_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4358_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__28_));
AOI21X1 AOI21X1_129 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4366_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4363_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__29_));
AOI21X1 AOI21X1_13 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_6_), .C(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n199_));
AOI21X1 AOI21X1_130 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4371_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4368_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__30_));
AOI21X1 AOI21X1_131 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4373_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4374_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__31_));
AOI21X1 AOI21X1_132 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3873_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4378_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__1_));
AOI21X1 AOI21X1_133 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3878_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4380_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__2_));
AOI21X1 AOI21X1_134 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3883_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4382_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__3_));
AOI21X1 AOI21X1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3888_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4384_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__4_));
AOI21X1 AOI21X1_136 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3893_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4386_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__5_));
AOI21X1 AOI21X1_137 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3898_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4388_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__6_));
AOI21X1 AOI21X1_138 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3903_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4390_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__7_));
AOI21X1 AOI21X1_139 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3908_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4392_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__8_));
AOI21X1 AOI21X1_14 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n179_), .C(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n204_));
AOI21X1 AOI21X1_140 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3913_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4394_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__9_));
AOI21X1 AOI21X1_141 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3918_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4396_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__10_));
AOI21X1 AOI21X1_142 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3923_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4398_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__11_));
AOI21X1 AOI21X1_143 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3928_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4400_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__12_));
AOI21X1 AOI21X1_144 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3933_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4402_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__13_));
AOI21X1 AOI21X1_145 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3938_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4404_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__14_));
AOI21X1 AOI21X1_146 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3943_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4406_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__15_));
AOI21X1 AOI21X1_147 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3948_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4408_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__16_));
AOI21X1 AOI21X1_148 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3953_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4410_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__17_));
AOI21X1 AOI21X1_149 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3958_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4412_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__18_));
AOI21X1 AOI21X1_15 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_3_), .C(AES_CORE_DATAPATH_col_en_host_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2460_));
AOI21X1 AOI21X1_150 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3963_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4414_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__19_));
AOI21X1 AOI21X1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3968_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4416_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__20_));
AOI21X1 AOI21X1_152 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3973_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4418_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__21_));
AOI21X1 AOI21X1_153 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3978_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4420_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__22_));
AOI21X1 AOI21X1_154 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3983_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4422_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__23_));
AOI21X1 AOI21X1_155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3988_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4424_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__24_));
AOI21X1 AOI21X1_156 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3993_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4426_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__25_));
AOI21X1 AOI21X1_157 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3998_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4428_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__26_));
AOI21X1 AOI21X1_158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4003_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4430_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__27_));
AOI21X1 AOI21X1_159 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4008_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4432_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__28_));
AOI21X1 AOI21X1_16 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_2_), .C(AES_CORE_DATAPATH_col_en_host_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2465_));
AOI21X1 AOI21X1_160 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4013_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4434_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__29_));
AOI21X1 AOI21X1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4018_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4436_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__30_));
AOI21X1 AOI21X1_162 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4025_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4438_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__31_));
AOI21X1 AOI21X1_163 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2712_), .B(AES_CORE_DATAPATH_key_en_pp1_2_), .C(start), .Y(AES_CORE_DATAPATH__abc_15863_new_n4440_));
AOI21X1 AOI21X1_164 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_2_), .C(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4441_));
AOI21X1 AOI21X1_165 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2740_), .B(AES_CORE_DATAPATH__abc_15863_new_n3104_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4589_));
AOI21X1 AOI21X1_166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4617_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4619_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4620_));
AOI21X1 AOI21X1_167 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4660_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4661_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4662_));
AOI21X1 AOI21X1_168 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2764_), .B(AES_CORE_DATAPATH__abc_15863_new_n3150_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4676_));
AOI21X1 AOI21X1_169 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4699_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4700_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4701_));
AOI21X1 AOI21X1_17 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_1_), .C(AES_CORE_DATAPATH_col_en_host_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2472_));
AOI21X1 AOI21X1_170 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4737_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4738_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4739_));
AOI21X1 AOI21X1_171 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2784_), .B(AES_CORE_DATAPATH__abc_15863_new_n3195_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4755_));
AOI21X1 AOI21X1_172 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_bkp_1__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4761_));
AOI21X1 AOI21X1_173 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n4763_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4764_));
AOI21X1 AOI21X1_174 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4775_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4776_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4777_));
AOI21X1 AOI21X1_175 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2794_), .B(AES_CORE_DATAPATH__abc_15863_new_n3217_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4791_));
AOI21X1 AOI21X1_176 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4814_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4815_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4816_));
AOI21X1 AOI21X1_177 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2804_), .B(AES_CORE_DATAPATH__abc_15863_new_n3239_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4830_));
AOI21X1 AOI21X1_178 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_bkp_1__6_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4836_));
AOI21X1 AOI21X1_179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n4838_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4839_));
AOI21X1 AOI21X1_18 ( .A(AES_CORE_CONTROL_UNIT_col_en_0_), .B(AES_CORE_CONTROL_UNIT_bypass_rk), .C(AES_CORE_DATAPATH_col_en_host_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2477_));
AOI21X1 AOI21X1_180 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4849_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4850_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4851_));
AOI21X1 AOI21X1_181 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4888_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4889_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4890_));
AOI21X1 AOI21X1_182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2828_), .B(AES_CORE_DATAPATH__abc_15863_new_n3283_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4904_));
AOI21X1 AOI21X1_183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_bkp_1__8_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4910_));
AOI21X1 AOI21X1_184 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n4912_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4913_));
AOI21X1 AOI21X1_185 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4923_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4924_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4925_));
AOI21X1 AOI21X1_186 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4961_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n4962_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4963_));
AOI21X1 AOI21X1_187 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2851_), .B(AES_CORE_DATAPATH__abc_15863_new_n3327_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4978_));
AOI21X1 AOI21X1_188 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5001_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5002_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5003_));
AOI21X1 AOI21X1_189 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5039_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5040_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5041_));
AOI21X1 AOI21X1_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2481_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2483_));
AOI21X1 AOI21X1_190 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2870_), .B(AES_CORE_DATAPATH__abc_15863_new_n3371_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5056_));
AOI21X1 AOI21X1_191 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5079_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5081_));
AOI21X1 AOI21X1_192 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5117_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5118_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5119_));
AOI21X1 AOI21X1_193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2890_), .B(AES_CORE_DATAPATH__abc_15863_new_n3415_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5134_));
AOI21X1 AOI21X1_194 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_bkp_1__14_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5140_));
AOI21X1 AOI21X1_195 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n5142_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5143_));
AOI21X1 AOI21X1_196 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5154_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5155_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5156_));
AOI21X1 AOI21X1_197 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5192_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5193_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5194_));
AOI21X1 AOI21X1_198 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2911_), .B(AES_CORE_DATAPATH__abc_15863_new_n3459_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5209_));
AOI21X1 AOI21X1_199 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5232_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5233_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5234_));
AOI21X1 AOI21X1_2 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n93_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n88_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n85_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_5_));
AOI21X1 AOI21X1_20 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__1_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2488_));
AOI21X1 AOI21X1_200 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5270_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5271_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5272_));
AOI21X1 AOI21X1_201 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5309_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5310_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5311_));
AOI21X1 AOI21X1_202 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5348_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5349_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5350_));
AOI21X1 AOI21X1_203 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2951_), .B(AES_CORE_DATAPATH__abc_15863_new_n3547_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5365_));
AOI21X1 AOI21X1_204 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5388_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5389_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5390_));
AOI21X1 AOI21X1_205 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5426_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5427_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5428_));
AOI21X1 AOI21X1_206 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2973_), .B(AES_CORE_DATAPATH__abc_15863_new_n3591_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5443_));
AOI21X1 AOI21X1_207 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_bkp_1__22_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5449_));
AOI21X1 AOI21X1_208 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n5451_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5452_));
AOI21X1 AOI21X1_209 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5463_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5464_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5465_));
AOI21X1 AOI21X1_21 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2490_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2491_));
AOI21X1 AOI21X1_210 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5502_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5503_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5504_));
AOI21X1 AOI21X1_211 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2997_), .B(AES_CORE_DATAPATH__abc_15863_new_n3635_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5518_));
AOI21X1 AOI21X1_212 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5541_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5542_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5543_));
AOI21X1 AOI21X1_213 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5579_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5581_));
AOI21X1 AOI21X1_214 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5618_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5619_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5620_));
AOI21X1 AOI21X1_215 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3029_), .B(AES_CORE_DATAPATH__abc_15863_new_n3701_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5635_));
AOI21X1 AOI21X1_216 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5658_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5659_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5660_));
AOI21X1 AOI21X1_217 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5696_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5697_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5698_));
AOI21X1 AOI21X1_218 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3050_), .B(AES_CORE_DATAPATH__abc_15863_new_n3745_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5713_));
AOI21X1 AOI21X1_219 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_bkp_1__29_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5719_));
AOI21X1 AOI21X1_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__2_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2496_));
AOI21X1 AOI21X1_220 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n5721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5722_));
AOI21X1 AOI21X1_221 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5733_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5734_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5735_));
AOI21X1 AOI21X1_222 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3060_), .B(AES_CORE_DATAPATH__abc_15863_new_n3767_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5749_));
AOI21X1 AOI21X1_223 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5772_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5773_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5774_));
AOI21X1 AOI21X1_224 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5810_), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_DATAPATH__abc_15863_new_n5811_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5812_));
AOI21X1 AOI21X1_225 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2712_), .B(AES_CORE_DATAPATH_key_en_pp1_3_), .C(start), .Y(AES_CORE_DATAPATH__abc_15863_new_n5823_));
AOI21X1 AOI21X1_226 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_3_), .C(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5824_));
AOI21X1 AOI21X1_227 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5831_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n5989_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__1_));
AOI21X1 AOI21X1_228 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5836_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n5991_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__2_));
AOI21X1 AOI21X1_229 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5841_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n5993_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__3_));
AOI21X1 AOI21X1_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__3_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2502_));
AOI21X1 AOI21X1_230 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5846_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n5995_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__4_));
AOI21X1 AOI21X1_231 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5851_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n5997_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__5_));
AOI21X1 AOI21X1_232 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5856_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n5999_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__6_));
AOI21X1 AOI21X1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5861_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6001_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__7_));
AOI21X1 AOI21X1_234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6003_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__8_));
AOI21X1 AOI21X1_235 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5871_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6005_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__9_));
AOI21X1 AOI21X1_236 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5876_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6007_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__10_));
AOI21X1 AOI21X1_237 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5881_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6009_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__11_));
AOI21X1 AOI21X1_238 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5886_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6011_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__12_));
AOI21X1 AOI21X1_239 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5891_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6013_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__13_));
AOI21X1 AOI21X1_24 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2504_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2505_));
AOI21X1 AOI21X1_240 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5896_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6015_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__14_));
AOI21X1 AOI21X1_241 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5901_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6017_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__15_));
AOI21X1 AOI21X1_242 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5906_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6019_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__16_));
AOI21X1 AOI21X1_243 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5911_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6021_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__17_));
AOI21X1 AOI21X1_244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5916_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6023_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__18_));
AOI21X1 AOI21X1_245 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5921_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6025_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__19_));
AOI21X1 AOI21X1_246 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5926_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6027_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__20_));
AOI21X1 AOI21X1_247 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5931_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6029_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__21_));
AOI21X1 AOI21X1_248 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5936_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6031_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__22_));
AOI21X1 AOI21X1_249 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5941_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6033_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__23_));
AOI21X1 AOI21X1_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2510_));
AOI21X1 AOI21X1_250 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5946_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6035_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__24_));
AOI21X1 AOI21X1_251 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5951_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6037_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__25_));
AOI21X1 AOI21X1_252 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5956_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6039_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__26_));
AOI21X1 AOI21X1_253 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5961_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6041_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__27_));
AOI21X1 AOI21X1_254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5966_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6043_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__28_));
AOI21X1 AOI21X1_255 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5971_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6045_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__29_));
AOI21X1 AOI21X1_256 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5976_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6047_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__30_));
AOI21X1 AOI21X1_257 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5982_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6049_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__31_));
AOI21X1 AOI21X1_258 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6779_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6780_));
AOI21X1 AOI21X1_259 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6785_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6786_));
AOI21X1 AOI21X1_26 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__5_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2516_));
AOI21X1 AOI21X1_260 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6791_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6792_));
AOI21X1 AOI21X1_261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6797_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6798_));
AOI21X1 AOI21X1_262 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6804_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6805_));
AOI21X1 AOI21X1_263 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6810_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6811_));
AOI21X1 AOI21X1_264 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6817_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6818_));
AOI21X1 AOI21X1_265 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6823_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6824_));
AOI21X1 AOI21X1_266 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6830_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6831_));
AOI21X1 AOI21X1_267 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6836_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6837_));
AOI21X1 AOI21X1_268 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6842_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6843_));
AOI21X1 AOI21X1_269 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6848_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6849_));
AOI21X1 AOI21X1_27 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2524_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2525_));
AOI21X1 AOI21X1_270 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6854_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6855_));
AOI21X1 AOI21X1_271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6860_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6861_));
AOI21X1 AOI21X1_272 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6867_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6868_));
AOI21X1 AOI21X1_273 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6873_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6874_));
AOI21X1 AOI21X1_274 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6879_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6880_));
AOI21X1 AOI21X1_275 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6885_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6886_));
AOI21X1 AOI21X1_276 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6891_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6892_));
AOI21X1 AOI21X1_277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6897_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6898_));
AOI21X1 AOI21X1_278 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6903_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6904_));
AOI21X1 AOI21X1_279 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6909_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6910_));
AOI21X1 AOI21X1_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2532_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2533_));
AOI21X1 AOI21X1_280 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6916_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6917_));
AOI21X1 AOI21X1_281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6922_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6923_));
AOI21X1 AOI21X1_282 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6928_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6929_));
AOI21X1 AOI21X1_283 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6934_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6935_));
AOI21X1 AOI21X1_284 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6940_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6941_));
AOI21X1 AOI21X1_285 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6946_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6947_));
AOI21X1 AOI21X1_286 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6952_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6953_));
AOI21X1 AOI21X1_287 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6959_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6960_));
AOI21X1 AOI21X1_288 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6965_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6966_));
AOI21X1 AOI21X1_289 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6971_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n6972_));
AOI21X1 AOI21X1_29 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2540_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2541_));
AOI21X1 AOI21X1_290 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7013_), .B(AES_CORE_DATAPATH__abc_15863_new_n2514_), .C(AES_CORE_DATAPATH__abc_15863_new_n7015_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7016_));
AOI21X1 AOI21X1_291 ( .A(\bus_in[9] ), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .C(AES_CORE_DATAPATH__abc_15863_new_n6977_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7045_));
AOI21X1 AOI21X1_292 ( .A(\bus_in[10] ), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .C(AES_CORE_DATAPATH__abc_15863_new_n6977_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7052_));
AOI21X1 AOI21X1_293 ( .A(\bus_in[11] ), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .C(AES_CORE_DATAPATH__abc_15863_new_n6977_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7058_));
AOI21X1 AOI21X1_294 ( .A(AES_CORE_DATAPATH_iv_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7063_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7064_));
AOI21X1 AOI21X1_295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7060_), .B(AES_CORE_DATAPATH__abc_15863_new_n2574_), .C(AES_CORE_DATAPATH__abc_15863_new_n6982_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7066_));
AOI21X1 AOI21X1_296 ( .A(AES_CORE_DATAPATH_iv_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7068_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7069_));
AOI21X1 AOI21X1_297 ( .A(AES_CORE_DATAPATH_iv_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7075_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7076_));
AOI21X1 AOI21X1_298 ( .A(AES_CORE_DATAPATH_iv_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7081_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7082_));
AOI21X1 AOI21X1_299 ( .A(AES_CORE_DATAPATH_iv_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7088_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7089_));
AOI21X1 AOI21X1_3 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n116_), .B(AES_CORE_CONTROL_UNIT_key_gen), .C(AES_CORE_CONTROL_UNIT_state_15_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n117_));
AOI21X1 AOI21X1_30 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2548_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2549_));
AOI21X1 AOI21X1_300 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7084_), .B(AES_CORE_DATAPATH__abc_15863_new_n2602_), .C(AES_CORE_DATAPATH__abc_15863_new_n6982_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7091_));
AOI21X1 AOI21X1_301 ( .A(AES_CORE_DATAPATH_iv_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7093_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7094_));
AOI21X1 AOI21X1_302 ( .A(AES_CORE_DATAPATH_iv_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7100_));
AOI21X1 AOI21X1_303 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7097_), .B(AES_CORE_DATAPATH__abc_15863_new_n2618_), .C(AES_CORE_DATAPATH__abc_15863_new_n6982_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7102_));
AOI21X1 AOI21X1_304 ( .A(AES_CORE_DATAPATH_iv_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7104_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7105_));
AOI21X1 AOI21X1_305 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7112_), .B(AES_CORE_DATAPATH__abc_15863_new_n7115_), .C(AES_CORE_DATAPATH__abc_15863_new_n2626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7116_));
AOI21X1 AOI21X1_306 ( .A(AES_CORE_DATAPATH_iv_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7120_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7121_));
AOI21X1 AOI21X1_307 ( .A(AES_CORE_DATAPATH_iv_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7127_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7128_));
AOI21X1 AOI21X1_308 ( .A(AES_CORE_DATAPATH_iv_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7135_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7136_));
AOI21X1 AOI21X1_309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7131_), .B(AES_CORE_DATAPATH_iv_3__22_), .C(AES_CORE_DATAPATH__abc_15863_new_n2646_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7138_));
AOI21X1 AOI21X1_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2556_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2557_));
AOI21X1 AOI21X1_310 ( .A(AES_CORE_DATAPATH_iv_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7142_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7143_));
AOI21X1 AOI21X1_311 ( .A(AES_CORE_DATAPATH_iv_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7153_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7154_));
AOI21X1 AOI21X1_312 ( .A(AES_CORE_DATAPATH_iv_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7160_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7161_));
AOI21X1 AOI21X1_313 ( .A(AES_CORE_DATAPATH_iv_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7169_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7170_));
AOI21X1 AOI21X1_314 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7165_), .B(AES_CORE_DATAPATH_iv_3__26_), .C(AES_CORE_DATAPATH__abc_15863_new_n2676_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7172_));
AOI21X1 AOI21X1_315 ( .A(AES_CORE_DATAPATH_iv_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7176_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7177_));
AOI21X1 AOI21X1_316 ( .A(AES_CORE_DATAPATH_iv_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7185_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7186_));
AOI21X1 AOI21X1_317 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7180_), .B(AES_CORE_DATAPATH_iv_3__28_), .C(AES_CORE_DATAPATH__abc_15863_new_n2690_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7188_));
AOI21X1 AOI21X1_318 ( .A(AES_CORE_DATAPATH_iv_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7192_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7193_));
AOI21X1 AOI21X1_319 ( .A(AES_CORE_DATAPATH_iv_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7200_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7201_));
AOI21X1 AOI21X1_32 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2564_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2565_));
AOI21X1 AOI21X1_320 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7196_), .B(AES_CORE_DATAPATH_iv_3__30_), .C(AES_CORE_DATAPATH__abc_15863_new_n2702_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7203_));
AOI21X1 AOI21X1_321 ( .A(AES_CORE_DATAPATH_iv_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .C(AES_CORE_DATAPATH__abc_15863_new_n7207_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7208_));
AOI21X1 AOI21X1_322 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4241_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7214_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__2_));
AOI21X1 AOI21X1_323 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4251_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7218_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__4_));
AOI21X1 AOI21X1_324 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4256_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7220_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__5_));
AOI21X1 AOI21X1_325 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4279_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7234_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__12_));
AOI21X1 AOI21X1_326 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4289_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7238_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__14_));
AOI21X1 AOI21X1_327 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4299_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7242_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__16_));
AOI21X1 AOI21X1_328 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4319_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7250_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__20_));
AOI21X1 AOI21X1_329 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4329_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7254_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__22_));
AOI21X1 AOI21X1_33 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__12_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2570_));
AOI21X1 AOI21X1_330 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4339_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7258_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__24_));
AOI21X1 AOI21X1_331 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4354_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7264_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__27_));
AOI21X1 AOI21X1_332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4364_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7268_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__29_));
AOI21X1 AOI21X1_333 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4369_), .B(\iv_en[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7270_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__30_));
AOI21X1 AOI21X1_334 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7339_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7340_));
AOI21X1 AOI21X1_335 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7344_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7345_));
AOI21X1 AOI21X1_336 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7349_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7350_));
AOI21X1 AOI21X1_337 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7354_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7355_));
AOI21X1 AOI21X1_338 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7359_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7360_));
AOI21X1 AOI21X1_339 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7364_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7365_));
AOI21X1 AOI21X1_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__13_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2576_));
AOI21X1 AOI21X1_340 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7369_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7370_));
AOI21X1 AOI21X1_341 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7374_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7375_));
AOI21X1 AOI21X1_342 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7379_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7380_));
AOI21X1 AOI21X1_343 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7384_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7385_));
AOI21X1 AOI21X1_344 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7389_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7390_));
AOI21X1 AOI21X1_345 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7394_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7395_));
AOI21X1 AOI21X1_346 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7399_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7400_));
AOI21X1 AOI21X1_347 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7404_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7405_));
AOI21X1 AOI21X1_348 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7409_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7410_));
AOI21X1 AOI21X1_349 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7414_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7415_));
AOI21X1 AOI21X1_35 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2578_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2579_));
AOI21X1 AOI21X1_350 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7419_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7420_));
AOI21X1 AOI21X1_351 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7424_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7425_));
AOI21X1 AOI21X1_352 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7429_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7430_));
AOI21X1 AOI21X1_353 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7434_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7435_));
AOI21X1 AOI21X1_354 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7439_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7440_));
AOI21X1 AOI21X1_355 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7444_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7445_));
AOI21X1 AOI21X1_356 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7449_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7450_));
AOI21X1 AOI21X1_357 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7454_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7455_));
AOI21X1 AOI21X1_358 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7459_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7460_));
AOI21X1 AOI21X1_359 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7464_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7465_));
AOI21X1 AOI21X1_36 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__14_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2584_));
AOI21X1 AOI21X1_360 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7469_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7470_));
AOI21X1 AOI21X1_361 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7474_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7475_));
AOI21X1 AOI21X1_362 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7479_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7480_));
AOI21X1 AOI21X1_363 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7484_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7485_));
AOI21X1 AOI21X1_364 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7489_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7490_));
AOI21X1 AOI21X1_365 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7494_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7495_));
AOI21X1 AOI21X1_366 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4236_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7501_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__1_));
AOI21X1 AOI21X1_367 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4241_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7503_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__2_));
AOI21X1 AOI21X1_368 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4246_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7505_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__3_));
AOI21X1 AOI21X1_369 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4251_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7507_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__4_));
AOI21X1 AOI21X1_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__15_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2590_));
AOI21X1 AOI21X1_370 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4256_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7509_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__5_));
AOI21X1 AOI21X1_371 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4279_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7523_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__12_));
AOI21X1 AOI21X1_372 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4284_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7525_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__13_));
AOI21X1 AOI21X1_373 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4289_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7527_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__14_));
AOI21X1 AOI21X1_374 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4294_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7529_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__15_));
AOI21X1 AOI21X1_375 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4299_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7531_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__16_));
AOI21X1 AOI21X1_376 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4304_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7533_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__17_));
AOI21X1 AOI21X1_377 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4309_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7535_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__18_));
AOI21X1 AOI21X1_378 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4314_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7537_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__19_));
AOI21X1 AOI21X1_379 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4319_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7539_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__20_));
AOI21X1 AOI21X1_38 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2592_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2593_));
AOI21X1 AOI21X1_380 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4324_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7541_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__21_));
AOI21X1 AOI21X1_381 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4329_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7543_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__22_));
AOI21X1 AOI21X1_382 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4334_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7545_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__23_));
AOI21X1 AOI21X1_383 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4339_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7547_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__24_));
AOI21X1 AOI21X1_384 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4344_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7549_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__25_));
AOI21X1 AOI21X1_385 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4349_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7551_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__26_));
AOI21X1 AOI21X1_386 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4354_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7553_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__27_));
AOI21X1 AOI21X1_387 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4359_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7555_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__28_));
AOI21X1 AOI21X1_388 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4364_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7557_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__29_));
AOI21X1 AOI21X1_389 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4369_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7559_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__30_));
AOI21X1 AOI21X1_39 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__16_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2598_));
AOI21X1 AOI21X1_390 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4023_), .B(\iv_en[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7561_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__31_));
AOI21X1 AOI21X1_391 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7566_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7567_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__1_));
AOI21X1 AOI21X1_392 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7571_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7572_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__3_));
AOI21X1 AOI21X1_393 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7580_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7581_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__7_));
AOI21X1 AOI21X1_394 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7585_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7586_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__9_));
AOI21X1 AOI21X1_395 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7590_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7591_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__11_));
AOI21X1 AOI21X1_396 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7595_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7596_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__13_));
AOI21X1 AOI21X1_397 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7600_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7601_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__15_));
AOI21X1 AOI21X1_398 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7605_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7606_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__17_));
AOI21X1 AOI21X1_399 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7608_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7609_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__18_));
AOI21X1 AOI21X1_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n136_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n135_), .C(disable_core), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_4_));
AOI21X1 AOI21X1_40 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__17_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2604_));
AOI21X1 AOI21X1_400 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7611_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7612_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__19_));
AOI21X1 AOI21X1_401 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7616_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7617_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__21_));
AOI21X1 AOI21X1_402 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7621_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7622_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__23_));
AOI21X1 AOI21X1_403 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7626_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7627_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__25_));
AOI21X1 AOI21X1_404 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7629_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7630_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__26_));
AOI21X1 AOI21X1_405 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7634_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7635_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__28_));
AOI21X1 AOI21X1_406 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7641_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7642_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__31_));
AOI21X1 AOI21X1_407 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7645_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7646_));
AOI21X1 AOI21X1_408 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7566_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7651_));
AOI21X1 AOI21X1_409 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7656_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7657_));
AOI21X1 AOI21X1_41 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2606_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2607_));
AOI21X1 AOI21X1_410 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7571_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7662_));
AOI21X1 AOI21X1_411 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7667_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7668_));
AOI21X1 AOI21X1_412 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7673_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7674_));
AOI21X1 AOI21X1_413 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7679_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7680_));
AOI21X1 AOI21X1_414 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7580_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7685_));
AOI21X1 AOI21X1_415 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7690_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7691_));
AOI21X1 AOI21X1_416 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7585_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7696_));
AOI21X1 AOI21X1_417 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7701_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7702_));
AOI21X1 AOI21X1_418 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7590_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7707_));
AOI21X1 AOI21X1_419 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7712_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7713_));
AOI21X1 AOI21X1_42 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__18_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2612_));
AOI21X1 AOI21X1_420 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7595_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7718_));
AOI21X1 AOI21X1_421 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7723_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7724_));
AOI21X1 AOI21X1_422 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7600_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7729_));
AOI21X1 AOI21X1_423 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7734_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7735_));
AOI21X1 AOI21X1_424 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7605_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7740_));
AOI21X1 AOI21X1_425 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7608_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7745_));
AOI21X1 AOI21X1_426 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7611_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7750_));
AOI21X1 AOI21X1_427 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7755_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7756_));
AOI21X1 AOI21X1_428 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7616_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7761_));
AOI21X1 AOI21X1_429 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7766_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7767_));
AOI21X1 AOI21X1_43 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2614_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2615_));
AOI21X1 AOI21X1_430 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7621_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7772_));
AOI21X1 AOI21X1_431 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7777_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7778_));
AOI21X1 AOI21X1_432 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7626_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7783_));
AOI21X1 AOI21X1_433 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7629_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7788_));
AOI21X1 AOI21X1_434 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7793_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7794_));
AOI21X1 AOI21X1_435 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7634_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7799_));
AOI21X1 AOI21X1_436 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7804_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7805_));
AOI21X1 AOI21X1_437 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7810_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7811_));
AOI21X1 AOI21X1_438 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7641_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7816_));
AOI21X1 AOI21X1_439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4231_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7820_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__0_));
AOI21X1 AOI21X1_44 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__19_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2620_));
AOI21X1 AOI21X1_440 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4236_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7822_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__1_));
AOI21X1 AOI21X1_441 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4241_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7824_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__2_));
AOI21X1 AOI21X1_442 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4246_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7826_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__3_));
AOI21X1 AOI21X1_443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4251_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7828_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__4_));
AOI21X1 AOI21X1_444 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4256_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7830_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__5_));
AOI21X1 AOI21X1_445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4279_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7850_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__12_));
AOI21X1 AOI21X1_446 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4284_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7852_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__13_));
AOI21X1 AOI21X1_447 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4289_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7854_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__14_));
AOI21X1 AOI21X1_448 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4294_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7856_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__15_));
AOI21X1 AOI21X1_449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4299_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7858_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__16_));
AOI21X1 AOI21X1_45 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2622_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2623_));
AOI21X1 AOI21X1_450 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4304_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7860_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__17_));
AOI21X1 AOI21X1_451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4309_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7862_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__18_));
AOI21X1 AOI21X1_452 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4314_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7864_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__19_));
AOI21X1 AOI21X1_453 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4319_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7866_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__20_));
AOI21X1 AOI21X1_454 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4324_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7868_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__21_));
AOI21X1 AOI21X1_455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4329_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7870_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__22_));
AOI21X1 AOI21X1_456 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4334_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7872_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__23_));
AOI21X1 AOI21X1_457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4339_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7874_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__24_));
AOI21X1 AOI21X1_458 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4344_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7876_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__25_));
AOI21X1 AOI21X1_459 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4349_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7878_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__26_));
AOI21X1 AOI21X1_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__20_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2628_));
AOI21X1 AOI21X1_460 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4354_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7880_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__27_));
AOI21X1 AOI21X1_461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4359_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7882_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__28_));
AOI21X1 AOI21X1_462 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4364_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7884_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__29_));
AOI21X1 AOI21X1_463 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4369_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7886_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__30_));
AOI21X1 AOI21X1_464 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4023_), .B(\iv_en[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n7888_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__31_));
AOI21X1 AOI21X1_465 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7956_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7957_));
AOI21X1 AOI21X1_466 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7962_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7963_));
AOI21X1 AOI21X1_467 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7968_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7969_));
AOI21X1 AOI21X1_468 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7974_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7975_));
AOI21X1 AOI21X1_469 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7980_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7981_));
AOI21X1 AOI21X1_47 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__21_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2634_));
AOI21X1 AOI21X1_470 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7986_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7987_));
AOI21X1 AOI21X1_471 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7992_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7993_));
AOI21X1 AOI21X1_472 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n7998_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n7999_));
AOI21X1 AOI21X1_473 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8004_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8005_));
AOI21X1 AOI21X1_474 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8010_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8011_));
AOI21X1 AOI21X1_475 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8016_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8017_));
AOI21X1 AOI21X1_476 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8022_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8023_));
AOI21X1 AOI21X1_477 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8028_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8029_));
AOI21X1 AOI21X1_478 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8034_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8035_));
AOI21X1 AOI21X1_479 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8040_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8041_));
AOI21X1 AOI21X1_48 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2636_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2637_));
AOI21X1 AOI21X1_480 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8046_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8047_));
AOI21X1 AOI21X1_481 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8052_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8053_));
AOI21X1 AOI21X1_482 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8058_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8059_));
AOI21X1 AOI21X1_483 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8064_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8065_));
AOI21X1 AOI21X1_484 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8070_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8071_));
AOI21X1 AOI21X1_485 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8076_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8077_));
AOI21X1 AOI21X1_486 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8082_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8083_));
AOI21X1 AOI21X1_487 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8088_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8089_));
AOI21X1 AOI21X1_488 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8094_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8095_));
AOI21X1 AOI21X1_489 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8100_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8101_));
AOI21X1 AOI21X1_49 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__22_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2642_));
AOI21X1 AOI21X1_490 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8106_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8107_));
AOI21X1 AOI21X1_491 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8112_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8113_));
AOI21X1 AOI21X1_492 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8118_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8119_));
AOI21X1 AOI21X1_493 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8124_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8125_));
AOI21X1 AOI21X1_494 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8130_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8131_));
AOI21X1 AOI21X1_495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8136_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8137_));
AOI21X1 AOI21X1_496 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n8142_), .C(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n8143_));
AOI21X1 AOI21X1_497 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n404_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n406_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n402_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n407_));
AOI21X1 AOI21X1_498 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n414_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n401_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n415_));
AOI21X1 AOI21X1_499 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n412_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n441_));
AOI21X1 AOI21X1_5 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT_state_7_), .C(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_));
AOI21X1 AOI21X1_50 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__23_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2648_));
AOI21X1 AOI21X1_500 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n216_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n221_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n259_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n260_));
AOI21X1 AOI21X1_501 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n262_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n214_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n144_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n263_));
AOI21X1 AOI21X1_502 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n303_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n304_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n305_));
AOI21X1 AOI21X1_503 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n306_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n307_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n299_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n308_));
AOI21X1 AOI21X1_504 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n113_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n119_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n366_));
AOI21X1 AOI21X1_505 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n209_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n212_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n259_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n387_));
AOI21X1 AOI21X1_506 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n424_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n425_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n421_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n426_));
AOI21X1 AOI21X1_507 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n427_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n428_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n429_));
AOI21X1 AOI21X1_508 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n424_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n425_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n523_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n524_));
AOI21X1 AOI21X1_509 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n427_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n428_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n525_));
AOI21X1 AOI21X1_51 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2650_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2651_));
AOI21X1 AOI21X1_510 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n66_));
AOI21X1 AOI21X1_511 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n77_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n78_));
AOI21X1 AOI21X1_512 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n88_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_));
AOI21X1 AOI21X1_513 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n71_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n90_));
AOI21X1 AOI21X1_514 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n75_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n86_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n92_));
AOI21X1 AOI21X1_515 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n91_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n93_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_));
AOI21X1 AOI21X1_516 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n115_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n117_));
AOI21X1 AOI21X1_517 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n122_));
AOI21X1 AOI21X1_518 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n157_));
AOI21X1 AOI21X1_519 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n175_));
AOI21X1 AOI21X1_52 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__24_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2656_));
AOI21X1 AOI21X1_520 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n231_));
AOI21X1 AOI21X1_521 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n181_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n240_));
AOI21X1 AOI21X1_522 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n237_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n212_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n270_));
AOI21X1 AOI21X1_523 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n245_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n226_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n271_));
AOI21X1 AOI21X1_524 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n293_));
AOI21X1 AOI21X1_525 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n302_));
AOI21X1 AOI21X1_526 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n307_));
AOI21X1 AOI21X1_527 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n311_));
AOI21X1 AOI21X1_528 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n312_));
AOI21X1 AOI21X1_529 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n387_));
AOI21X1 AOI21X1_53 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__25_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2662_));
AOI21X1 AOI21X1_530 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n395_));
AOI21X1 AOI21X1_531 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n445_));
AOI21X1 AOI21X1_532 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n446_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n447_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n448_));
AOI21X1 AOI21X1_533 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n435_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n450_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n451_));
AOI21X1 AOI21X1_534 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n66_));
AOI21X1 AOI21X1_535 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n77_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n78_));
AOI21X1 AOI21X1_536 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n88_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_));
AOI21X1 AOI21X1_537 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n71_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n90_));
AOI21X1 AOI21X1_538 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n75_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n86_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n92_));
AOI21X1 AOI21X1_539 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n91_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n93_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_));
AOI21X1 AOI21X1_54 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2664_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2665_));
AOI21X1 AOI21X1_540 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n115_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n117_));
AOI21X1 AOI21X1_541 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n122_));
AOI21X1 AOI21X1_542 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n157_));
AOI21X1 AOI21X1_543 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n175_));
AOI21X1 AOI21X1_544 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n231_));
AOI21X1 AOI21X1_545 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n181_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n240_));
AOI21X1 AOI21X1_546 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n237_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n212_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n270_));
AOI21X1 AOI21X1_547 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n245_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n226_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n271_));
AOI21X1 AOI21X1_548 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n293_));
AOI21X1 AOI21X1_549 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n302_));
AOI21X1 AOI21X1_55 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__26_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2670_));
AOI21X1 AOI21X1_550 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n307_));
AOI21X1 AOI21X1_551 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n311_));
AOI21X1 AOI21X1_552 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n312_));
AOI21X1 AOI21X1_553 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n387_));
AOI21X1 AOI21X1_554 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n395_));
AOI21X1 AOI21X1_555 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n445_));
AOI21X1 AOI21X1_556 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n446_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n447_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n448_));
AOI21X1 AOI21X1_557 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n435_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n450_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n451_));
AOI21X1 AOI21X1_558 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n66_));
AOI21X1 AOI21X1_559 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n77_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n78_));
AOI21X1 AOI21X1_56 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2672_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2673_));
AOI21X1 AOI21X1_560 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n88_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_));
AOI21X1 AOI21X1_561 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n71_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n90_));
AOI21X1 AOI21X1_562 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n75_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n86_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n92_));
AOI21X1 AOI21X1_563 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n91_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n93_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_));
AOI21X1 AOI21X1_564 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n115_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n117_));
AOI21X1 AOI21X1_565 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n122_));
AOI21X1 AOI21X1_566 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n157_));
AOI21X1 AOI21X1_567 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n175_));
AOI21X1 AOI21X1_568 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n231_));
AOI21X1 AOI21X1_569 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n181_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n240_));
AOI21X1 AOI21X1_57 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__27_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2678_));
AOI21X1 AOI21X1_570 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n237_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n212_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n270_));
AOI21X1 AOI21X1_571 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n245_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n226_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n271_));
AOI21X1 AOI21X1_572 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n293_));
AOI21X1 AOI21X1_573 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n302_));
AOI21X1 AOI21X1_574 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n307_));
AOI21X1 AOI21X1_575 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n311_));
AOI21X1 AOI21X1_576 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n312_));
AOI21X1 AOI21X1_577 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n387_));
AOI21X1 AOI21X1_578 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n395_));
AOI21X1 AOI21X1_579 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n445_));
AOI21X1 AOI21X1_58 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__28_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2684_));
AOI21X1 AOI21X1_580 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n446_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n447_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n448_));
AOI21X1 AOI21X1_581 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n435_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n450_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n451_));
AOI21X1 AOI21X1_582 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n66_));
AOI21X1 AOI21X1_583 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n77_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n78_));
AOI21X1 AOI21X1_584 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n88_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_));
AOI21X1 AOI21X1_585 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n71_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n90_));
AOI21X1 AOI21X1_586 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n75_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n86_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n92_));
AOI21X1 AOI21X1_587 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n91_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n93_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_));
AOI21X1 AOI21X1_588 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n115_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n117_));
AOI21X1 AOI21X1_589 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n122_));
AOI21X1 AOI21X1_59 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2686_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2687_));
AOI21X1 AOI21X1_590 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n157_));
AOI21X1 AOI21X1_591 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n175_));
AOI21X1 AOI21X1_592 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n231_));
AOI21X1 AOI21X1_593 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n181_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n240_));
AOI21X1 AOI21X1_594 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n237_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n212_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n270_));
AOI21X1 AOI21X1_595 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n245_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n226_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n271_));
AOI21X1 AOI21X1_596 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n149_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n293_));
AOI21X1 AOI21X1_597 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n302_));
AOI21X1 AOI21X1_598 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n307_));
AOI21X1 AOI21X1_599 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n303_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n301_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n311_));
AOI21X1 AOI21X1_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n146_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n148_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__0_));
AOI21X1 AOI21X1_60 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__29_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2692_));
AOI21X1 AOI21X1_600 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n295_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n312_));
AOI21X1 AOI21X1_601 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n65_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n387_));
AOI21X1 AOI21X1_602 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n395_));
AOI21X1 AOI21X1_603 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n445_));
AOI21X1 AOI21X1_604 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n446_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n447_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n448_));
AOI21X1 AOI21X1_605 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n435_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n450_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n451_));
AOI21X1 AOI21X1_61 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__30_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2698_));
AOI21X1 AOI21X1_62 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__31_), .C(AES_CORE_DATAPATH__abc_15863_new_n2468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2704_));
AOI21X1 AOI21X1_63 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2706_), .C(AES_CORE_DATAPATH__abc_15863_new_n2482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2707_));
AOI21X1 AOI21X1_64 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_out_sel_1_), .C(\key_sel_rd[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2720_));
AOI21X1 AOI21X1_65 ( .A(AES_CORE_CONTROL_UNIT_key_out_sel_0_), .B(AES_CORE_CONTROL_UNIT_bypass_key_en), .C(\key_sel_rd[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2727_));
AOI21X1 AOI21X1_66 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2733_), .B(AES_CORE_DATAPATH__abc_15863_new_n2712_), .C(AES_CORE_DATAPATH__abc_15863_new_n2734_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2735_));
AOI21X1 AOI21X1_67 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .B(AES_CORE_DATAPATH_last_round_pp2), .C(AES_CORE_DATAPATH__abc_15863_new_n3109_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3110_));
AOI21X1 AOI21X1_68 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .C(AES_CORE_DATAPATH__abc_15863_new_n3132_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3133_));
AOI21X1 AOI21X1_69 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .C(AES_CORE_DATAPATH__abc_15863_new_n3154_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3155_));
AOI21X1 AOI21X1_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n151_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n152_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__1_));
AOI21X1 AOI21X1_70 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .C(AES_CORE_DATAPATH__abc_15863_new_n3177_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3178_));
AOI21X1 AOI21X1_71 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n3199_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3200_));
AOI21X1 AOI21X1_72 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .C(AES_CORE_DATAPATH__abc_15863_new_n3221_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3222_));
AOI21X1 AOI21X1_73 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .C(AES_CORE_DATAPATH__abc_15863_new_n3243_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3244_));
AOI21X1 AOI21X1_74 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .C(AES_CORE_DATAPATH__abc_15863_new_n3265_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3266_));
AOI21X1 AOI21X1_75 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .C(AES_CORE_DATAPATH__abc_15863_new_n3287_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3288_));
AOI21X1 AOI21X1_76 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .C(AES_CORE_DATAPATH__abc_15863_new_n3309_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3310_));
AOI21X1 AOI21X1_77 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .C(AES_CORE_DATAPATH__abc_15863_new_n3331_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3332_));
AOI21X1 AOI21X1_78 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .C(AES_CORE_DATAPATH__abc_15863_new_n3353_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3354_));
AOI21X1 AOI21X1_79 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n3375_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3376_));
AOI21X1 AOI21X1_8 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n154_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n155_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__2_));
AOI21X1 AOI21X1_80 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .C(AES_CORE_DATAPATH__abc_15863_new_n3397_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3398_));
AOI21X1 AOI21X1_81 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .C(AES_CORE_DATAPATH__abc_15863_new_n3419_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3420_));
AOI21X1 AOI21X1_82 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .C(AES_CORE_DATAPATH__abc_15863_new_n3441_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3442_));
AOI21X1 AOI21X1_83 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .C(AES_CORE_DATAPATH__abc_15863_new_n3463_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3464_));
AOI21X1 AOI21X1_84 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .C(AES_CORE_DATAPATH__abc_15863_new_n3485_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3486_));
AOI21X1 AOI21X1_85 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .C(AES_CORE_DATAPATH__abc_15863_new_n3507_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3508_));
AOI21X1 AOI21X1_86 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .C(AES_CORE_DATAPATH__abc_15863_new_n3529_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3530_));
AOI21X1 AOI21X1_87 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n3551_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3552_));
AOI21X1 AOI21X1_88 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .C(AES_CORE_DATAPATH__abc_15863_new_n3573_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3574_));
AOI21X1 AOI21X1_89 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .C(AES_CORE_DATAPATH__abc_15863_new_n3595_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3596_));
AOI21X1 AOI21X1_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n172_), .B(AES_CORE_CONTROL_UNIT_state_6_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n171_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_));
AOI21X1 AOI21X1_90 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .C(AES_CORE_DATAPATH__abc_15863_new_n3617_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3618_));
AOI21X1 AOI21X1_91 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .C(AES_CORE_DATAPATH__abc_15863_new_n3639_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3640_));
AOI21X1 AOI21X1_92 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .C(AES_CORE_DATAPATH__abc_15863_new_n3661_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3662_));
AOI21X1 AOI21X1_93 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .C(AES_CORE_DATAPATH__abc_15863_new_n3683_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3684_));
AOI21X1 AOI21X1_94 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .C(AES_CORE_DATAPATH__abc_15863_new_n3705_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3706_));
AOI21X1 AOI21X1_95 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n3727_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3728_));
AOI21X1 AOI21X1_96 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .C(AES_CORE_DATAPATH__abc_15863_new_n3749_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3750_));
AOI21X1 AOI21X1_97 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .C(AES_CORE_DATAPATH__abc_15863_new_n3771_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3772_));
AOI21X1 AOI21X1_98 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .C(AES_CORE_DATAPATH__abc_15863_new_n3793_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3794_));
AOI21X1 AOI21X1_99 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2712_), .B(AES_CORE_DATAPATH_key_en_pp1_1_), .C(start), .Y(AES_CORE_DATAPATH__abc_15863_new_n3864_));
AOI22X1 AOI22X1_1 ( .A(AES_CORE_CONTROL_UNIT_rd_count_3_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n167_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n77_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n80_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n168_));
AOI22X1 AOI22X1_10 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3192_));
AOI22X1 AOI22X1_100 ( .A(AES_CORE_DATAPATH_bkp_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2482_), .C(AES_CORE_DATAPATH__abc_15863_new_n5450_), .D(AES_CORE_DATAPATH__abc_15863_new_n5452_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5453_));
AOI22X1 AOI22X1_101 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5456_), .D(AES_CORE_DATAPATH__abc_15863_new_n5462_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5466_));
AOI22X1 AOI22X1_102 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n5497_), .D(AES_CORE_DATAPATH__abc_15863_new_n5496_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5498_));
AOI22X1 AOI22X1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5493_), .D(AES_CORE_DATAPATH__abc_15863_new_n5501_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5505_));
AOI22X1 AOI22X1_104 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5534_), .D(AES_CORE_DATAPATH__abc_15863_new_n5540_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5544_));
AOI22X1 AOI22X1_105 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5558_), .D(AES_CORE_DATAPATH__abc_15863_new_n5557_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5559_));
AOI22X1 AOI22X1_106 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3663_), .D(AES_CORE_DATAPATH__abc_15863_new_n3659_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5575_));
AOI22X1 AOI22X1_107 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5574_), .D(AES_CORE_DATAPATH__abc_15863_new_n5578_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5582_));
AOI22X1 AOI22X1_108 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5597_), .D(AES_CORE_DATAPATH__abc_15863_new_n5596_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5598_));
AOI22X1 AOI22X1_109 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3685_), .D(AES_CORE_DATAPATH__abc_15863_new_n3681_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5614_));
AOI22X1 AOI22X1_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3196_), .D(AES_CORE_DATAPATH__abc_15863_new_n3194_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3197_));
AOI22X1 AOI22X1_110 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5613_), .D(AES_CORE_DATAPATH__abc_15863_new_n5617_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5621_));
AOI22X1 AOI22X1_111 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5651_), .D(AES_CORE_DATAPATH__abc_15863_new_n5657_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5661_));
AOI22X1 AOI22X1_112 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5675_), .D(AES_CORE_DATAPATH__abc_15863_new_n5674_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5676_));
AOI22X1 AOI22X1_113 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3729_), .D(AES_CORE_DATAPATH__abc_15863_new_n3725_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5692_));
AOI22X1 AOI22X1_114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5691_), .D(AES_CORE_DATAPATH__abc_15863_new_n5695_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5699_));
AOI22X1 AOI22X1_115 ( .A(AES_CORE_DATAPATH_bkp_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2482_), .C(AES_CORE_DATAPATH__abc_15863_new_n5720_), .D(AES_CORE_DATAPATH__abc_15863_new_n5722_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5723_));
AOI22X1 AOI22X1_116 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5726_), .D(AES_CORE_DATAPATH__abc_15863_new_n5732_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5736_));
AOI22X1 AOI22X1_117 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5765_), .D(AES_CORE_DATAPATH__abc_15863_new_n5771_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5775_));
AOI22X1 AOI22X1_118 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5789_), .D(AES_CORE_DATAPATH__abc_15863_new_n5788_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5790_));
AOI22X1 AOI22X1_119 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3795_), .D(AES_CORE_DATAPATH__abc_15863_new_n3791_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5806_));
AOI22X1 AOI22X1_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3214_));
AOI22X1 AOI22X1_120 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5805_), .D(AES_CORE_DATAPATH__abc_15863_new_n5809_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5813_));
AOI22X1 AOI22X1_121 ( .A(AES_CORE_DATAPATH_col_en_host_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n6709_), .C(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .D(AES_CORE_DATAPATH__abc_15863_new_n6712_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6713_));
AOI22X1 AOI22X1_122 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4605_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6783_), .D(AES_CORE_DATAPATH__abc_15863_new_n6781_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__0_));
AOI22X1 AOI22X1_123 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4646_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6789_), .D(AES_CORE_DATAPATH__abc_15863_new_n6787_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__1_));
AOI22X1 AOI22X1_124 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4687_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6795_), .D(AES_CORE_DATAPATH__abc_15863_new_n6793_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__2_));
AOI22X1 AOI22X1_125 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4727_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6801_), .D(AES_CORE_DATAPATH__abc_15863_new_n6799_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__3_));
AOI22X1 AOI22X1_126 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6803_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6808_), .D(AES_CORE_DATAPATH__abc_15863_new_n6806_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__4_));
AOI22X1 AOI22X1_127 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4802_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6814_), .D(AES_CORE_DATAPATH__abc_15863_new_n6812_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__5_));
AOI22X1 AOI22X1_128 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6816_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6821_), .D(AES_CORE_DATAPATH__abc_15863_new_n6819_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__6_));
AOI22X1 AOI22X1_129 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4874_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6827_), .D(AES_CORE_DATAPATH__abc_15863_new_n6825_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__7_));
AOI22X1 AOI22X1_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3218_), .D(AES_CORE_DATAPATH__abc_15863_new_n3216_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3219_));
AOI22X1 AOI22X1_130 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6829_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6834_), .D(AES_CORE_DATAPATH__abc_15863_new_n6832_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__8_));
AOI22X1 AOI22X1_131 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4951_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6840_), .D(AES_CORE_DATAPATH__abc_15863_new_n6838_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__9_));
AOI22X1 AOI22X1_132 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4989_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6846_), .D(AES_CORE_DATAPATH__abc_15863_new_n6844_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__10_));
AOI22X1 AOI22X1_133 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5029_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6852_), .D(AES_CORE_DATAPATH__abc_15863_new_n6850_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__11_));
AOI22X1 AOI22X1_134 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5067_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6858_), .D(AES_CORE_DATAPATH__abc_15863_new_n6856_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__12_));
AOI22X1 AOI22X1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5107_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6864_), .D(AES_CORE_DATAPATH__abc_15863_new_n6862_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__13_));
AOI22X1 AOI22X1_136 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6866_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6871_), .D(AES_CORE_DATAPATH__abc_15863_new_n6869_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__14_));
AOI22X1 AOI22X1_137 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5182_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6877_), .D(AES_CORE_DATAPATH__abc_15863_new_n6875_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__15_));
AOI22X1 AOI22X1_138 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5220_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6883_), .D(AES_CORE_DATAPATH__abc_15863_new_n6881_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__16_));
AOI22X1 AOI22X1_139 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5260_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6889_), .D(AES_CORE_DATAPATH__abc_15863_new_n6887_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__17_));
AOI22X1 AOI22X1_14 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3236_));
AOI22X1 AOI22X1_140 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5299_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6895_), .D(AES_CORE_DATAPATH__abc_15863_new_n6893_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__18_));
AOI22X1 AOI22X1_141 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5338_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6901_), .D(AES_CORE_DATAPATH__abc_15863_new_n6899_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__19_));
AOI22X1 AOI22X1_142 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5376_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6907_), .D(AES_CORE_DATAPATH__abc_15863_new_n6905_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__20_));
AOI22X1 AOI22X1_143 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5416_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6913_), .D(AES_CORE_DATAPATH__abc_15863_new_n6911_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__21_));
AOI22X1 AOI22X1_144 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6915_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6920_), .D(AES_CORE_DATAPATH__abc_15863_new_n6918_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__22_));
AOI22X1 AOI22X1_145 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5488_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6926_), .D(AES_CORE_DATAPATH__abc_15863_new_n6924_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__23_));
AOI22X1 AOI22X1_146 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5529_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6932_), .D(AES_CORE_DATAPATH__abc_15863_new_n6930_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__24_));
AOI22X1 AOI22X1_147 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5569_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6938_), .D(AES_CORE_DATAPATH__abc_15863_new_n6936_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__25_));
AOI22X1 AOI22X1_148 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5608_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6944_), .D(AES_CORE_DATAPATH__abc_15863_new_n6942_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__26_));
AOI22X1 AOI22X1_149 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5646_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6950_), .D(AES_CORE_DATAPATH__abc_15863_new_n6948_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__27_));
AOI22X1 AOI22X1_15 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3240_), .D(AES_CORE_DATAPATH__abc_15863_new_n3238_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3241_));
AOI22X1 AOI22X1_150 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5686_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6956_), .D(AES_CORE_DATAPATH__abc_15863_new_n6954_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__28_));
AOI22X1 AOI22X1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6958_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6963_), .D(AES_CORE_DATAPATH__abc_15863_new_n6961_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__29_));
AOI22X1 AOI22X1_152 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5760_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6969_), .D(AES_CORE_DATAPATH__abc_15863_new_n6967_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__30_));
AOI22X1 AOI22X1_153 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5800_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .C(AES_CORE_DATAPATH__abc_15863_new_n6975_), .D(AES_CORE_DATAPATH__abc_15863_new_n6973_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__31_));
AOI22X1 AOI22X1_154 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6980_), .B(AES_CORE_DATAPATH__abc_15863_new_n2457_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .D(AES_CORE_DATAPATH__abc_15863_new_n6983_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__0_));
AOI22X1 AOI22X1_155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2486_), .B(AES_CORE_DATAPATH__abc_15863_new_n6991_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .D(AES_CORE_DATAPATH__abc_15863_new_n6989_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__1_));
AOI22X1 AOI22X1_156 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2494_), .B(AES_CORE_DATAPATH__abc_15863_new_n6994_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .D(AES_CORE_DATAPATH__abc_15863_new_n6997_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__2_));
AOI22X1 AOI22X1_157 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2500_), .B(AES_CORE_DATAPATH__abc_15863_new_n6999_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .D(AES_CORE_DATAPATH__abc_15863_new_n7005_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__3_));
AOI22X1 AOI22X1_158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2508_), .B(AES_CORE_DATAPATH__abc_15863_new_n7007_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .D(AES_CORE_DATAPATH__abc_15863_new_n7011_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__4_));
AOI22X1 AOI22X1_159 ( .A(\bus_in[7] ), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .C(AES_CORE_DATAPATH__abc_15863_new_n7027_), .D(AES_CORE_DATAPATH__abc_15863_new_n7030_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7031_));
AOI22X1 AOI22X1_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3258_));
AOI22X1 AOI22X1_160 ( .A(\bus_in[8] ), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .C(AES_CORE_DATAPATH__abc_15863_new_n7029_), .D(AES_CORE_DATAPATH__abc_15863_new_n7035_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7036_));
AOI22X1 AOI22X1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2544_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7045_), .D(AES_CORE_DATAPATH__abc_15863_new_n7044_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__9_));
AOI22X1 AOI22X1_162 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2552_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7052_), .D(AES_CORE_DATAPATH__abc_15863_new_n7051_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__10_));
AOI22X1 AOI22X1_163 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2560_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7058_), .D(AES_CORE_DATAPATH__abc_15863_new_n7057_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__11_));
AOI22X1 AOI22X1_164 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2568_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7064_), .D(AES_CORE_DATAPATH__abc_15863_new_n7062_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__12_));
AOI22X1 AOI22X1_165 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2574_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7069_), .D(AES_CORE_DATAPATH__abc_15863_new_n7067_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__13_));
AOI22X1 AOI22X1_166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2582_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7076_), .D(AES_CORE_DATAPATH__abc_15863_new_n7074_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__14_));
AOI22X1 AOI22X1_167 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2588_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7082_), .D(AES_CORE_DATAPATH__abc_15863_new_n7080_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__15_));
AOI22X1 AOI22X1_168 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2596_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7089_), .D(AES_CORE_DATAPATH__abc_15863_new_n7087_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__16_));
AOI22X1 AOI22X1_169 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2602_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7094_), .D(AES_CORE_DATAPATH__abc_15863_new_n7092_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__17_));
AOI22X1 AOI22X1_17 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3262_), .D(AES_CORE_DATAPATH__abc_15863_new_n3260_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3263_));
AOI22X1 AOI22X1_170 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2610_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7100_), .D(AES_CORE_DATAPATH__abc_15863_new_n7098_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__18_));
AOI22X1 AOI22X1_171 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2618_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7105_), .D(AES_CORE_DATAPATH__abc_15863_new_n7103_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__19_));
AOI22X1 AOI22X1_172 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2626_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7121_), .D(AES_CORE_DATAPATH__abc_15863_new_n7119_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__20_));
AOI22X1 AOI22X1_173 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2632_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7128_), .D(AES_CORE_DATAPATH__abc_15863_new_n7126_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__21_));
AOI22X1 AOI22X1_174 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2640_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7136_), .D(AES_CORE_DATAPATH__abc_15863_new_n7134_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__22_));
AOI22X1 AOI22X1_175 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2646_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7143_), .D(AES_CORE_DATAPATH__abc_15863_new_n7141_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__23_));
AOI22X1 AOI22X1_176 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2654_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7154_), .D(AES_CORE_DATAPATH__abc_15863_new_n7152_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__24_));
AOI22X1 AOI22X1_177 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2660_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7161_), .D(AES_CORE_DATAPATH__abc_15863_new_n7159_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__25_));
AOI22X1 AOI22X1_178 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2668_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7170_), .D(AES_CORE_DATAPATH__abc_15863_new_n7168_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__26_));
AOI22X1 AOI22X1_179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2676_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7177_), .D(AES_CORE_DATAPATH__abc_15863_new_n7175_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__27_));
AOI22X1 AOI22X1_18 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3280_));
AOI22X1 AOI22X1_180 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2682_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7186_), .D(AES_CORE_DATAPATH__abc_15863_new_n7184_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__28_));
AOI22X1 AOI22X1_181 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2690_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7193_), .D(AES_CORE_DATAPATH__abc_15863_new_n7191_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__29_));
AOI22X1 AOI22X1_182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2696_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7201_), .D(AES_CORE_DATAPATH__abc_15863_new_n7199_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__30_));
AOI22X1 AOI22X1_183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2702_), .B(AES_CORE_DATAPATH__abc_15863_new_n6977_), .C(AES_CORE_DATAPATH__abc_15863_new_n7208_), .D(AES_CORE_DATAPATH__abc_15863_new_n7206_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__31_));
AOI22X1 AOI22X1_184 ( .A(AES_CORE_DATAPATH_col_en_host_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n6709_), .C(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .D(AES_CORE_DATAPATH__abc_15863_new_n6712_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7274_));
AOI22X1 AOI22X1_185 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4599_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7342_), .D(AES_CORE_DATAPATH__abc_15863_new_n7341_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__0_));
AOI22X1 AOI22X1_186 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4640_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7347_), .D(AES_CORE_DATAPATH__abc_15863_new_n7346_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__1_));
AOI22X1 AOI22X1_187 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4681_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7352_), .D(AES_CORE_DATAPATH__abc_15863_new_n7351_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__2_));
AOI22X1 AOI22X1_188 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4721_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7357_), .D(AES_CORE_DATAPATH__abc_15863_new_n7356_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__3_));
AOI22X1 AOI22X1_189 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4763_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7362_), .D(AES_CORE_DATAPATH__abc_15863_new_n7361_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__4_));
AOI22X1 AOI22X1_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3284_), .D(AES_CORE_DATAPATH__abc_15863_new_n3282_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3285_));
AOI22X1 AOI22X1_190 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4796_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7367_), .D(AES_CORE_DATAPATH__abc_15863_new_n7366_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__5_));
AOI22X1 AOI22X1_191 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4838_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7372_), .D(AES_CORE_DATAPATH__abc_15863_new_n7371_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__6_));
AOI22X1 AOI22X1_192 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4868_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7377_), .D(AES_CORE_DATAPATH__abc_15863_new_n7376_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__7_));
AOI22X1 AOI22X1_193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4912_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7382_), .D(AES_CORE_DATAPATH__abc_15863_new_n7381_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__8_));
AOI22X1 AOI22X1_194 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4945_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7387_), .D(AES_CORE_DATAPATH__abc_15863_new_n7386_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__9_));
AOI22X1 AOI22X1_195 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4983_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7392_), .D(AES_CORE_DATAPATH__abc_15863_new_n7391_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__10_));
AOI22X1 AOI22X1_196 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5023_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7397_), .D(AES_CORE_DATAPATH__abc_15863_new_n7396_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__11_));
AOI22X1 AOI22X1_197 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5061_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7402_), .D(AES_CORE_DATAPATH__abc_15863_new_n7401_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__12_));
AOI22X1 AOI22X1_198 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5101_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7407_), .D(AES_CORE_DATAPATH__abc_15863_new_n7406_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__13_));
AOI22X1 AOI22X1_199 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5142_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7412_), .D(AES_CORE_DATAPATH__abc_15863_new_n7411_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__14_));
AOI22X1 AOI22X1_2 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_CONTROL_UNIT_last_round), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n182_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n183_));
AOI22X1 AOI22X1_20 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3302_));
AOI22X1 AOI22X1_200 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5176_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7417_), .D(AES_CORE_DATAPATH__abc_15863_new_n7416_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__15_));
AOI22X1 AOI22X1_201 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5214_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7422_), .D(AES_CORE_DATAPATH__abc_15863_new_n7421_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__16_));
AOI22X1 AOI22X1_202 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5254_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7427_), .D(AES_CORE_DATAPATH__abc_15863_new_n7426_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__17_));
AOI22X1 AOI22X1_203 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5293_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7432_), .D(AES_CORE_DATAPATH__abc_15863_new_n7431_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__18_));
AOI22X1 AOI22X1_204 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5332_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7437_), .D(AES_CORE_DATAPATH__abc_15863_new_n7436_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__19_));
AOI22X1 AOI22X1_205 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5370_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7442_), .D(AES_CORE_DATAPATH__abc_15863_new_n7441_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__20_));
AOI22X1 AOI22X1_206 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5410_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7447_), .D(AES_CORE_DATAPATH__abc_15863_new_n7446_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__21_));
AOI22X1 AOI22X1_207 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5451_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7452_), .D(AES_CORE_DATAPATH__abc_15863_new_n7451_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__22_));
AOI22X1 AOI22X1_208 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5482_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7457_), .D(AES_CORE_DATAPATH__abc_15863_new_n7456_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__23_));
AOI22X1 AOI22X1_209 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5523_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7462_), .D(AES_CORE_DATAPATH__abc_15863_new_n7461_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__24_));
AOI22X1 AOI22X1_21 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3324_));
AOI22X1 AOI22X1_210 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5563_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7467_), .D(AES_CORE_DATAPATH__abc_15863_new_n7466_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__25_));
AOI22X1 AOI22X1_211 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5602_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7472_), .D(AES_CORE_DATAPATH__abc_15863_new_n7471_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__26_));
AOI22X1 AOI22X1_212 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5640_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7477_), .D(AES_CORE_DATAPATH__abc_15863_new_n7476_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__27_));
AOI22X1 AOI22X1_213 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5680_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7482_), .D(AES_CORE_DATAPATH__abc_15863_new_n7481_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__28_));
AOI22X1 AOI22X1_214 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5721_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7487_), .D(AES_CORE_DATAPATH__abc_15863_new_n7486_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__29_));
AOI22X1 AOI22X1_215 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5754_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7492_), .D(AES_CORE_DATAPATH__abc_15863_new_n7491_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__30_));
AOI22X1 AOI22X1_216 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5794_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .C(AES_CORE_DATAPATH__abc_15863_new_n7497_), .D(AES_CORE_DATAPATH__abc_15863_new_n7496_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__31_));
AOI22X1 AOI22X1_217 ( .A(AES_CORE_DATAPATH_col_en_host_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n6709_), .C(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .D(AES_CORE_DATAPATH__abc_15863_new_n6712_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7563_));
AOI22X1 AOI22X1_218 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7644_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7648_), .D(AES_CORE_DATAPATH__abc_15863_new_n7647_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__0_));
AOI22X1 AOI22X1_219 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7650_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7653_), .D(AES_CORE_DATAPATH__abc_15863_new_n7652_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__1_));
AOI22X1 AOI22X1_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3328_), .D(AES_CORE_DATAPATH__abc_15863_new_n3326_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3329_));
AOI22X1 AOI22X1_220 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7655_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7659_), .D(AES_CORE_DATAPATH__abc_15863_new_n7658_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__2_));
AOI22X1 AOI22X1_221 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7661_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7664_), .D(AES_CORE_DATAPATH__abc_15863_new_n7663_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__3_));
AOI22X1 AOI22X1_222 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7666_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7670_), .D(AES_CORE_DATAPATH__abc_15863_new_n7669_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__4_));
AOI22X1 AOI22X1_223 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7672_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7676_), .D(AES_CORE_DATAPATH__abc_15863_new_n7675_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__5_));
AOI22X1 AOI22X1_224 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7678_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7682_), .D(AES_CORE_DATAPATH__abc_15863_new_n7681_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__6_));
AOI22X1 AOI22X1_225 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7684_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7687_), .D(AES_CORE_DATAPATH__abc_15863_new_n7686_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__7_));
AOI22X1 AOI22X1_226 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7689_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7693_), .D(AES_CORE_DATAPATH__abc_15863_new_n7692_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__8_));
AOI22X1 AOI22X1_227 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7695_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7698_), .D(AES_CORE_DATAPATH__abc_15863_new_n7697_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__9_));
AOI22X1 AOI22X1_228 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7700_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7704_), .D(AES_CORE_DATAPATH__abc_15863_new_n7703_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__10_));
AOI22X1 AOI22X1_229 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7706_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7709_), .D(AES_CORE_DATAPATH__abc_15863_new_n7708_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__11_));
AOI22X1 AOI22X1_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3346_));
AOI22X1 AOI22X1_230 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7711_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7715_), .D(AES_CORE_DATAPATH__abc_15863_new_n7714_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__12_));
AOI22X1 AOI22X1_231 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7717_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7720_), .D(AES_CORE_DATAPATH__abc_15863_new_n7719_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__13_));
AOI22X1 AOI22X1_232 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7722_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7726_), .D(AES_CORE_DATAPATH__abc_15863_new_n7725_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__14_));
AOI22X1 AOI22X1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7728_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7731_), .D(AES_CORE_DATAPATH__abc_15863_new_n7730_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__15_));
AOI22X1 AOI22X1_234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7733_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7737_), .D(AES_CORE_DATAPATH__abc_15863_new_n7736_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__16_));
AOI22X1 AOI22X1_235 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7739_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7742_), .D(AES_CORE_DATAPATH__abc_15863_new_n7741_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__17_));
AOI22X1 AOI22X1_236 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7744_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7747_), .D(AES_CORE_DATAPATH__abc_15863_new_n7746_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__18_));
AOI22X1 AOI22X1_237 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7749_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7752_), .D(AES_CORE_DATAPATH__abc_15863_new_n7751_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__19_));
AOI22X1 AOI22X1_238 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7754_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7758_), .D(AES_CORE_DATAPATH__abc_15863_new_n7757_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__20_));
AOI22X1 AOI22X1_239 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7760_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7763_), .D(AES_CORE_DATAPATH__abc_15863_new_n7762_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__21_));
AOI22X1 AOI22X1_24 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3368_));
AOI22X1 AOI22X1_240 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7765_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7769_), .D(AES_CORE_DATAPATH__abc_15863_new_n7768_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__22_));
AOI22X1 AOI22X1_241 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7771_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7774_), .D(AES_CORE_DATAPATH__abc_15863_new_n7773_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__23_));
AOI22X1 AOI22X1_242 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7776_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7780_), .D(AES_CORE_DATAPATH__abc_15863_new_n7779_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__24_));
AOI22X1 AOI22X1_243 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7782_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7785_), .D(AES_CORE_DATAPATH__abc_15863_new_n7784_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__25_));
AOI22X1 AOI22X1_244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7787_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7790_), .D(AES_CORE_DATAPATH__abc_15863_new_n7789_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__26_));
AOI22X1 AOI22X1_245 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7792_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7796_), .D(AES_CORE_DATAPATH__abc_15863_new_n7795_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__27_));
AOI22X1 AOI22X1_246 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7798_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7801_), .D(AES_CORE_DATAPATH__abc_15863_new_n7800_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__28_));
AOI22X1 AOI22X1_247 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7803_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7807_), .D(AES_CORE_DATAPATH__abc_15863_new_n7806_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__29_));
AOI22X1 AOI22X1_248 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7809_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7813_), .D(AES_CORE_DATAPATH__abc_15863_new_n7812_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__30_));
AOI22X1 AOI22X1_249 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7815_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7818_), .D(AES_CORE_DATAPATH__abc_15863_new_n7817_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__31_));
AOI22X1 AOI22X1_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3372_), .D(AES_CORE_DATAPATH__abc_15863_new_n3370_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3373_));
AOI22X1 AOI22X1_250 ( .A(AES_CORE_DATAPATH_col_en_host_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n6709_), .C(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .D(AES_CORE_DATAPATH__abc_15863_new_n6712_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7890_));
AOI22X1 AOI22X1_251 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7955_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7959_), .D(AES_CORE_DATAPATH__abc_15863_new_n7958_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__0_));
AOI22X1 AOI22X1_252 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7961_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7965_), .D(AES_CORE_DATAPATH__abc_15863_new_n7964_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__1_));
AOI22X1 AOI22X1_253 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7967_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7971_), .D(AES_CORE_DATAPATH__abc_15863_new_n7970_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__2_));
AOI22X1 AOI22X1_254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7973_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7977_), .D(AES_CORE_DATAPATH__abc_15863_new_n7976_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__3_));
AOI22X1 AOI22X1_255 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7979_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7983_), .D(AES_CORE_DATAPATH__abc_15863_new_n7982_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__4_));
AOI22X1 AOI22X1_256 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7985_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7989_), .D(AES_CORE_DATAPATH__abc_15863_new_n7988_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__5_));
AOI22X1 AOI22X1_257 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7991_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n7995_), .D(AES_CORE_DATAPATH__abc_15863_new_n7994_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__6_));
AOI22X1 AOI22X1_258 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7997_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8001_), .D(AES_CORE_DATAPATH__abc_15863_new_n8000_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__7_));
AOI22X1 AOI22X1_259 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8003_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8007_), .D(AES_CORE_DATAPATH__abc_15863_new_n8006_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__8_));
AOI22X1 AOI22X1_26 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3390_));
AOI22X1 AOI22X1_260 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8009_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8013_), .D(AES_CORE_DATAPATH__abc_15863_new_n8012_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__9_));
AOI22X1 AOI22X1_261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8015_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8019_), .D(AES_CORE_DATAPATH__abc_15863_new_n8018_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__10_));
AOI22X1 AOI22X1_262 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8021_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8025_), .D(AES_CORE_DATAPATH__abc_15863_new_n8024_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__11_));
AOI22X1 AOI22X1_263 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8027_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8031_), .D(AES_CORE_DATAPATH__abc_15863_new_n8030_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__12_));
AOI22X1 AOI22X1_264 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8033_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8037_), .D(AES_CORE_DATAPATH__abc_15863_new_n8036_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__13_));
AOI22X1 AOI22X1_265 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8039_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8043_), .D(AES_CORE_DATAPATH__abc_15863_new_n8042_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__14_));
AOI22X1 AOI22X1_266 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8045_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8049_), .D(AES_CORE_DATAPATH__abc_15863_new_n8048_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__15_));
AOI22X1 AOI22X1_267 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8051_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8055_), .D(AES_CORE_DATAPATH__abc_15863_new_n8054_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__16_));
AOI22X1 AOI22X1_268 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8057_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8061_), .D(AES_CORE_DATAPATH__abc_15863_new_n8060_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__17_));
AOI22X1 AOI22X1_269 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8063_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8067_), .D(AES_CORE_DATAPATH__abc_15863_new_n8066_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__18_));
AOI22X1 AOI22X1_27 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3412_));
AOI22X1 AOI22X1_270 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8069_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8073_), .D(AES_CORE_DATAPATH__abc_15863_new_n8072_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__19_));
AOI22X1 AOI22X1_271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8075_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8079_), .D(AES_CORE_DATAPATH__abc_15863_new_n8078_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__20_));
AOI22X1 AOI22X1_272 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8081_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8085_), .D(AES_CORE_DATAPATH__abc_15863_new_n8084_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__21_));
AOI22X1 AOI22X1_273 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8087_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8091_), .D(AES_CORE_DATAPATH__abc_15863_new_n8090_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__22_));
AOI22X1 AOI22X1_274 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8093_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8097_), .D(AES_CORE_DATAPATH__abc_15863_new_n8096_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__23_));
AOI22X1 AOI22X1_275 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8099_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8103_), .D(AES_CORE_DATAPATH__abc_15863_new_n8102_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__24_));
AOI22X1 AOI22X1_276 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8105_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8109_), .D(AES_CORE_DATAPATH__abc_15863_new_n8108_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__25_));
AOI22X1 AOI22X1_277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8111_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8115_), .D(AES_CORE_DATAPATH__abc_15863_new_n8114_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__26_));
AOI22X1 AOI22X1_278 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8117_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8121_), .D(AES_CORE_DATAPATH__abc_15863_new_n8120_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__27_));
AOI22X1 AOI22X1_279 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8123_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8127_), .D(AES_CORE_DATAPATH__abc_15863_new_n8126_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__28_));
AOI22X1 AOI22X1_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3416_), .D(AES_CORE_DATAPATH__abc_15863_new_n3414_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3417_));
AOI22X1 AOI22X1_280 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8129_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8133_), .D(AES_CORE_DATAPATH__abc_15863_new_n8132_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__29_));
AOI22X1 AOI22X1_281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8135_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8139_), .D(AES_CORE_DATAPATH__abc_15863_new_n8138_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__30_));
AOI22X1 AOI22X1_282 ( .A(AES_CORE_DATAPATH__abc_15863_new_n8141_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .C(AES_CORE_DATAPATH__abc_15863_new_n8145_), .D(AES_CORE_DATAPATH__abc_15863_new_n8144_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__31_));
AOI22X1 AOI22X1_283 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n441_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n478_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n415_), .D(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n477_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n479_));
AOI22X1 AOI22X1_284 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n101_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n102_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n129_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n131_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n132_));
AOI22X1 AOI22X1_285 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n135_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n136_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n133_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n134_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n137_));
AOI22X1 AOI22X1_286 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n133_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n134_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n129_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n131_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n148_));
AOI22X1 AOI22X1_287 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n101_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n102_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n135_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n136_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n149_));
AOI22X1 AOI22X1_288 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n253_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n257_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n245_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n246_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n258_));
AOI22X1 AOI22X1_289 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n267_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n268_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n269_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n270_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n271_));
AOI22X1 AOI22X1_29 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3434_));
AOI22X1 AOI22X1_290 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n272_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n255_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n172_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n173_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n273_));
AOI22X1 AOI22X1_291 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n295_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n297_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n314_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n315_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n318_));
AOI22X1 AOI22X1_292 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n311_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n312_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n309_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n319_));
AOI22X1 AOI22X1_293 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n253_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n257_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n225_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n226_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n386_));
AOI22X1 AOI22X1_294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n139_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n141_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_));
AOI22X1 AOI22X1_295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n139_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n147_));
AOI22X1 AOI22X1_296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n169_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n176_));
AOI22X1 AOI22X1_297 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n161_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n186_));
AOI22X1 AOI22X1_298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n155_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n187_));
AOI22X1 AOI22X1_299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n144_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n190_));
AOI22X1 AOI22X1_3 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3101_));
AOI22X1 AOI22X1_30 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3456_));
AOI22X1 AOI22X1_300 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n210_));
AOI22X1 AOI22X1_301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n249_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n181_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n250_));
AOI22X1 AOI22X1_302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n251_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n252_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n253_));
AOI22X1 AOI22X1_303 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n289_));
AOI22X1 AOI22X1_304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n291_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n292_));
AOI22X1 AOI22X1_305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n232_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n233_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n294_));
AOI22X1 AOI22X1_306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n229_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n304_));
AOI22X1 AOI22X1_307 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n290_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n309_));
AOI22X1 AOI22X1_308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n310_));
AOI22X1 AOI22X1_309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n330_));
AOI22X1 AOI22X1_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3460_), .D(AES_CORE_DATAPATH__abc_15863_new_n3458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3461_));
AOI22X1 AOI22X1_310 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n332_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n331_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n333_));
AOI22X1 AOI22X1_311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n331_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n332_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n335_));
AOI22X1 AOI22X1_312 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n336_));
AOI22X1 AOI22X1_313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n491_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n492_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n381_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n493_));
AOI22X1 AOI22X1_314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n494_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n495_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n377_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n496_));
AOI22X1 AOI22X1_315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n139_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n141_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_));
AOI22X1 AOI22X1_316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n139_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n147_));
AOI22X1 AOI22X1_317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n169_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n176_));
AOI22X1 AOI22X1_318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n161_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n186_));
AOI22X1 AOI22X1_319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n155_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n187_));
AOI22X1 AOI22X1_32 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3478_));
AOI22X1 AOI22X1_320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n144_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n190_));
AOI22X1 AOI22X1_321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n210_));
AOI22X1 AOI22X1_322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n249_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n181_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n250_));
AOI22X1 AOI22X1_323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n251_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n252_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n253_));
AOI22X1 AOI22X1_324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n289_));
AOI22X1 AOI22X1_325 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n291_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n292_));
AOI22X1 AOI22X1_326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n232_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n233_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n294_));
AOI22X1 AOI22X1_327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n229_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n304_));
AOI22X1 AOI22X1_328 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n290_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n309_));
AOI22X1 AOI22X1_329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n310_));
AOI22X1 AOI22X1_33 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3500_));
AOI22X1 AOI22X1_330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n330_));
AOI22X1 AOI22X1_331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n332_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n331_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n333_));
AOI22X1 AOI22X1_332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n331_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n332_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n335_));
AOI22X1 AOI22X1_333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n336_));
AOI22X1 AOI22X1_334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n491_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n492_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n381_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n493_));
AOI22X1 AOI22X1_335 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n494_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n495_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n377_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n496_));
AOI22X1 AOI22X1_336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n139_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n141_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_));
AOI22X1 AOI22X1_337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n139_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n147_));
AOI22X1 AOI22X1_338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n169_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n176_));
AOI22X1 AOI22X1_339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n161_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n186_));
AOI22X1 AOI22X1_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3522_));
AOI22X1 AOI22X1_340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n155_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n187_));
AOI22X1 AOI22X1_341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n144_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n190_));
AOI22X1 AOI22X1_342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n210_));
AOI22X1 AOI22X1_343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n249_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n181_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n250_));
AOI22X1 AOI22X1_344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n251_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n252_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n253_));
AOI22X1 AOI22X1_345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n289_));
AOI22X1 AOI22X1_346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n291_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n292_));
AOI22X1 AOI22X1_347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n232_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n233_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n294_));
AOI22X1 AOI22X1_348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n229_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n304_));
AOI22X1 AOI22X1_349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n290_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n309_));
AOI22X1 AOI22X1_35 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3544_));
AOI22X1 AOI22X1_350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n310_));
AOI22X1 AOI22X1_351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n330_));
AOI22X1 AOI22X1_352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n332_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n331_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n333_));
AOI22X1 AOI22X1_353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n331_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n332_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n335_));
AOI22X1 AOI22X1_354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n336_));
AOI22X1 AOI22X1_355 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n491_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n492_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n381_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n493_));
AOI22X1 AOI22X1_356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n494_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n495_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n377_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n496_));
AOI22X1 AOI22X1_357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n139_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n141_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_));
AOI22X1 AOI22X1_358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n139_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n147_));
AOI22X1 AOI22X1_359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n169_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n176_));
AOI22X1 AOI22X1_36 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3548_), .D(AES_CORE_DATAPATH__abc_15863_new_n3546_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3549_));
AOI22X1 AOI22X1_360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n161_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n186_));
AOI22X1 AOI22X1_361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n155_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n187_));
AOI22X1 AOI22X1_362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n144_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n190_));
AOI22X1 AOI22X1_363 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n210_));
AOI22X1 AOI22X1_364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n249_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n181_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n250_));
AOI22X1 AOI22X1_365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n251_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n252_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n253_));
AOI22X1 AOI22X1_366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n289_));
AOI22X1 AOI22X1_367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n291_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n292_));
AOI22X1 AOI22X1_368 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n232_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n233_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n294_));
AOI22X1 AOI22X1_369 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n229_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n304_));
AOI22X1 AOI22X1_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3566_));
AOI22X1 AOI22X1_370 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n290_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n284_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n309_));
AOI22X1 AOI22X1_371 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n285_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n288_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n179_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n310_));
AOI22X1 AOI22X1_372 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n330_));
AOI22X1 AOI22X1_373 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n332_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n331_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n333_));
AOI22X1 AOI22X1_374 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n331_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n332_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n303_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n305_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n335_));
AOI22X1 AOI22X1_375 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n329_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n295_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n336_));
AOI22X1 AOI22X1_376 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n491_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n492_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n381_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n493_));
AOI22X1 AOI22X1_377 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n494_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n495_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n377_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n496_));
AOI22X1 AOI22X1_378 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[0] ), .C(\bus_in[31] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n73_));
AOI22X1 AOI22X1_379 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[1] ), .C(\bus_in[30] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n77_));
AOI22X1 AOI22X1_38 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3588_));
AOI22X1 AOI22X1_380 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[2] ), .C(\bus_in[29] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n81_));
AOI22X1 AOI22X1_381 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[3] ), .C(\bus_in[28] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n85_));
AOI22X1 AOI22X1_382 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[4] ), .C(\bus_in[27] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n89_));
AOI22X1 AOI22X1_383 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[5] ), .C(\bus_in[26] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n93_));
AOI22X1 AOI22X1_384 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[6] ), .C(\bus_in[25] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n97_));
AOI22X1 AOI22X1_385 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[7] ), .C(\bus_in[24] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n101_));
AOI22X1 AOI22X1_386 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[8] ), .C(\bus_in[23] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n105_));
AOI22X1 AOI22X1_387 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[9] ), .C(\bus_in[22] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n109_));
AOI22X1 AOI22X1_388 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[10] ), .C(\bus_in[21] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n113_));
AOI22X1 AOI22X1_389 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[11] ), .C(\bus_in[20] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n117_));
AOI22X1 AOI22X1_39 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3592_), .D(AES_CORE_DATAPATH__abc_15863_new_n3590_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3593_));
AOI22X1 AOI22X1_390 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[12] ), .C(\bus_in[19] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n121_));
AOI22X1 AOI22X1_391 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[13] ), .C(\bus_in[18] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n125_));
AOI22X1 AOI22X1_392 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[14] ), .C(\bus_in[17] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n129_));
AOI22X1 AOI22X1_393 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[15] ), .C(\bus_in[16] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n133_));
AOI22X1 AOI22X1_394 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[16] ), .C(\bus_in[15] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n137_));
AOI22X1 AOI22X1_395 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[17] ), .C(\bus_in[14] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n141_));
AOI22X1 AOI22X1_396 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[18] ), .C(\bus_in[13] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n145_));
AOI22X1 AOI22X1_397 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[19] ), .C(\bus_in[12] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n149_));
AOI22X1 AOI22X1_398 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[20] ), .C(\bus_in[11] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n153_));
AOI22X1 AOI22X1_399 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[21] ), .C(\bus_in[10] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n157_));
AOI22X1 AOI22X1_4 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3105_), .D(AES_CORE_DATAPATH__abc_15863_new_n3103_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3106_));
AOI22X1 AOI22X1_40 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3610_));
AOI22X1 AOI22X1_400 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[22] ), .C(\bus_in[9] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n161_));
AOI22X1 AOI22X1_401 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[23] ), .C(\bus_in[8] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n165_));
AOI22X1 AOI22X1_402 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[24] ), .C(\bus_in[7] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n169_));
AOI22X1 AOI22X1_403 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[25] ), .C(\bus_in[6] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n173_));
AOI22X1 AOI22X1_404 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[26] ), .C(\bus_in[5] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n177_));
AOI22X1 AOI22X1_405 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[27] ), .C(\bus_in[4] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n181_));
AOI22X1 AOI22X1_406 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[28] ), .C(\bus_in[3] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n185_));
AOI22X1 AOI22X1_407 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[29] ), .C(\bus_in[2] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n189_));
AOI22X1 AOI22X1_408 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[30] ), .C(\bus_in[1] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n193_));
AOI22X1 AOI22X1_409 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_), .B(\bus_in[31] ), .C(\bus_in[0] ), .D(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n197_));
AOI22X1 AOI22X1_41 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3614_), .D(AES_CORE_DATAPATH__abc_15863_new_n3612_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3615_));
AOI22X1 AOI22X1_410 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n73_));
AOI22X1 AOI22X1_411 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n77_));
AOI22X1 AOI22X1_412 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n81_));
AOI22X1 AOI22X1_413 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n85_));
AOI22X1 AOI22X1_414 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n89_));
AOI22X1 AOI22X1_415 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n93_));
AOI22X1 AOI22X1_416 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n97_));
AOI22X1 AOI22X1_417 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n101_));
AOI22X1 AOI22X1_418 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n105_));
AOI22X1 AOI22X1_419 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n109_));
AOI22X1 AOI22X1_42 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3632_));
AOI22X1 AOI22X1_420 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n113_));
AOI22X1 AOI22X1_421 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n117_));
AOI22X1 AOI22X1_422 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n121_));
AOI22X1 AOI22X1_423 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n125_));
AOI22X1 AOI22X1_424 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n129_));
AOI22X1 AOI22X1_425 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n133_));
AOI22X1 AOI22X1_426 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n137_));
AOI22X1 AOI22X1_427 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n141_));
AOI22X1 AOI22X1_428 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n145_));
AOI22X1 AOI22X1_429 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n149_));
AOI22X1 AOI22X1_43 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3636_), .D(AES_CORE_DATAPATH__abc_15863_new_n3634_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3637_));
AOI22X1 AOI22X1_430 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n153_));
AOI22X1 AOI22X1_431 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n157_));
AOI22X1 AOI22X1_432 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n161_));
AOI22X1 AOI22X1_433 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n165_));
AOI22X1 AOI22X1_434 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n169_));
AOI22X1 AOI22X1_435 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n173_));
AOI22X1 AOI22X1_436 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n177_));
AOI22X1 AOI22X1_437 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n181_));
AOI22X1 AOI22X1_438 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n185_));
AOI22X1 AOI22X1_439 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n189_));
AOI22X1 AOI22X1_44 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3654_));
AOI22X1 AOI22X1_440 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n193_));
AOI22X1 AOI22X1_441 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .D(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n197_));
AOI22X1 AOI22X1_45 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3676_));
AOI22X1 AOI22X1_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3698_));
AOI22X1 AOI22X1_47 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3702_), .D(AES_CORE_DATAPATH__abc_15863_new_n3700_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3703_));
AOI22X1 AOI22X1_48 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3720_));
AOI22X1 AOI22X1_49 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3742_));
AOI22X1 AOI22X1_5 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3125_));
AOI22X1 AOI22X1_50 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3746_), .D(AES_CORE_DATAPATH__abc_15863_new_n3744_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3747_));
AOI22X1 AOI22X1_51 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3764_));
AOI22X1 AOI22X1_52 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3768_), .D(AES_CORE_DATAPATH__abc_15863_new_n3766_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3769_));
AOI22X1 AOI22X1_53 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3786_));
AOI22X1 AOI22X1_54 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4610_), .D(AES_CORE_DATAPATH__abc_15863_new_n4616_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4622_));
AOI22X1 AOI22X1_55 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n4655_), .D(AES_CORE_DATAPATH__abc_15863_new_n4654_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4656_));
AOI22X1 AOI22X1_56 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4651_), .D(AES_CORE_DATAPATH__abc_15863_new_n4659_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4663_));
AOI22X1 AOI22X1_57 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4692_), .D(AES_CORE_DATAPATH__abc_15863_new_n4698_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4702_));
AOI22X1 AOI22X1_58 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n4716_), .D(AES_CORE_DATAPATH__abc_15863_new_n4715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4717_));
AOI22X1 AOI22X1_59 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3179_), .D(AES_CORE_DATAPATH__abc_15863_new_n3175_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4733_));
AOI22X1 AOI22X1_6 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3129_), .D(AES_CORE_DATAPATH__abc_15863_new_n3127_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3130_));
AOI22X1 AOI22X1_60 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4732_), .D(AES_CORE_DATAPATH__abc_15863_new_n4736_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4740_));
AOI22X1 AOI22X1_61 ( .A(AES_CORE_DATAPATH_bkp_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2482_), .C(AES_CORE_DATAPATH__abc_15863_new_n4762_), .D(AES_CORE_DATAPATH__abc_15863_new_n4764_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4765_));
AOI22X1 AOI22X1_62 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4768_), .D(AES_CORE_DATAPATH__abc_15863_new_n4774_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4778_));
AOI22X1 AOI22X1_63 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4807_), .D(AES_CORE_DATAPATH__abc_15863_new_n4813_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4817_));
AOI22X1 AOI22X1_64 ( .A(AES_CORE_DATAPATH_bkp_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n2482_), .C(AES_CORE_DATAPATH__abc_15863_new_n4837_), .D(AES_CORE_DATAPATH__abc_15863_new_n4839_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4840_));
AOI22X1 AOI22X1_65 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4843_), .D(AES_CORE_DATAPATH__abc_15863_new_n4848_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4852_));
AOI22X1 AOI22X1_66 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n4883_), .D(AES_CORE_DATAPATH__abc_15863_new_n4882_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4884_));
AOI22X1 AOI22X1_67 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4879_), .D(AES_CORE_DATAPATH__abc_15863_new_n4887_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4891_));
AOI22X1 AOI22X1_68 ( .A(AES_CORE_DATAPATH_bkp_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n2482_), .C(AES_CORE_DATAPATH__abc_15863_new_n4911_), .D(AES_CORE_DATAPATH__abc_15863_new_n4913_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4914_));
AOI22X1 AOI22X1_69 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4917_), .D(AES_CORE_DATAPATH__abc_15863_new_n4922_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4926_));
AOI22X1 AOI22X1_7 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3147_));
AOI22X1 AOI22X1_70 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n4940_), .D(AES_CORE_DATAPATH__abc_15863_new_n4939_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4941_));
AOI22X1 AOI22X1_71 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3311_), .D(AES_CORE_DATAPATH__abc_15863_new_n3307_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4957_));
AOI22X1 AOI22X1_72 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4956_), .D(AES_CORE_DATAPATH__abc_15863_new_n4960_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4964_));
AOI22X1 AOI22X1_73 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n4994_), .D(AES_CORE_DATAPATH__abc_15863_new_n5000_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5004_));
AOI22X1 AOI22X1_74 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5018_), .D(AES_CORE_DATAPATH__abc_15863_new_n5017_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5019_));
AOI22X1 AOI22X1_75 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3355_), .D(AES_CORE_DATAPATH__abc_15863_new_n3351_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5035_));
AOI22X1 AOI22X1_76 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5034_), .D(AES_CORE_DATAPATH__abc_15863_new_n5038_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5042_));
AOI22X1 AOI22X1_77 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5072_), .D(AES_CORE_DATAPATH__abc_15863_new_n5078_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5082_));
AOI22X1 AOI22X1_78 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5096_), .D(AES_CORE_DATAPATH__abc_15863_new_n5095_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5097_));
AOI22X1 AOI22X1_79 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3399_), .D(AES_CORE_DATAPATH__abc_15863_new_n3395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5113_));
AOI22X1 AOI22X1_8 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n3151_), .D(AES_CORE_DATAPATH__abc_15863_new_n3149_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3152_));
AOI22X1 AOI22X1_80 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5112_), .D(AES_CORE_DATAPATH__abc_15863_new_n5116_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5120_));
AOI22X1 AOI22X1_81 ( .A(AES_CORE_DATAPATH_bkp_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2482_), .C(AES_CORE_DATAPATH__abc_15863_new_n5141_), .D(AES_CORE_DATAPATH__abc_15863_new_n5143_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5144_));
AOI22X1 AOI22X1_82 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5147_), .D(AES_CORE_DATAPATH__abc_15863_new_n5153_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5157_));
AOI22X1 AOI22X1_83 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5171_), .D(AES_CORE_DATAPATH__abc_15863_new_n5170_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5172_));
AOI22X1 AOI22X1_84 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3443_), .D(AES_CORE_DATAPATH__abc_15863_new_n3439_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5188_));
AOI22X1 AOI22X1_85 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5187_), .D(AES_CORE_DATAPATH__abc_15863_new_n5191_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5195_));
AOI22X1 AOI22X1_86 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5225_), .D(AES_CORE_DATAPATH__abc_15863_new_n5231_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5235_));
AOI22X1 AOI22X1_87 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5249_), .D(AES_CORE_DATAPATH__abc_15863_new_n5248_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5250_));
AOI22X1 AOI22X1_88 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3487_), .D(AES_CORE_DATAPATH__abc_15863_new_n3483_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5266_));
AOI22X1 AOI22X1_89 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5265_), .D(AES_CORE_DATAPATH__abc_15863_new_n5269_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5273_));
AOI22X1 AOI22X1_9 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3100_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_), .D(AES_CORE_DATAPATH__abc_15863_new_n3099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3170_));
AOI22X1 AOI22X1_90 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5288_), .D(AES_CORE_DATAPATH__abc_15863_new_n5287_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5289_));
AOI22X1 AOI22X1_91 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3509_), .D(AES_CORE_DATAPATH__abc_15863_new_n3505_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5305_));
AOI22X1 AOI22X1_92 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5304_), .D(AES_CORE_DATAPATH__abc_15863_new_n5308_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5312_));
AOI22X1 AOI22X1_93 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5327_), .D(AES_CORE_DATAPATH__abc_15863_new_n5326_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5328_));
AOI22X1 AOI22X1_94 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3531_), .D(AES_CORE_DATAPATH__abc_15863_new_n3527_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5344_));
AOI22X1 AOI22X1_95 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5343_), .D(AES_CORE_DATAPATH__abc_15863_new_n5347_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5351_));
AOI22X1 AOI22X1_96 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5381_), .D(AES_CORE_DATAPATH__abc_15863_new_n5387_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5391_));
AOI22X1 AOI22X1_97 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n3073_), .C(AES_CORE_DATAPATH__abc_15863_new_n5405_), .D(AES_CORE_DATAPATH__abc_15863_new_n5404_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5406_));
AOI22X1 AOI22X1_98 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3575_), .D(AES_CORE_DATAPATH__abc_15863_new_n3571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5422_));
AOI22X1 AOI22X1_99 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5421_), .D(AES_CORE_DATAPATH__abc_15863_new_n5425_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5429_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__0_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__9_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__1_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__10_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__2_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__11_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__3_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__12_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__4_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__13_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__5_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__14_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__6_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__15_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__7_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__16_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__0_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__17_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__1_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__18_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__1_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__19_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__3_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__20_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__4_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__21_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__5_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__22_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__6_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__23_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__7_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__24_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__0_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__25_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__1_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__26_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__2_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__27_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__3_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__28_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__4_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__2_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__29_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__5_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__30_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__6_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__31_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__7_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__3_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__4_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__5_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__6_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__6_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__7_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__7_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__8_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__0_));
DFFSR DFFSR_1 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_0_), .Q(AES_CORE_CONTROL_UNIT_state_0_), .R(1'h1), .S(rst_n));
DFFSR DFFSR_10 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_9_), .Q(AES_CORE_CONTROL_UNIT_state_9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_101 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_102 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_103 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_104 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_105 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_106 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_107 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_108 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_109 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_10_), .Q(AES_CORE_CONTROL_UNIT_key_gen), .R(rst_n), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1897), .Q(AES_CORE_CONTROL_UNIT_state_11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_120 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_12_), .Q(AES_CORE_CONTROL_UNIT_state_12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_130 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_134 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_14 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_13_), .Q(AES_CORE_CONTROL_UNIT_state_13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_140 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_149 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_14_), .Q(AES_CORE_CONTROL_UNIT_state_14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_150 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_153 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1928), .Q(AES_CORE_CONTROL_UNIT_state_15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_160 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__0_), .Q(AES_CORE_CONTROL_UNIT_rd_count_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_170 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_177 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__1_), .Q(AES_CORE_CONTROL_UNIT_rd_count_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_180 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__2_), .Q(AES_CORE_CONTROL_UNIT_rd_count_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_190 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_1_), .Q(AES_CORE_CONTROL_UNIT_state_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__3_), .Q(AES_CORE_CONTROL_UNIT_rd_count_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_200 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_210 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_220 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_230 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_240 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_248 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_25 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_250 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_251 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_252 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_253 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_254 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_260 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_270 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_273 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_276 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_277 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__0_), .Q(AES_CORE_DATAPATH_col_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_278 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__1_), .Q(AES_CORE_DATAPATH_col_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__2_), .Q(AES_CORE_DATAPATH_col_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_28 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_280 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__3_), .Q(AES_CORE_DATAPATH_col_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_281 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__4_), .Q(AES_CORE_DATAPATH_col_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_282 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__5_), .Q(AES_CORE_DATAPATH_col_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__6_), .Q(AES_CORE_DATAPATH_col_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__7_), .Q(AES_CORE_DATAPATH_col_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__8_), .Q(AES_CORE_DATAPATH_col_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__9_), .Q(AES_CORE_DATAPATH_col_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__10_), .Q(AES_CORE_DATAPATH_col_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__11_), .Q(AES_CORE_DATAPATH_col_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_289 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__12_), .Q(AES_CORE_DATAPATH_col_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_290 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__13_), .Q(AES_CORE_DATAPATH_col_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__14_), .Q(AES_CORE_DATAPATH_col_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__15_), .Q(AES_CORE_DATAPATH_col_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__16_), .Q(AES_CORE_DATAPATH_col_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__17_), .Q(AES_CORE_DATAPATH_col_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__18_), .Q(AES_CORE_DATAPATH_col_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__19_), .Q(AES_CORE_DATAPATH_col_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__20_), .Q(AES_CORE_DATAPATH_col_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__21_), .Q(AES_CORE_DATAPATH_col_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__22_), .Q(AES_CORE_DATAPATH_col_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_3 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_2_), .Q(AES_CORE_CONTROL_UNIT_state_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_300 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__23_), .Q(AES_CORE_DATAPATH_col_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_301 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__24_), .Q(AES_CORE_DATAPATH_col_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_302 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__25_), .Q(AES_CORE_DATAPATH_col_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_303 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__26_), .Q(AES_CORE_DATAPATH_col_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_304 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__27_), .Q(AES_CORE_DATAPATH_col_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_305 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__28_), .Q(AES_CORE_DATAPATH_col_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_306 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__29_), .Q(AES_CORE_DATAPATH_col_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_307 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__30_), .Q(AES_CORE_DATAPATH_col_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_308 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__31_), .Q(AES_CORE_DATAPATH_col_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_309 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__0_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_310 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__1_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_311 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__2_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_312 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__3_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_313 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__4_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_314 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__5_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_315 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__6_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_316 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__7_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_317 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__8_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_318 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__9_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_319 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__10_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_32 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_320 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__11_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_321 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__12_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_322 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__13_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_323 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__14_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_324 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__15_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_325 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__16_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_326 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__17_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_327 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__18_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_328 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__19_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_329 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__20_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_33 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_330 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__21_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_331 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__22_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_332 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__23_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_333 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__24_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_334 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__25_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_335 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__26_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_336 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__27_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_337 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__28_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_338 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__29_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_339 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__30_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_34 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_340 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__31_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_341 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__0_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_342 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__1_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_343 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__2_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_344 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__3_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_345 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__4_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_346 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__5_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_347 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__6_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_348 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__7_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_349 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__8_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_35 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_350 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__9_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_351 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__10_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_352 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__11_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_353 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__12_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_354 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__13_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_355 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__14_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_356 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__15_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_357 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__16_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_358 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__17_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_359 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__18_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_36 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_360 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__19_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_361 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__20_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_362 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__21_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_363 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__22_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_364 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__23_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_365 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__24_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_366 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__25_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_367 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__26_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_368 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__27_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_369 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__28_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_37 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_370 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__29_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_371 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__30_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_372 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__31_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_373 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__0_), .Q(AES_CORE_DATAPATH_col_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_374 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__1_), .Q(AES_CORE_DATAPATH_col_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_375 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__2_), .Q(AES_CORE_DATAPATH_col_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_376 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__3_), .Q(AES_CORE_DATAPATH_col_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_377 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__4_), .Q(AES_CORE_DATAPATH_col_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_378 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__5_), .Q(AES_CORE_DATAPATH_col_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_379 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__6_), .Q(AES_CORE_DATAPATH_col_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_38 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_380 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__7_), .Q(AES_CORE_DATAPATH_col_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_381 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__8_), .Q(AES_CORE_DATAPATH_col_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_382 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__9_), .Q(AES_CORE_DATAPATH_col_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_383 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__10_), .Q(AES_CORE_DATAPATH_col_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_384 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__11_), .Q(AES_CORE_DATAPATH_col_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_385 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__12_), .Q(AES_CORE_DATAPATH_col_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_386 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__13_), .Q(AES_CORE_DATAPATH_col_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_387 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__14_), .Q(AES_CORE_DATAPATH_col_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_388 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__15_), .Q(AES_CORE_DATAPATH_col_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_389 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__16_), .Q(AES_CORE_DATAPATH_col_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_39 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_390 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__17_), .Q(AES_CORE_DATAPATH_col_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_391 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__18_), .Q(AES_CORE_DATAPATH_col_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_392 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__19_), .Q(AES_CORE_DATAPATH_col_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_393 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__20_), .Q(AES_CORE_DATAPATH_col_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_394 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__21_), .Q(AES_CORE_DATAPATH_col_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_395 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__22_), .Q(AES_CORE_DATAPATH_col_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_396 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__23_), .Q(AES_CORE_DATAPATH_col_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_397 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__24_), .Q(AES_CORE_DATAPATH_col_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_398 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__25_), .Q(AES_CORE_DATAPATH_col_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_399 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__26_), .Q(AES_CORE_DATAPATH_col_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_4 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1817), .Q(AES_CORE_CONTROL_UNIT_state_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_400 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__27_), .Q(AES_CORE_DATAPATH_col_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_401 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__28_), .Q(AES_CORE_DATAPATH_col_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_402 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__29_), .Q(AES_CORE_DATAPATH_col_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_403 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__30_), .Q(AES_CORE_DATAPATH_col_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_404 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__31_), .Q(AES_CORE_DATAPATH_col_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_405 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__0_), .Q(AES_CORE_DATAPATH_iv_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_406 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__1_), .Q(AES_CORE_DATAPATH_iv_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_407 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__2_), .Q(AES_CORE_DATAPATH_iv_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_408 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__3_), .Q(AES_CORE_DATAPATH_iv_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_409 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__4_), .Q(AES_CORE_DATAPATH_iv_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_410 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__5_), .Q(AES_CORE_DATAPATH_iv_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_411 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__6_), .Q(AES_CORE_DATAPATH_iv_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_412 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__7_), .Q(AES_CORE_DATAPATH_iv_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_413 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__8_), .Q(AES_CORE_DATAPATH_iv_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_414 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__9_), .Q(AES_CORE_DATAPATH_iv_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_415 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__10_), .Q(AES_CORE_DATAPATH_iv_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_416 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__11_), .Q(AES_CORE_DATAPATH_iv_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_417 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__12_), .Q(AES_CORE_DATAPATH_iv_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_418 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__13_), .Q(AES_CORE_DATAPATH_iv_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_419 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__14_), .Q(AES_CORE_DATAPATH_iv_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_420 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__15_), .Q(AES_CORE_DATAPATH_iv_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_421 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__16_), .Q(AES_CORE_DATAPATH_iv_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_422 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__17_), .Q(AES_CORE_DATAPATH_iv_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_423 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__18_), .Q(AES_CORE_DATAPATH_iv_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_424 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__19_), .Q(AES_CORE_DATAPATH_iv_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_425 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__20_), .Q(AES_CORE_DATAPATH_iv_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_426 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__21_), .Q(AES_CORE_DATAPATH_iv_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_427 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__22_), .Q(AES_CORE_DATAPATH_iv_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_428 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__23_), .Q(AES_CORE_DATAPATH_iv_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_429 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__24_), .Q(AES_CORE_DATAPATH_iv_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_430 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__25_), .Q(AES_CORE_DATAPATH_iv_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_431 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__26_), .Q(AES_CORE_DATAPATH_iv_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_432 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__27_), .Q(AES_CORE_DATAPATH_iv_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_433 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__28_), .Q(AES_CORE_DATAPATH_iv_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_434 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__29_), .Q(AES_CORE_DATAPATH_iv_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_435 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__30_), .Q(AES_CORE_DATAPATH_iv_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_436 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__31_), .Q(AES_CORE_DATAPATH_iv_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_437 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_438 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_439 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_440 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_441 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_442 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_443 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_444 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_445 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_446 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_447 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_448 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_449 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_450 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_451 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_452 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_453 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_454 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_455 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_456 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_457 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_458 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_459 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_460 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_461 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_462 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_463 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_464 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_465 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_466 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_467 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_468 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_469 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_470 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_471 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_472 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_473 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_474 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_475 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_476 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_477 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_478 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_479 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_480 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_481 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_482 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_483 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_484 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_485 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_486 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_487 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_488 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_489 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_490 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_491 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_492 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_493 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_494 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_495 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_496 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_497 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_498 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_499 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_5 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_4_), .Q(AES_CORE_CONTROL_UNIT_state_4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_500 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_501 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__0_), .Q(AES_CORE_DATAPATH_iv_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_502 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__1_), .Q(AES_CORE_DATAPATH_iv_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_503 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__2_), .Q(AES_CORE_DATAPATH_iv_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_504 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__3_), .Q(AES_CORE_DATAPATH_iv_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_505 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__4_), .Q(AES_CORE_DATAPATH_iv_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_506 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__5_), .Q(AES_CORE_DATAPATH_iv_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_507 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__6_), .Q(AES_CORE_DATAPATH_iv_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_508 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__7_), .Q(AES_CORE_DATAPATH_iv_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_509 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__8_), .Q(AES_CORE_DATAPATH_iv_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_51 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_510 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__9_), .Q(AES_CORE_DATAPATH_iv_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_511 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__10_), .Q(AES_CORE_DATAPATH_iv_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_512 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__11_), .Q(AES_CORE_DATAPATH_iv_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_513 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__12_), .Q(AES_CORE_DATAPATH_iv_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_514 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__13_), .Q(AES_CORE_DATAPATH_iv_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_515 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__14_), .Q(AES_CORE_DATAPATH_iv_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_516 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__15_), .Q(AES_CORE_DATAPATH_iv_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_517 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__16_), .Q(AES_CORE_DATAPATH_iv_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_518 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__17_), .Q(AES_CORE_DATAPATH_iv_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_519 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__18_), .Q(AES_CORE_DATAPATH_iv_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_52 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_520 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__19_), .Q(AES_CORE_DATAPATH_iv_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_521 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__20_), .Q(AES_CORE_DATAPATH_iv_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_522 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__21_), .Q(AES_CORE_DATAPATH_iv_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_523 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__22_), .Q(AES_CORE_DATAPATH_iv_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_524 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__23_), .Q(AES_CORE_DATAPATH_iv_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_525 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__24_), .Q(AES_CORE_DATAPATH_iv_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_526 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__25_), .Q(AES_CORE_DATAPATH_iv_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_527 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__26_), .Q(AES_CORE_DATAPATH_iv_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_528 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__27_), .Q(AES_CORE_DATAPATH_iv_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_529 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__28_), .Q(AES_CORE_DATAPATH_iv_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_53 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_530 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__29_), .Q(AES_CORE_DATAPATH_iv_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_531 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__30_), .Q(AES_CORE_DATAPATH_iv_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_532 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__31_), .Q(AES_CORE_DATAPATH_iv_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_533 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_534 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_535 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_536 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_537 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_538 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_539 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_54 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_540 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_541 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_542 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_543 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_544 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_545 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_546 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_547 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_548 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_549 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_55 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_550 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_551 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_552 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_553 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_554 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_555 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_556 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_557 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_558 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_559 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_56 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_560 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_561 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_562 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_563 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_564 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_565 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_566 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_567 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_568 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_569 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_57 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_570 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_571 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_572 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_573 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_574 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_575 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_576 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_577 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_578 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_579 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_58 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_580 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_581 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_582 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_583 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_584 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_585 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_586 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_587 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_588 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_589 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_59 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_590 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_591 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_592 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_593 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_594 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_595 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_596 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_597 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__0_), .Q(AES_CORE_DATAPATH_iv_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_598 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__1_), .Q(AES_CORE_DATAPATH_iv_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_599 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__2_), .Q(AES_CORE_DATAPATH_iv_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_6 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_5_), .Q(end_aes), .R(rst_n), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_600 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__3_), .Q(AES_CORE_DATAPATH_iv_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_601 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__4_), .Q(AES_CORE_DATAPATH_iv_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_602 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__5_), .Q(AES_CORE_DATAPATH_iv_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_603 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__6_), .Q(AES_CORE_DATAPATH_iv_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_604 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__7_), .Q(AES_CORE_DATAPATH_iv_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_605 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__8_), .Q(AES_CORE_DATAPATH_iv_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_606 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__9_), .Q(AES_CORE_DATAPATH_iv_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_607 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__10_), .Q(AES_CORE_DATAPATH_iv_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_608 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__11_), .Q(AES_CORE_DATAPATH_iv_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_609 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__12_), .Q(AES_CORE_DATAPATH_iv_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_61 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_610 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__13_), .Q(AES_CORE_DATAPATH_iv_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_611 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__14_), .Q(AES_CORE_DATAPATH_iv_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_612 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__15_), .Q(AES_CORE_DATAPATH_iv_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_613 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__16_), .Q(AES_CORE_DATAPATH_iv_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_614 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__17_), .Q(AES_CORE_DATAPATH_iv_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_615 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__18_), .Q(AES_CORE_DATAPATH_iv_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_616 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__19_), .Q(AES_CORE_DATAPATH_iv_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_617 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__20_), .Q(AES_CORE_DATAPATH_iv_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_618 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__21_), .Q(AES_CORE_DATAPATH_iv_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_619 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__22_), .Q(AES_CORE_DATAPATH_iv_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_62 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_620 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__23_), .Q(AES_CORE_DATAPATH_iv_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_621 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__24_), .Q(AES_CORE_DATAPATH_iv_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_622 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__25_), .Q(AES_CORE_DATAPATH_iv_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_623 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__26_), .Q(AES_CORE_DATAPATH_iv_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_624 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__27_), .Q(AES_CORE_DATAPATH_iv_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_625 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__28_), .Q(AES_CORE_DATAPATH_iv_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_626 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__29_), .Q(AES_CORE_DATAPATH_iv_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_627 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__30_), .Q(AES_CORE_DATAPATH_iv_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_628 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__31_), .Q(AES_CORE_DATAPATH_iv_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_629 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_63 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_630 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_631 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_632 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_633 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_634 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_635 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_636 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_637 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_638 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_639 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_64 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_640 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_641 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_642 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_643 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_644 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_645 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_646 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_647 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_648 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_649 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_65 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_650 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_651 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_652 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_653 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_654 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_655 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_656 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_657 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_658 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_659 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_66 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_660 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_661 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_662 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_663 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_664 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_665 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_666 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_667 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_668 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_669 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_67 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_670 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_671 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_672 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_673 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_674 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_675 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_676 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_677 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_678 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_679 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_68 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_680 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_681 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_682 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_683 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_684 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_685 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_686 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_687 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_688 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_689 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_69 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_690 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_691 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_692 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_693 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__0_), .Q(AES_CORE_DATAPATH_iv_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_694 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__1_), .Q(AES_CORE_DATAPATH_iv_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_695 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__2_), .Q(AES_CORE_DATAPATH_iv_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_696 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__3_), .Q(AES_CORE_DATAPATH_iv_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_697 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__4_), .Q(AES_CORE_DATAPATH_iv_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_698 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__5_), .Q(AES_CORE_DATAPATH_iv_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_699 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__6_), .Q(AES_CORE_DATAPATH_iv_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_7 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_6_), .Q(AES_CORE_CONTROL_UNIT_state_6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_700 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__7_), .Q(AES_CORE_DATAPATH_iv_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_701 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__8_), .Q(AES_CORE_DATAPATH_iv_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_702 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__9_), .Q(AES_CORE_DATAPATH_iv_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_703 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__10_), .Q(AES_CORE_DATAPATH_iv_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_704 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__11_), .Q(AES_CORE_DATAPATH_iv_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_705 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__12_), .Q(AES_CORE_DATAPATH_iv_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_706 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__13_), .Q(AES_CORE_DATAPATH_iv_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_707 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__14_), .Q(AES_CORE_DATAPATH_iv_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_708 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__15_), .Q(AES_CORE_DATAPATH_iv_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_709 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__16_), .Q(AES_CORE_DATAPATH_iv_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_71 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_710 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__17_), .Q(AES_CORE_DATAPATH_iv_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_711 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__18_), .Q(AES_CORE_DATAPATH_iv_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_712 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__19_), .Q(AES_CORE_DATAPATH_iv_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_713 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__20_), .Q(AES_CORE_DATAPATH_iv_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_714 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__21_), .Q(AES_CORE_DATAPATH_iv_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_715 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__22_), .Q(AES_CORE_DATAPATH_iv_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_716 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__23_), .Q(AES_CORE_DATAPATH_iv_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_717 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__24_), .Q(AES_CORE_DATAPATH_iv_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_718 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__25_), .Q(AES_CORE_DATAPATH_iv_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_719 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__26_), .Q(AES_CORE_DATAPATH_iv_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_72 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_720 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__27_), .Q(AES_CORE_DATAPATH_iv_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_721 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__28_), .Q(AES_CORE_DATAPATH_iv_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_722 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__29_), .Q(AES_CORE_DATAPATH_iv_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_723 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__30_), .Q(AES_CORE_DATAPATH_iv_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_724 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__31_), .Q(AES_CORE_DATAPATH_iv_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_725 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_726 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_727 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_728 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_729 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_73 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_730 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_731 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_732 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_733 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_734 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_735 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_736 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_737 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_738 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_739 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_74 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_740 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_741 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_742 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_743 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_744 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_745 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_746 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_747 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_748 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_749 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_75 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_750 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_751 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_752 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_753 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_754 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_755 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_756 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_757 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_758 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_759 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_76 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_760 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_761 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_762 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_763 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_764 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_765 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_766 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_767 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_768 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_769 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_77 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_770 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_771 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_772 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_773 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_774 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_775 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_776 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_777 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_778 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_779 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_780 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_781 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_782 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_783 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_784 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_785 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_786 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_787 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_788 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_789 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__0_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_790 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__1_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_791 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__2_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_792 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__3_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_793 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__0_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_794 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__1_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_795 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__2_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_796 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__3_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_797 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__0_), .Q(AES_CORE_DATAPATH_key_en_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_798 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__1_), .Q(AES_CORE_DATAPATH_key_en_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_799 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__2_), .Q(AES_CORE_DATAPATH_key_en_pp1_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1856), .Q(AES_CORE_CONTROL_UNIT_state_7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_800 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__3_), .Q(AES_CORE_DATAPATH_key_en_pp1_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_801 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_802 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_803 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_804 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_805 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_col_sel_0_), .Q(AES_CORE_DATAPATH_col_sel_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_806 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_col_sel_1_), .Q(AES_CORE_DATAPATH_col_sel_pp1_1_), .R(1'h1), .S(rst_n));
DFFSR DFFSR_807 ( .CLK(clk), .D(AES_CORE_DATAPATH_col_sel_pp1_0_), .Q(AES_CORE_DATAPATH_col_sel_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_808 ( .CLK(clk), .D(AES_CORE_DATAPATH_col_sel_pp1_1_), .Q(AES_CORE_DATAPATH_col_sel_pp2_1_), .R(1'h1), .S(rst_n));
DFFSR DFFSR_809 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_key_out_sel_0_), .Q(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_810 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_key_out_sel_1_), .Q(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_811 ( .CLK(clk), .D(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Q(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_812 ( .CLK(clk), .D(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Q(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_813 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rk_sel_0_), .Q(AES_CORE_DATAPATH_rk_sel_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_814 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rk_sel_1_), .Q(AES_CORE_DATAPATH_rk_sel_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_815 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_sel_pp1_0_), .Q(AES_CORE_DATAPATH_rk_sel_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_816 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_sel_pp1_1_), .Q(AES_CORE_DATAPATH_rk_sel_pp2_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_817 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_key_sel), .Q(AES_CORE_DATAPATH_key_sel_pp1), .R(rst_n), .S(1'h1));
DFFSR DFFSR_818 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_out_sel), .Q(AES_CORE_DATAPATH_rk_out_sel_pp1), .R(1'h1), .S(rst_n));
DFFSR DFFSR_819 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_out_sel_pp1), .Q(AES_CORE_DATAPATH_rk_out_sel_pp2), .R(1'h1), .S(rst_n));
DFFSR DFFSR_82 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_820 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_last_round), .Q(AES_CORE_DATAPATH_last_round_pp1), .R(1'h1), .S(rst_n));
DFFSR DFFSR_821 ( .CLK(clk), .D(AES_CORE_DATAPATH_last_round_pp1), .Q(AES_CORE_DATAPATH_last_round_pp2), .R(rst_n), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_8_), .Q(AES_CORE_CONTROL_UNIT_state_8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_97 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_98 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_99 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_1__14_), .R(rst_n), .S(1'h1));
INVX1 INVX1_1 ( .A(write_en), .Y(_abc_15574_new_n11_));
INVX1 INVX1_10 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_));
INVX1 INVX1_100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2749_));
INVX1 INVX1_1000 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n363_));
INVX1 INVX1_1001 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n364_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n365_));
INVX1 INVX1_1002 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n366_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n368_));
INVX1 INVX1_1003 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n384_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_));
INVX1 INVX1_1004 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n411_));
INVX1 INVX1_1005 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n421_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_));
INVX1 INVX1_1006 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n349_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n423_));
INVX1 INVX1_1007 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n469_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_));
INVX1 INVX1_1008 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n476_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_));
INVX1 INVX1_1009 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n492_));
INVX1 INVX1_101 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2751_), .Y(\key_out[1] ));
INVX1 INVX1_1010 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n502_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_));
INVX1 INVX1_1011 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n516_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_));
INVX1 INVX1_1012 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n523_));
INVX1 INVX1_1013 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_));
INVX1 INVX1_1014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_));
INVX1 INVX1_1015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n62_));
INVX1 INVX1_1016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_));
INVX1 INVX1_1017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n69_));
INVX1 INVX1_1018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n80_));
INVX1 INVX1_1019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n82_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_));
INVX1 INVX1_102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2754_));
INVX1 INVX1_1020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n86_));
INVX1 INVX1_1021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n90_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n91_));
INVX1 INVX1_1022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n92_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n93_));
INVX1 INVX1_1023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_));
INVX1 INVX1_1024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n99_));
INVX1 INVX1_1025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n106_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n107_));
INVX1 INVX1_1026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n118_));
INVX1 INVX1_1027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n121_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n128_));
INVX1 INVX1_1028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_));
INVX1 INVX1_1029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_));
INVX1 INVX1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2755_));
INVX1 INVX1_1030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n138_));
INVX1 INVX1_1031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n143_));
INVX1 INVX1_1032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n152_));
INVX1 INVX1_1033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_));
INVX1 INVX1_1034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n158_));
INVX1 INVX1_1035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n159_));
INVX1 INVX1_1036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n166_));
INVX1 INVX1_1037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_));
INVX1 INVX1_1038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n170_));
INVX1 INVX1_1039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n182_));
INVX1 INVX1_104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2762_));
INVX1 INVX1_1040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n201_));
INVX1 INVX1_1041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n206_));
INVX1 INVX1_1042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n207_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n208_));
INVX1 INVX1_1043 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n213_));
INVX1 INVX1_1044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n216_));
INVX1 INVX1_1045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n220_));
INVX1 INVX1_1046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n227_));
INVX1 INVX1_1047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n235_));
INVX1 INVX1_1048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n238_));
INVX1 INVX1_1049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n162_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n255_));
INVX1 INVX1_105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2768_));
INVX1 INVX1_1050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n260_));
INVX1 INVX1_1051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n279_));
INVX1 INVX1_1052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n319_));
INVX1 INVX1_1053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n373_));
INVX1 INVX1_1054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n385_));
INVX1 INVX1_1055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n403_));
INVX1 INVX1_1056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n407_));
INVX1 INVX1_1057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n428_));
INVX1 INVX1_1058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n440_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n442_));
INVX1 INVX1_1059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n462_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n463_));
INVX1 INVX1_106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2778_));
INVX1 INVX1_1060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n478_));
INVX1 INVX1_1061 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n302_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n491_));
INVX1 INVX1_1062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n492_));
INVX1 INVX1_1063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n494_));
INVX1 INVX1_1064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n495_));
INVX1 INVX1_1065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_));
INVX1 INVX1_1066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_));
INVX1 INVX1_1067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n62_));
INVX1 INVX1_1068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_));
INVX1 INVX1_1069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n69_));
INVX1 INVX1_107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2792_));
INVX1 INVX1_1070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n80_));
INVX1 INVX1_1071 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n82_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_));
INVX1 INVX1_1072 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n86_));
INVX1 INVX1_1073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n90_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n91_));
INVX1 INVX1_1074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n92_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n93_));
INVX1 INVX1_1075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_));
INVX1 INVX1_1076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n99_));
INVX1 INVX1_1077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n106_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n107_));
INVX1 INVX1_1078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n118_));
INVX1 INVX1_1079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n121_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n128_));
INVX1 INVX1_108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2798_));
INVX1 INVX1_1080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_));
INVX1 INVX1_1081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_));
INVX1 INVX1_1082 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n138_));
INVX1 INVX1_1083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n143_));
INVX1 INVX1_1084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n152_));
INVX1 INVX1_1085 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_));
INVX1 INVX1_1086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n158_));
INVX1 INVX1_1087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n159_));
INVX1 INVX1_1088 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n166_));
INVX1 INVX1_1089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_));
INVX1 INVX1_109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2813_));
INVX1 INVX1_1090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n170_));
INVX1 INVX1_1091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n182_));
INVX1 INVX1_1092 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n201_));
INVX1 INVX1_1093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n206_));
INVX1 INVX1_1094 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n207_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n208_));
INVX1 INVX1_1095 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n213_));
INVX1 INVX1_1096 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n216_));
INVX1 INVX1_1097 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n220_));
INVX1 INVX1_1098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n227_));
INVX1 INVX1_1099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n235_));
INVX1 INVX1_11 ( .A(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n108_));
INVX1 INVX1_110 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2815_), .Y(\key_out[7] ));
INVX1 INVX1_1100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n238_));
INVX1 INVX1_1101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n162_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n255_));
INVX1 INVX1_1102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n260_));
INVX1 INVX1_1103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n279_));
INVX1 INVX1_1104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n319_));
INVX1 INVX1_1105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n373_));
INVX1 INVX1_1106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n385_));
INVX1 INVX1_1107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n403_));
INVX1 INVX1_1108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n407_));
INVX1 INVX1_1109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n428_));
INVX1 INVX1_111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2818_));
INVX1 INVX1_1110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n440_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n442_));
INVX1 INVX1_1111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n462_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n463_));
INVX1 INVX1_1112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n478_));
INVX1 INVX1_1113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n302_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n491_));
INVX1 INVX1_1114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n492_));
INVX1 INVX1_1115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n494_));
INVX1 INVX1_1116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n495_));
INVX1 INVX1_1117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_));
INVX1 INVX1_1118 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_));
INVX1 INVX1_1119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n62_));
INVX1 INVX1_112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2826_));
INVX1 INVX1_1120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_));
INVX1 INVX1_1121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n69_));
INVX1 INVX1_1122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n80_));
INVX1 INVX1_1123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n82_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_));
INVX1 INVX1_1124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n86_));
INVX1 INVX1_1125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n90_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n91_));
INVX1 INVX1_1126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n92_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n93_));
INVX1 INVX1_1127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_));
INVX1 INVX1_1128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n99_));
INVX1 INVX1_1129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n106_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n107_));
INVX1 INVX1_113 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2828_), .Y(\key_out[8] ));
INVX1 INVX1_1130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n118_));
INVX1 INVX1_1131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n121_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n128_));
INVX1 INVX1_1132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_));
INVX1 INVX1_1133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_));
INVX1 INVX1_1134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n138_));
INVX1 INVX1_1135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n143_));
INVX1 INVX1_1136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n152_));
INVX1 INVX1_1137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_));
INVX1 INVX1_1138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n158_));
INVX1 INVX1_1139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n159_));
INVX1 INVX1_114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2831_));
INVX1 INVX1_1140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n166_));
INVX1 INVX1_1141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_));
INVX1 INVX1_1142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n170_));
INVX1 INVX1_1143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n182_));
INVX1 INVX1_1144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n201_));
INVX1 INVX1_1145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n206_));
INVX1 INVX1_1146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n207_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n208_));
INVX1 INVX1_1147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n213_));
INVX1 INVX1_1148 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n216_));
INVX1 INVX1_1149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n220_));
INVX1 INVX1_115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2838_));
INVX1 INVX1_1150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n227_));
INVX1 INVX1_1151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n235_));
INVX1 INVX1_1152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n238_));
INVX1 INVX1_1153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n162_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n255_));
INVX1 INVX1_1154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n260_));
INVX1 INVX1_1155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n279_));
INVX1 INVX1_1156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n319_));
INVX1 INVX1_1157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n373_));
INVX1 INVX1_1158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n385_));
INVX1 INVX1_1159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n403_));
INVX1 INVX1_116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2849_));
INVX1 INVX1_1160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n407_));
INVX1 INVX1_1161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n428_));
INVX1 INVX1_1162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n440_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n442_));
INVX1 INVX1_1163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n462_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n463_));
INVX1 INVX1_1164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n478_));
INVX1 INVX1_1165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n302_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n491_));
INVX1 INVX1_1166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n492_));
INVX1 INVX1_1167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n494_));
INVX1 INVX1_1168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n495_));
INVX1 INVX1_1169 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_));
INVX1 INVX1_117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2858_));
INVX1 INVX1_1170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_));
INVX1 INVX1_1171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n62_));
INVX1 INVX1_1172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_));
INVX1 INVX1_1173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n69_));
INVX1 INVX1_1174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n80_));
INVX1 INVX1_1175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n82_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_));
INVX1 INVX1_1176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n86_));
INVX1 INVX1_1177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n90_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n91_));
INVX1 INVX1_1178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n92_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n93_));
INVX1 INVX1_1179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_));
INVX1 INVX1_118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2868_));
INVX1 INVX1_1180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n99_));
INVX1 INVX1_1181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n106_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n107_));
INVX1 INVX1_1182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n118_));
INVX1 INVX1_1183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n121_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n128_));
INVX1 INVX1_1184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_));
INVX1 INVX1_1185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_));
INVX1 INVX1_1186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n137_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n138_));
INVX1 INVX1_1187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n143_));
INVX1 INVX1_1188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n152_));
INVX1 INVX1_1189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_));
INVX1 INVX1_119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2874_));
INVX1 INVX1_1190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n158_));
INVX1 INVX1_1191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n159_));
INVX1 INVX1_1192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n166_));
INVX1 INVX1_1193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_));
INVX1 INVX1_1194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n170_));
INVX1 INVX1_1195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n182_));
INVX1 INVX1_1196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n201_));
INVX1 INVX1_1197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n206_));
INVX1 INVX1_1198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n207_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n208_));
INVX1 INVX1_1199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n213_));
INVX1 INVX1_12 ( .A(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_));
INVX1 INVX1_120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2888_));
INVX1 INVX1_1200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n216_));
INVX1 INVX1_1201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n220_));
INVX1 INVX1_1202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n227_));
INVX1 INVX1_1203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n234_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n235_));
INVX1 INVX1_1204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n238_));
INVX1 INVX1_1205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n162_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n255_));
INVX1 INVX1_1206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n260_));
INVX1 INVX1_1207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n279_));
INVX1 INVX1_1208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n319_));
INVX1 INVX1_1209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n373_));
INVX1 INVX1_121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2894_));
INVX1 INVX1_1210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n385_));
INVX1 INVX1_1211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n403_));
INVX1 INVX1_1212 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n407_));
INVX1 INVX1_1213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n428_));
INVX1 INVX1_1214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n440_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n442_));
INVX1 INVX1_1215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n462_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n463_));
INVX1 INVX1_1216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n478_));
INVX1 INVX1_1217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n302_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n491_));
INVX1 INVX1_1218 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n492_));
INVX1 INVX1_1219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n494_));
INVX1 INVX1_122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2905_));
INVX1 INVX1_1220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n495_));
INVX1 INVX1_1221 ( .A(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_));
INVX1 INVX1_1222 ( .A(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_));
INVX1 INVX1_1223 ( .A(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_));
INVX1 INVX1_1224 ( .A(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_));
INVX1 INVX1_123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2914_));
INVX1 INVX1_124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2924_));
INVX1 INVX1_125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2934_));
INVX1 INVX1_126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2945_));
INVX1 INVX1_127 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2951_), .Y(\key_out[20] ));
INVX1 INVX1_128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2954_));
INVX1 INVX1_129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2957_));
INVX1 INVX1_13 ( .A(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n119_));
INVX1 INVX1_130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2967_));
INVX1 INVX1_131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2978_));
INVX1 INVX1_132 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2984_), .Y(\key_out[23] ));
INVX1 INVX1_133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2987_));
INVX1 INVX1_134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2995_));
INVX1 INVX1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2997_), .Y(\key_out[24] ));
INVX1 INVX1_136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3000_));
INVX1 INVX1_137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3007_));
INVX1 INVX1_138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3017_));
INVX1 INVX1_139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3027_));
INVX1 INVX1_14 ( .A(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_));
INVX1 INVX1_140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3038_));
INVX1 INVX1_141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3048_));
INVX1 INVX1_142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3058_));
INVX1 INVX1_143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3063_));
INVX1 INVX1_144 ( .A(AES_CORE_DATAPATH_rk_out_sel_pp2), .Y(AES_CORE_DATAPATH__abc_15863_new_n3073_));
INVX1 INVX1_145 ( .A(AES_CORE_DATAPATH_rk_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3074_));
INVX1 INVX1_146 ( .A(AES_CORE_DATAPATH_rk_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3077_));
INVX1 INVX1_147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3081_));
INVX1 INVX1_148 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3083_));
INVX1 INVX1_149 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3079_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3098_));
INVX1 INVX1_15 ( .A(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n122_));
INVX1 INVX1_150 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3107_));
INVX1 INVX1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3111_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3112_));
INVX1 INVX1_152 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3115_));
INVX1 INVX1_153 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3116_));
INVX1 INVX1_154 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3131_));
INVX1 INVX1_155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3134_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3135_));
INVX1 INVX1_156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3138_));
INVX1 INVX1_157 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3153_));
INVX1 INVX1_158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3156_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3157_));
INVX1 INVX1_159 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3160_));
INVX1 INVX1_16 ( .A(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_));
INVX1 INVX1_160 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3161_));
INVX1 INVX1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3168_));
INVX1 INVX1_162 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3176_));
INVX1 INVX1_163 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3178_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3179_));
INVX1 INVX1_164 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3183_));
INVX1 INVX1_165 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3198_));
INVX1 INVX1_166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3201_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3202_));
INVX1 INVX1_167 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3205_));
INVX1 INVX1_168 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3220_));
INVX1 INVX1_169 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3223_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3224_));
INVX1 INVX1_17 ( .A(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_));
INVX1 INVX1_170 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3227_));
INVX1 INVX1_171 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3242_));
INVX1 INVX1_172 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3245_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3246_));
INVX1 INVX1_173 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3249_));
INVX1 INVX1_174 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3250_));
INVX1 INVX1_175 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3264_));
INVX1 INVX1_176 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3267_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3268_));
INVX1 INVX1_177 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3271_));
INVX1 INVX1_178 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3286_));
INVX1 INVX1_179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3289_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3290_));
INVX1 INVX1_18 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_), .Y(AES_CORE_CONTROL_UNIT_mode_cbc));
INVX1 INVX1_180 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3293_));
INVX1 INVX1_181 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3294_));
INVX1 INVX1_182 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3308_));
INVX1 INVX1_183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3310_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3311_));
INVX1 INVX1_184 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3315_));
INVX1 INVX1_185 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3330_));
INVX1 INVX1_186 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3333_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3334_));
INVX1 INVX1_187 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3337_));
INVX1 INVX1_188 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3338_));
INVX1 INVX1_189 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3352_));
INVX1 INVX1_19 ( .A(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_));
INVX1 INVX1_190 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3354_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3355_));
INVX1 INVX1_191 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3359_));
INVX1 INVX1_192 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3374_));
INVX1 INVX1_193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3377_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3378_));
INVX1 INVX1_194 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3381_));
INVX1 INVX1_195 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3382_));
INVX1 INVX1_196 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3396_));
INVX1 INVX1_197 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3398_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3399_));
INVX1 INVX1_198 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3403_));
INVX1 INVX1_199 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3418_));
INVX1 INVX1_2 ( .A(\addr[1] ), .Y(_abc_15574_new_n15_));
INVX1 INVX1_20 ( .A(AES_CORE_CONTROL_UNIT_rd_count_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_));
INVX1 INVX1_200 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3421_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3422_));
INVX1 INVX1_201 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3425_));
INVX1 INVX1_202 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3426_));
INVX1 INVX1_203 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3440_));
INVX1 INVX1_204 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3443_));
INVX1 INVX1_205 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3447_));
INVX1 INVX1_206 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3462_));
INVX1 INVX1_207 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3465_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3466_));
INVX1 INVX1_208 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3469_));
INVX1 INVX1_209 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3470_));
INVX1 INVX1_21 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_));
INVX1 INVX1_210 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3484_));
INVX1 INVX1_211 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3486_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3487_));
INVX1 INVX1_212 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3491_));
INVX1 INVX1_213 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3492_));
INVX1 INVX1_214 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3506_));
INVX1 INVX1_215 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3508_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3509_));
INVX1 INVX1_216 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3513_));
INVX1 INVX1_217 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3514_));
INVX1 INVX1_218 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3528_));
INVX1 INVX1_219 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3530_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3531_));
INVX1 INVX1_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n161_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n162_));
INVX1 INVX1_220 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3535_));
INVX1 INVX1_221 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3550_));
INVX1 INVX1_222 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3553_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3554_));
INVX1 INVX1_223 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3557_));
INVX1 INVX1_224 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3558_));
INVX1 INVX1_225 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3572_));
INVX1 INVX1_226 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3574_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3575_));
INVX1 INVX1_227 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3579_));
INVX1 INVX1_228 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3594_));
INVX1 INVX1_229 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3597_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3598_));
INVX1 INVX1_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n179_));
INVX1 INVX1_230 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3601_));
INVX1 INVX1_231 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3602_));
INVX1 INVX1_232 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3616_));
INVX1 INVX1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3619_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3620_));
INVX1 INVX1_234 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3623_));
INVX1 INVX1_235 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3638_));
INVX1 INVX1_236 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3641_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3642_));
INVX1 INVX1_237 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3645_));
INVX1 INVX1_238 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3646_));
INVX1 INVX1_239 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3660_));
INVX1 INVX1_24 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n146_), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_2_));
INVX1 INVX1_240 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3662_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3663_));
INVX1 INVX1_241 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3667_));
INVX1 INVX1_242 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3668_));
INVX1 INVX1_243 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3682_));
INVX1 INVX1_244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3684_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3685_));
INVX1 INVX1_245 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3689_));
INVX1 INVX1_246 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3704_));
INVX1 INVX1_247 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3707_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3708_));
INVX1 INVX1_248 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3711_));
INVX1 INVX1_249 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3712_));
INVX1 INVX1_25 ( .A(end_aes), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n210_));
INVX1 INVX1_250 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3726_));
INVX1 INVX1_251 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3729_));
INVX1 INVX1_252 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3733_));
INVX1 INVX1_253 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3748_));
INVX1 INVX1_254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3751_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3752_));
INVX1 INVX1_255 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3755_));
INVX1 INVX1_256 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3770_));
INVX1 INVX1_257 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3773_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3774_));
INVX1 INVX1_258 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3777_));
INVX1 INVX1_259 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3778_));
INVX1 INVX1_26 ( .A(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2457_));
INVX1 INVX1_260 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3792_));
INVX1 INVX1_261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3794_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3795_));
INVX1 INVX1_262 ( .A(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4023_));
INVX1 INVX1_263 ( .A(AES_CORE_CONTROL_UNIT_key_en_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4030_));
INVX1 INVX1_264 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4035_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4036_));
INVX1 INVX1_265 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n4198_));
INVX1 INVX1_266 ( .A(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4231_));
INVX1 INVX1_267 ( .A(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4236_));
INVX1 INVX1_268 ( .A(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4241_));
INVX1 INVX1_269 ( .A(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4246_));
INVX1 INVX1_27 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_DATAPATH__abc_15863_new_n2458_));
INVX1 INVX1_270 ( .A(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4251_));
INVX1 INVX1_271 ( .A(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4256_));
INVX1 INVX1_272 ( .A(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4279_));
INVX1 INVX1_273 ( .A(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4284_));
INVX1 INVX1_274 ( .A(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4289_));
INVX1 INVX1_275 ( .A(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4294_));
INVX1 INVX1_276 ( .A(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4299_));
INVX1 INVX1_277 ( .A(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4304_));
INVX1 INVX1_278 ( .A(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4309_));
INVX1 INVX1_279 ( .A(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4314_));
INVX1 INVX1_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2462_));
INVX1 INVX1_280 ( .A(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4319_));
INVX1 INVX1_281 ( .A(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4324_));
INVX1 INVX1_282 ( .A(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4329_));
INVX1 INVX1_283 ( .A(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4334_));
INVX1 INVX1_284 ( .A(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4339_));
INVX1 INVX1_285 ( .A(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4344_));
INVX1 INVX1_286 ( .A(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4349_));
INVX1 INVX1_287 ( .A(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4354_));
INVX1 INVX1_288 ( .A(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4359_));
INVX1 INVX1_289 ( .A(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4364_));
INVX1 INVX1_29 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2468_));
INVX1 INVX1_290 ( .A(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4369_));
INVX1 INVX1_291 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2478_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4571_));
INVX1 INVX1_292 ( .A(AES_CORE_DATAPATH_col_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4573_));
INVX1 INVX1_293 ( .A(AES_CORE_DATAPATH_col_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4576_));
INVX1 INVX1_294 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4579_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4580_));
INVX1 INVX1_295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4582_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4583_));
INVX1 INVX1_296 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4578_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4584_));
INVX1 INVX1_297 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4587_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4588_));
INVX1 INVX1_298 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3110_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4591_));
INVX1 INVX1_299 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4593_));
INVX1 INVX1_3 ( .A(_abc_15574_new_n17_), .Y(AES_CORE_DATAPATH_col_en_host_3_));
INVX1 INVX1_30 ( .A(AES_CORE_DATAPATH_iv_1__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2469_));
INVX1 INVX1_300 ( .A(first_block), .Y(AES_CORE_DATAPATH__abc_15863_new_n4596_));
INVX1 INVX1_301 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4598_));
INVX1 INVX1_302 ( .A(AES_CORE_DATAPATH_bkp_2__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4599_));
INVX1 INVX1_303 ( .A(AES_CORE_DATAPATH_bkp_3__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4605_));
INVX1 INVX1_304 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4612_));
INVX1 INVX1_305 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_15863_new_n4621_));
INVX1 INVX1_306 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4623_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4624_));
INVX1 INVX1_307 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4630_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4631_));
INVX1 INVX1_308 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4635_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4636_));
INVX1 INVX1_309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4638_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4639_));
INVX1 INVX1_31 ( .A(\iv_sel_rd[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2470_));
INVX1 INVX1_310 ( .A(AES_CORE_DATAPATH_bkp_2__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4640_));
INVX1 INVX1_311 ( .A(AES_CORE_DATAPATH_bkp_3__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4646_));
INVX1 INVX1_312 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3133_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4655_));
INVX1 INVX1_313 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4669_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4670_));
INVX1 INVX1_314 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4674_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4675_));
INVX1 INVX1_315 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3155_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4678_));
INVX1 INVX1_316 ( .A(AES_CORE_DATAPATH_bkp_2__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4681_));
INVX1 INVX1_317 ( .A(AES_CORE_DATAPATH_bkp_3__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4687_));
INVX1 INVX1_318 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4694_));
INVX1 INVX1_319 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4708_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4709_));
INVX1 INVX1_32 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2473_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2474_));
INVX1 INVX1_320 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4714_));
INVX1 INVX1_321 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4719_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4720_));
INVX1 INVX1_322 ( .A(AES_CORE_DATAPATH_bkp_2__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4721_));
INVX1 INVX1_323 ( .A(AES_CORE_DATAPATH_bkp_3__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4727_));
INVX1 INVX1_324 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4745_));
INVX1 INVX1_325 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4746_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4747_));
INVX1 INVX1_326 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4748_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4749_));
INVX1 INVX1_327 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4753_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4754_));
INVX1 INVX1_328 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3200_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4757_));
INVX1 INVX1_329 ( .A(AES_CORE_DATAPATH_bkp_2__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4763_));
INVX1 INVX1_33 ( .A(AES_CORE_DATAPATH_iv_2__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2481_));
INVX1 INVX1_330 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4770_));
INVX1 INVX1_331 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4784_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4785_));
INVX1 INVX1_332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4789_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4790_));
INVX1 INVX1_333 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3222_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4793_));
INVX1 INVX1_334 ( .A(AES_CORE_DATAPATH_bkp_2__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4796_));
INVX1 INVX1_335 ( .A(AES_CORE_DATAPATH_bkp_3__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4802_));
INVX1 INVX1_336 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4809_));
INVX1 INVX1_337 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4823_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4824_));
INVX1 INVX1_338 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4828_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4829_));
INVX1 INVX1_339 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3244_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4832_));
INVX1 INVX1_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2482_));
INVX1 INVX1_340 ( .A(AES_CORE_DATAPATH_bkp_2__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4838_));
INVX1 INVX1_341 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4845_));
INVX1 INVX1_342 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4842_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4847_));
INVX1 INVX1_343 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4858_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4859_));
INVX1 INVX1_344 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4863_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4864_));
INVX1 INVX1_345 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4867_));
INVX1 INVX1_346 ( .A(AES_CORE_DATAPATH_bkp_2__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4868_));
INVX1 INVX1_347 ( .A(AES_CORE_DATAPATH_bkp_3__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4874_));
INVX1 INVX1_348 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3266_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4883_));
INVX1 INVX1_349 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4897_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4898_));
INVX1 INVX1_35 ( .A(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2486_));
INVX1 INVX1_350 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4902_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4903_));
INVX1 INVX1_351 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3288_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4906_));
INVX1 INVX1_352 ( .A(AES_CORE_DATAPATH_bkp_2__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4912_));
INVX1 INVX1_353 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4919_));
INVX1 INVX1_354 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4916_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4921_));
INVX1 INVX1_355 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4932_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4933_));
INVX1 INVX1_356 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4937_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4938_));
INVX1 INVX1_357 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4943_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4944_));
INVX1 INVX1_358 ( .A(AES_CORE_DATAPATH_bkp_2__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4945_));
INVX1 INVX1_359 ( .A(AES_CORE_DATAPATH_bkp_3__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4951_));
INVX1 INVX1_36 ( .A(AES_CORE_DATAPATH_iv_2__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2490_));
INVX1 INVX1_360 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4969_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4970_));
INVX1 INVX1_361 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4971_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4972_));
INVX1 INVX1_362 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4976_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4977_));
INVX1 INVX1_363 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3332_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4980_));
INVX1 INVX1_364 ( .A(AES_CORE_DATAPATH_bkp_2__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4983_));
INVX1 INVX1_365 ( .A(AES_CORE_DATAPATH_bkp_3__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4989_));
INVX1 INVX1_366 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4996_));
INVX1 INVX1_367 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5010_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5011_));
INVX1 INVX1_368 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5015_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5016_));
INVX1 INVX1_369 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5021_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5022_));
INVX1 INVX1_37 ( .A(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2494_));
INVX1 INVX1_370 ( .A(AES_CORE_DATAPATH_bkp_2__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5023_));
INVX1 INVX1_371 ( .A(AES_CORE_DATAPATH_bkp_3__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5029_));
INVX1 INVX1_372 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5047_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5048_));
INVX1 INVX1_373 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5049_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5050_));
INVX1 INVX1_374 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5054_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5055_));
INVX1 INVX1_375 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3376_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5058_));
INVX1 INVX1_376 ( .A(AES_CORE_DATAPATH_bkp_2__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5061_));
INVX1 INVX1_377 ( .A(AES_CORE_DATAPATH_bkp_3__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5067_));
INVX1 INVX1_378 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5074_));
INVX1 INVX1_379 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5088_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5089_));
INVX1 INVX1_38 ( .A(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2500_));
INVX1 INVX1_380 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5093_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5094_));
INVX1 INVX1_381 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5099_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5100_));
INVX1 INVX1_382 ( .A(AES_CORE_DATAPATH_bkp_2__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5101_));
INVX1 INVX1_383 ( .A(AES_CORE_DATAPATH_bkp_3__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5107_));
INVX1 INVX1_384 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5125_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5126_));
INVX1 INVX1_385 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5127_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5128_));
INVX1 INVX1_386 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5132_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5133_));
INVX1 INVX1_387 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3420_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5136_));
INVX1 INVX1_388 ( .A(AES_CORE_DATAPATH_bkp_2__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5142_));
INVX1 INVX1_389 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5149_));
INVX1 INVX1_39 ( .A(AES_CORE_DATAPATH_iv_2__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2504_));
INVX1 INVX1_390 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5163_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5164_));
INVX1 INVX1_391 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5168_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5169_));
INVX1 INVX1_392 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5174_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5175_));
INVX1 INVX1_393 ( .A(AES_CORE_DATAPATH_bkp_2__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5176_));
INVX1 INVX1_394 ( .A(AES_CORE_DATAPATH_bkp_3__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5182_));
INVX1 INVX1_395 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5200_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5201_));
INVX1 INVX1_396 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5202_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5203_));
INVX1 INVX1_397 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5207_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5208_));
INVX1 INVX1_398 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3464_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5211_));
INVX1 INVX1_399 ( .A(AES_CORE_DATAPATH_bkp_2__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5214_));
INVX1 INVX1_4 ( .A(\aes_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_));
INVX1 INVX1_40 ( .A(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2508_));
INVX1 INVX1_400 ( .A(AES_CORE_DATAPATH_bkp_3__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5220_));
INVX1 INVX1_401 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5227_));
INVX1 INVX1_402 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5241_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5242_));
INVX1 INVX1_403 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5246_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5247_));
INVX1 INVX1_404 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5252_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5253_));
INVX1 INVX1_405 ( .A(AES_CORE_DATAPATH_bkp_2__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5254_));
INVX1 INVX1_406 ( .A(AES_CORE_DATAPATH_bkp_3__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5260_));
INVX1 INVX1_407 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5278_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5279_));
INVX1 INVX1_408 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5280_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5281_));
INVX1 INVX1_409 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5285_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5286_));
INVX1 INVX1_41 ( .A(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2514_));
INVX1 INVX1_410 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5291_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5292_));
INVX1 INVX1_411 ( .A(AES_CORE_DATAPATH_bkp_2__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5293_));
INVX1 INVX1_412 ( .A(AES_CORE_DATAPATH_bkp_3__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5299_));
INVX1 INVX1_413 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5317_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5318_));
INVX1 INVX1_414 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5319_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5320_));
INVX1 INVX1_415 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5324_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5325_));
INVX1 INVX1_416 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5330_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5331_));
INVX1 INVX1_417 ( .A(AES_CORE_DATAPATH_bkp_2__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5332_));
INVX1 INVX1_418 ( .A(AES_CORE_DATAPATH_bkp_3__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5338_));
INVX1 INVX1_419 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5356_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5357_));
INVX1 INVX1_42 ( .A(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2520_));
INVX1 INVX1_420 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5358_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5359_));
INVX1 INVX1_421 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5363_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5364_));
INVX1 INVX1_422 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3552_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5367_));
INVX1 INVX1_423 ( .A(AES_CORE_DATAPATH_bkp_2__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5370_));
INVX1 INVX1_424 ( .A(AES_CORE_DATAPATH_bkp_3__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5376_));
INVX1 INVX1_425 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5383_));
INVX1 INVX1_426 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5397_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5398_));
INVX1 INVX1_427 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5402_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5403_));
INVX1 INVX1_428 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5408_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5409_));
INVX1 INVX1_429 ( .A(AES_CORE_DATAPATH_bkp_2__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5410_));
INVX1 INVX1_43 ( .A(AES_CORE_DATAPATH_iv_1__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2521_));
INVX1 INVX1_430 ( .A(AES_CORE_DATAPATH_bkp_3__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5416_));
INVX1 INVX1_431 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5434_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5435_));
INVX1 INVX1_432 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5436_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5437_));
INVX1 INVX1_433 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5441_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5442_));
INVX1 INVX1_434 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3596_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5445_));
INVX1 INVX1_435 ( .A(AES_CORE_DATAPATH_bkp_2__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5451_));
INVX1 INVX1_436 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5458_));
INVX1 INVX1_437 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5472_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5473_));
INVX1 INVX1_438 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5477_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5478_));
INVX1 INVX1_439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5480_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5481_));
INVX1 INVX1_44 ( .A(AES_CORE_DATAPATH_iv_2__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2524_));
INVX1 INVX1_440 ( .A(AES_CORE_DATAPATH_bkp_2__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5482_));
INVX1 INVX1_441 ( .A(AES_CORE_DATAPATH_bkp_3__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5488_));
INVX1 INVX1_442 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5497_));
INVX1 INVX1_443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5511_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5512_));
INVX1 INVX1_444 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5516_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5517_));
INVX1 INVX1_445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3640_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5520_));
INVX1 INVX1_446 ( .A(AES_CORE_DATAPATH_bkp_2__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5523_));
INVX1 INVX1_447 ( .A(AES_CORE_DATAPATH_bkp_3__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5529_));
INVX1 INVX1_448 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5536_));
INVX1 INVX1_449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5550_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5551_));
INVX1 INVX1_45 ( .A(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2528_));
INVX1 INVX1_450 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5555_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5556_));
INVX1 INVX1_451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5561_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5562_));
INVX1 INVX1_452 ( .A(AES_CORE_DATAPATH_bkp_2__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5563_));
INVX1 INVX1_453 ( .A(AES_CORE_DATAPATH_bkp_3__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5569_));
INVX1 INVX1_454 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5587_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5588_));
INVX1 INVX1_455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5589_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5590_));
INVX1 INVX1_456 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5594_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5595_));
INVX1 INVX1_457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5600_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5601_));
INVX1 INVX1_458 ( .A(AES_CORE_DATAPATH_bkp_2__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5602_));
INVX1 INVX1_459 ( .A(AES_CORE_DATAPATH_bkp_3__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5608_));
INVX1 INVX1_46 ( .A(AES_CORE_DATAPATH_iv_1__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2529_));
INVX1 INVX1_460 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5627_));
INVX1 INVX1_461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5628_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5629_));
INVX1 INVX1_462 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5633_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5634_));
INVX1 INVX1_463 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3706_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5637_));
INVX1 INVX1_464 ( .A(AES_CORE_DATAPATH_bkp_2__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5640_));
INVX1 INVX1_465 ( .A(AES_CORE_DATAPATH_bkp_3__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5646_));
INVX1 INVX1_466 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5653_));
INVX1 INVX1_467 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5667_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5668_));
INVX1 INVX1_468 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5672_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5673_));
INVX1 INVX1_469 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5678_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5679_));
INVX1 INVX1_47 ( .A(AES_CORE_DATAPATH_iv_2__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2532_));
INVX1 INVX1_470 ( .A(AES_CORE_DATAPATH_bkp_2__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5680_));
INVX1 INVX1_471 ( .A(AES_CORE_DATAPATH_bkp_3__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5686_));
INVX1 INVX1_472 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5704_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5705_));
INVX1 INVX1_473 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5706_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5707_));
INVX1 INVX1_474 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5711_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5712_));
INVX1 INVX1_475 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3750_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5715_));
INVX1 INVX1_476 ( .A(AES_CORE_DATAPATH_bkp_2__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5721_));
INVX1 INVX1_477 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5728_));
INVX1 INVX1_478 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5742_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5743_));
INVX1 INVX1_479 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5747_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5748_));
INVX1 INVX1_48 ( .A(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2536_));
INVX1 INVX1_480 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3772_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5751_));
INVX1 INVX1_481 ( .A(AES_CORE_DATAPATH_bkp_2__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5754_));
INVX1 INVX1_482 ( .A(AES_CORE_DATAPATH_bkp_3__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5760_));
INVX1 INVX1_483 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5767_));
INVX1 INVX1_484 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5781_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5782_));
INVX1 INVX1_485 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5786_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5787_));
INVX1 INVX1_486 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5792_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5793_));
INVX1 INVX1_487 ( .A(AES_CORE_DATAPATH_bkp_2__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5794_));
INVX1 INVX1_488 ( .A(AES_CORE_DATAPATH_bkp_3__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5800_));
INVX1 INVX1_489 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5818_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5819_));
INVX1 INVX1_49 ( .A(AES_CORE_DATAPATH_iv_1__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2537_));
INVX1 INVX1_490 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5820_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5821_));
INVX1 INVX1_491 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6053_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6054_));
INVX1 INVX1_492 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6055_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6056_));
INVX1 INVX1_493 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6060_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6061_));
INVX1 INVX1_494 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6062_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6063_));
INVX1 INVX1_495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6067_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6068_));
INVX1 INVX1_496 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6069_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6070_));
INVX1 INVX1_497 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6074_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6075_));
INVX1 INVX1_498 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6076_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6077_));
INVX1 INVX1_499 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6081_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6082_));
INVX1 INVX1_5 ( .A(\aes_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n75_));
INVX1 INVX1_50 ( .A(AES_CORE_DATAPATH_iv_2__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2540_));
INVX1 INVX1_500 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6083_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6084_));
INVX1 INVX1_501 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6088_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6089_));
INVX1 INVX1_502 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6090_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6091_));
INVX1 INVX1_503 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6095_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6096_));
INVX1 INVX1_504 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6097_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6098_));
INVX1 INVX1_505 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6102_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6103_));
INVX1 INVX1_506 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6104_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6105_));
INVX1 INVX1_507 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6109_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6110_));
INVX1 INVX1_508 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6111_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6112_));
INVX1 INVX1_509 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6116_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6117_));
INVX1 INVX1_51 ( .A(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2544_));
INVX1 INVX1_510 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6118_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6119_));
INVX1 INVX1_511 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6123_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6124_));
INVX1 INVX1_512 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6125_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6126_));
INVX1 INVX1_513 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6130_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6131_));
INVX1 INVX1_514 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6132_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6133_));
INVX1 INVX1_515 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6137_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6138_));
INVX1 INVX1_516 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6139_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6140_));
INVX1 INVX1_517 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6144_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6145_));
INVX1 INVX1_518 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6146_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6147_));
INVX1 INVX1_519 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6151_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6152_));
INVX1 INVX1_52 ( .A(AES_CORE_DATAPATH_iv_1__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2545_));
INVX1 INVX1_520 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6153_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6154_));
INVX1 INVX1_521 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6158_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6159_));
INVX1 INVX1_522 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6160_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6161_));
INVX1 INVX1_523 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6165_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6166_));
INVX1 INVX1_524 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6167_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6168_));
INVX1 INVX1_525 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6172_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6173_));
INVX1 INVX1_526 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6174_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6175_));
INVX1 INVX1_527 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6179_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6180_));
INVX1 INVX1_528 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6181_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6182_));
INVX1 INVX1_529 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6186_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6187_));
INVX1 INVX1_53 ( .A(AES_CORE_DATAPATH_iv_2__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2548_));
INVX1 INVX1_530 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6188_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6189_));
INVX1 INVX1_531 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6193_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6194_));
INVX1 INVX1_532 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6195_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6196_));
INVX1 INVX1_533 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6200_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6201_));
INVX1 INVX1_534 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6202_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6203_));
INVX1 INVX1_535 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6207_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6208_));
INVX1 INVX1_536 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6209_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6210_));
INVX1 INVX1_537 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6214_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6215_));
INVX1 INVX1_538 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6216_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6217_));
INVX1 INVX1_539 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6221_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6222_));
INVX1 INVX1_54 ( .A(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2552_));
INVX1 INVX1_540 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6223_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6224_));
INVX1 INVX1_541 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6228_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6229_));
INVX1 INVX1_542 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6230_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6231_));
INVX1 INVX1_543 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6235_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6236_));
INVX1 INVX1_544 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6237_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6238_));
INVX1 INVX1_545 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6242_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6243_));
INVX1 INVX1_546 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6244_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6245_));
INVX1 INVX1_547 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6249_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6250_));
INVX1 INVX1_548 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6251_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6252_));
INVX1 INVX1_549 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6256_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6257_));
INVX1 INVX1_55 ( .A(AES_CORE_DATAPATH_iv_1__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2553_));
INVX1 INVX1_550 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6258_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6259_));
INVX1 INVX1_551 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6263_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6264_));
INVX1 INVX1_552 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6265_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6266_));
INVX1 INVX1_553 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6270_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6271_));
INVX1 INVX1_554 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6272_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6273_));
INVX1 INVX1_555 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6277_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6278_));
INVX1 INVX1_556 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6279_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6280_));
INVX1 INVX1_557 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6284_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6285_));
INVX1 INVX1_558 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6286_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6287_));
INVX1 INVX1_559 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6291_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6292_));
INVX1 INVX1_56 ( .A(AES_CORE_DATAPATH_iv_2__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2556_));
INVX1 INVX1_560 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6293_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6294_));
INVX1 INVX1_561 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6298_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6299_));
INVX1 INVX1_562 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6300_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6301_));
INVX1 INVX1_563 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6305_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6306_));
INVX1 INVX1_564 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6307_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6308_));
INVX1 INVX1_565 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6312_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6313_));
INVX1 INVX1_566 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6314_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6315_));
INVX1 INVX1_567 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6319_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6320_));
INVX1 INVX1_568 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6321_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6322_));
INVX1 INVX1_569 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6326_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6327_));
INVX1 INVX1_57 ( .A(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2560_));
INVX1 INVX1_570 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6328_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6329_));
INVX1 INVX1_571 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6333_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6334_));
INVX1 INVX1_572 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6335_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6336_));
INVX1 INVX1_573 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6340_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6341_));
INVX1 INVX1_574 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6342_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6343_));
INVX1 INVX1_575 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6347_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6348_));
INVX1 INVX1_576 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6349_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6350_));
INVX1 INVX1_577 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6354_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6355_));
INVX1 INVX1_578 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6356_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6357_));
INVX1 INVX1_579 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6361_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6362_));
INVX1 INVX1_58 ( .A(AES_CORE_DATAPATH_iv_1__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2561_));
INVX1 INVX1_580 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6363_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6364_));
INVX1 INVX1_581 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6368_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6369_));
INVX1 INVX1_582 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6370_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6371_));
INVX1 INVX1_583 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6375_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6376_));
INVX1 INVX1_584 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6377_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6378_));
INVX1 INVX1_585 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6382_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6383_));
INVX1 INVX1_586 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6384_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6385_));
INVX1 INVX1_587 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6389_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6390_));
INVX1 INVX1_588 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6391_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6392_));
INVX1 INVX1_589 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6396_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6397_));
INVX1 INVX1_59 ( .A(AES_CORE_DATAPATH_iv_2__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2564_));
INVX1 INVX1_590 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6398_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6399_));
INVX1 INVX1_591 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6403_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6404_));
INVX1 INVX1_592 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6405_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6406_));
INVX1 INVX1_593 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6410_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6411_));
INVX1 INVX1_594 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6412_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6413_));
INVX1 INVX1_595 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6417_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6418_));
INVX1 INVX1_596 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6419_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6420_));
INVX1 INVX1_597 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6424_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6425_));
INVX1 INVX1_598 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6426_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6427_));
INVX1 INVX1_599 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6431_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6432_));
INVX1 INVX1_6 ( .A(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_));
INVX1 INVX1_60 ( .A(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2568_));
INVX1 INVX1_600 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6433_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6434_));
INVX1 INVX1_601 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6438_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6439_));
INVX1 INVX1_602 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6440_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6441_));
INVX1 INVX1_603 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6445_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6446_));
INVX1 INVX1_604 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6447_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6448_));
INVX1 INVX1_605 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6452_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6453_));
INVX1 INVX1_606 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6454_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6455_));
INVX1 INVX1_607 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6459_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6460_));
INVX1 INVX1_608 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6462_));
INVX1 INVX1_609 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6466_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6467_));
INVX1 INVX1_61 ( .A(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2574_));
INVX1 INVX1_610 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6469_));
INVX1 INVX1_611 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6473_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6474_));
INVX1 INVX1_612 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6476_));
INVX1 INVX1_613 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6480_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6481_));
INVX1 INVX1_614 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6483_));
INVX1 INVX1_615 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6487_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6488_));
INVX1 INVX1_616 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6489_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6490_));
INVX1 INVX1_617 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6494_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6495_));
INVX1 INVX1_618 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6496_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6497_));
INVX1 INVX1_619 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6499_));
INVX1 INVX1_62 ( .A(AES_CORE_DATAPATH_iv_2__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2578_));
INVX1 INVX1_620 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6502_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6503_));
INVX1 INVX1_621 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6504_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6505_));
INVX1 INVX1_622 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6508_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6509_));
INVX1 INVX1_623 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6515_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6516_));
INVX1 INVX1_624 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6517_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6518_));
INVX1 INVX1_625 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6521_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6522_));
INVX1 INVX1_626 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6528_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6529_));
INVX1 INVX1_627 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6530_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6531_));
INVX1 INVX1_628 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6535_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6536_));
INVX1 INVX1_629 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6537_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6538_));
INVX1 INVX1_63 ( .A(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2582_));
INVX1 INVX1_630 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6542_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6543_));
INVX1 INVX1_631 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6544_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6545_));
INVX1 INVX1_632 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6548_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6549_));
INVX1 INVX1_633 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6555_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6556_));
INVX1 INVX1_634 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6557_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6558_));
INVX1 INVX1_635 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6561_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6562_));
INVX1 INVX1_636 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6568_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6569_));
INVX1 INVX1_637 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6570_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6571_));
INVX1 INVX1_638 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6574_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6575_));
INVX1 INVX1_639 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6581_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6582_));
INVX1 INVX1_64 ( .A(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2588_));
INVX1 INVX1_640 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6583_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6584_));
INVX1 INVX1_641 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6587_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6588_));
INVX1 INVX1_642 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6594_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6595_));
INVX1 INVX1_643 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6596_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6597_));
INVX1 INVX1_644 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6600_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6601_));
INVX1 INVX1_645 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6607_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6608_));
INVX1 INVX1_646 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6609_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6610_));
INVX1 INVX1_647 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6613_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6614_));
INVX1 INVX1_648 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6619_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6620_));
INVX1 INVX1_649 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6625_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6626_));
INVX1 INVX1_65 ( .A(AES_CORE_DATAPATH_iv_2__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2592_));
INVX1 INVX1_650 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6632_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6633_));
INVX1 INVX1_651 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6634_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6635_));
INVX1 INVX1_652 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6638_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6639_));
INVX1 INVX1_653 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6645_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6646_));
INVX1 INVX1_654 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6647_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6648_));
INVX1 INVX1_655 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6651_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6652_));
INVX1 INVX1_656 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6658_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6659_));
INVX1 INVX1_657 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6660_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6661_));
INVX1 INVX1_658 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6664_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6665_));
INVX1 INVX1_659 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6670_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6671_));
INVX1 INVX1_66 ( .A(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2596_));
INVX1 INVX1_660 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6677_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6678_));
INVX1 INVX1_661 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6679_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6680_));
INVX1 INVX1_662 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6683_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6684_));
INVX1 INVX1_663 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6690_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6691_));
INVX1 INVX1_664 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6692_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6693_));
INVX1 INVX1_665 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6697_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6698_));
INVX1 INVX1_666 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6699_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6700_));
INVX1 INVX1_667 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6703_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6704_));
INVX1 INVX1_668 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n6708_));
INVX1 INVX1_669 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6711_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6712_));
INVX1 INVX1_67 ( .A(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2602_));
INVX1 INVX1_670 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6710_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6778_));
INVX1 INVX1_671 ( .A(AES_CORE_DATAPATH_bkp_1_3__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6779_));
INVX1 INVX1_672 ( .A(AES_CORE_DATAPATH_bkp_1_3__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6785_));
INVX1 INVX1_673 ( .A(AES_CORE_DATAPATH_bkp_1_3__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6791_));
INVX1 INVX1_674 ( .A(AES_CORE_DATAPATH_bkp_1_3__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6797_));
INVX1 INVX1_675 ( .A(AES_CORE_DATAPATH_bkp_3__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6803_));
INVX1 INVX1_676 ( .A(AES_CORE_DATAPATH_bkp_1_3__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6804_));
INVX1 INVX1_677 ( .A(AES_CORE_DATAPATH_bkp_1_3__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6810_));
INVX1 INVX1_678 ( .A(AES_CORE_DATAPATH_bkp_3__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6816_));
INVX1 INVX1_679 ( .A(AES_CORE_DATAPATH_bkp_1_3__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6817_));
INVX1 INVX1_68 ( .A(AES_CORE_DATAPATH_iv_2__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2606_));
INVX1 INVX1_680 ( .A(AES_CORE_DATAPATH_bkp_1_3__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6823_));
INVX1 INVX1_681 ( .A(AES_CORE_DATAPATH_bkp_3__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6829_));
INVX1 INVX1_682 ( .A(AES_CORE_DATAPATH_bkp_1_3__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6830_));
INVX1 INVX1_683 ( .A(AES_CORE_DATAPATH_bkp_1_3__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6836_));
INVX1 INVX1_684 ( .A(AES_CORE_DATAPATH_bkp_1_3__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6842_));
INVX1 INVX1_685 ( .A(AES_CORE_DATAPATH_bkp_1_3__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6848_));
INVX1 INVX1_686 ( .A(AES_CORE_DATAPATH_bkp_1_3__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6854_));
INVX1 INVX1_687 ( .A(AES_CORE_DATAPATH_bkp_1_3__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6860_));
INVX1 INVX1_688 ( .A(AES_CORE_DATAPATH_bkp_3__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6866_));
INVX1 INVX1_689 ( .A(AES_CORE_DATAPATH_bkp_1_3__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6867_));
INVX1 INVX1_69 ( .A(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2610_));
INVX1 INVX1_690 ( .A(AES_CORE_DATAPATH_bkp_1_3__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6873_));
INVX1 INVX1_691 ( .A(AES_CORE_DATAPATH_bkp_1_3__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6879_));
INVX1 INVX1_692 ( .A(AES_CORE_DATAPATH_bkp_1_3__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6885_));
INVX1 INVX1_693 ( .A(AES_CORE_DATAPATH_bkp_1_3__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6891_));
INVX1 INVX1_694 ( .A(AES_CORE_DATAPATH_bkp_1_3__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6897_));
INVX1 INVX1_695 ( .A(AES_CORE_DATAPATH_bkp_1_3__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6903_));
INVX1 INVX1_696 ( .A(AES_CORE_DATAPATH_bkp_1_3__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6909_));
INVX1 INVX1_697 ( .A(AES_CORE_DATAPATH_bkp_3__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6915_));
INVX1 INVX1_698 ( .A(AES_CORE_DATAPATH_bkp_1_3__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6916_));
INVX1 INVX1_699 ( .A(AES_CORE_DATAPATH_bkp_1_3__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6922_));
INVX1 INVX1_7 ( .A(disable_core), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_));
INVX1 INVX1_70 ( .A(AES_CORE_DATAPATH_iv_2__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2614_));
INVX1 INVX1_700 ( .A(AES_CORE_DATAPATH_bkp_1_3__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6928_));
INVX1 INVX1_701 ( .A(AES_CORE_DATAPATH_bkp_1_3__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6934_));
INVX1 INVX1_702 ( .A(AES_CORE_DATAPATH_bkp_1_3__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6940_));
INVX1 INVX1_703 ( .A(AES_CORE_DATAPATH_bkp_1_3__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6946_));
INVX1 INVX1_704 ( .A(AES_CORE_DATAPATH_bkp_1_3__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6952_));
INVX1 INVX1_705 ( .A(AES_CORE_DATAPATH_bkp_3__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6958_));
INVX1 INVX1_706 ( .A(AES_CORE_DATAPATH_bkp_1_3__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6959_));
INVX1 INVX1_707 ( .A(AES_CORE_DATAPATH_bkp_1_3__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6965_));
INVX1 INVX1_708 ( .A(AES_CORE_DATAPATH_bkp_1_3__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6971_));
INVX1 INVX1_709 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6977_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6978_));
INVX1 INVX1_71 ( .A(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2618_));
INVX1 INVX1_710 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n6979_));
INVX1 INVX1_711 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6982_));
INVX1 INVX1_712 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6986_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6987_));
INVX1 INVX1_713 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6988_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6993_));
INVX1 INVX1_714 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7001_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7002_));
INVX1 INVX1_715 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7003_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7008_));
INVX1 INVX1_716 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7009_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7013_));
INVX1 INVX1_717 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7017_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7018_));
INVX1 INVX1_718 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7021_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7022_));
INVX1 INVX1_719 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7028_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7029_));
INVX1 INVX1_72 ( .A(AES_CORE_DATAPATH_iv_2__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2622_));
INVX1 INVX1_720 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7048_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7049_));
INVX1 INVX1_721 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7084_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7085_));
INVX1 INVX1_722 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7148_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7149_));
INVX1 INVX1_723 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7164_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7165_));
INVX1 INVX1_724 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7180_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7182_));
INVX1 INVX1_725 ( .A(AES_CORE_DATAPATH_bkp_1_2__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7339_));
INVX1 INVX1_726 ( .A(AES_CORE_DATAPATH_bkp_1_2__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7344_));
INVX1 INVX1_727 ( .A(AES_CORE_DATAPATH_bkp_1_2__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7349_));
INVX1 INVX1_728 ( .A(AES_CORE_DATAPATH_bkp_1_2__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7354_));
INVX1 INVX1_729 ( .A(AES_CORE_DATAPATH_bkp_1_2__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7359_));
INVX1 INVX1_73 ( .A(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2626_));
INVX1 INVX1_730 ( .A(AES_CORE_DATAPATH_bkp_1_2__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7364_));
INVX1 INVX1_731 ( .A(AES_CORE_DATAPATH_bkp_1_2__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7369_));
INVX1 INVX1_732 ( .A(AES_CORE_DATAPATH_bkp_1_2__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7374_));
INVX1 INVX1_733 ( .A(AES_CORE_DATAPATH_bkp_1_2__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7379_));
INVX1 INVX1_734 ( .A(AES_CORE_DATAPATH_bkp_1_2__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7384_));
INVX1 INVX1_735 ( .A(AES_CORE_DATAPATH_bkp_1_2__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7389_));
INVX1 INVX1_736 ( .A(AES_CORE_DATAPATH_bkp_1_2__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7394_));
INVX1 INVX1_737 ( .A(AES_CORE_DATAPATH_bkp_1_2__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7399_));
INVX1 INVX1_738 ( .A(AES_CORE_DATAPATH_bkp_1_2__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7404_));
INVX1 INVX1_739 ( .A(AES_CORE_DATAPATH_bkp_1_2__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7409_));
INVX1 INVX1_74 ( .A(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2632_));
INVX1 INVX1_740 ( .A(AES_CORE_DATAPATH_bkp_1_2__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7414_));
INVX1 INVX1_741 ( .A(AES_CORE_DATAPATH_bkp_1_2__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7419_));
INVX1 INVX1_742 ( .A(AES_CORE_DATAPATH_bkp_1_2__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7424_));
INVX1 INVX1_743 ( .A(AES_CORE_DATAPATH_bkp_1_2__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7429_));
INVX1 INVX1_744 ( .A(AES_CORE_DATAPATH_bkp_1_2__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7434_));
INVX1 INVX1_745 ( .A(AES_CORE_DATAPATH_bkp_1_2__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7439_));
INVX1 INVX1_746 ( .A(AES_CORE_DATAPATH_bkp_1_2__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7444_));
INVX1 INVX1_747 ( .A(AES_CORE_DATAPATH_bkp_1_2__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7449_));
INVX1 INVX1_748 ( .A(AES_CORE_DATAPATH_bkp_1_2__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7454_));
INVX1 INVX1_749 ( .A(AES_CORE_DATAPATH_bkp_1_2__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7459_));
INVX1 INVX1_75 ( .A(AES_CORE_DATAPATH_iv_2__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2636_));
INVX1 INVX1_750 ( .A(AES_CORE_DATAPATH_bkp_1_2__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7464_));
INVX1 INVX1_751 ( .A(AES_CORE_DATAPATH_bkp_1_2__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7469_));
INVX1 INVX1_752 ( .A(AES_CORE_DATAPATH_bkp_1_2__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7474_));
INVX1 INVX1_753 ( .A(AES_CORE_DATAPATH_bkp_1_2__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7479_));
INVX1 INVX1_754 ( .A(AES_CORE_DATAPATH_bkp_1_2__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7484_));
INVX1 INVX1_755 ( .A(AES_CORE_DATAPATH_bkp_1_2__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7489_));
INVX1 INVX1_756 ( .A(AES_CORE_DATAPATH_bkp_1_2__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7494_));
INVX1 INVX1_757 ( .A(AES_CORE_DATAPATH_bkp_1_1__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7566_));
INVX1 INVX1_758 ( .A(AES_CORE_DATAPATH_bkp_1_1__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7571_));
INVX1 INVX1_759 ( .A(AES_CORE_DATAPATH_bkp_1_1__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7580_));
INVX1 INVX1_76 ( .A(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2640_));
INVX1 INVX1_760 ( .A(AES_CORE_DATAPATH_bkp_1_1__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7585_));
INVX1 INVX1_761 ( .A(AES_CORE_DATAPATH_bkp_1_1__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7590_));
INVX1 INVX1_762 ( .A(AES_CORE_DATAPATH_bkp_1_1__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7595_));
INVX1 INVX1_763 ( .A(AES_CORE_DATAPATH_bkp_1_1__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7600_));
INVX1 INVX1_764 ( .A(AES_CORE_DATAPATH_bkp_1_1__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7605_));
INVX1 INVX1_765 ( .A(AES_CORE_DATAPATH_bkp_1_1__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7608_));
INVX1 INVX1_766 ( .A(AES_CORE_DATAPATH_bkp_1_1__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7611_));
INVX1 INVX1_767 ( .A(AES_CORE_DATAPATH_bkp_1_1__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7616_));
INVX1 INVX1_768 ( .A(AES_CORE_DATAPATH_bkp_1_1__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7621_));
INVX1 INVX1_769 ( .A(AES_CORE_DATAPATH_bkp_1_1__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7626_));
INVX1 INVX1_77 ( .A(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2646_));
INVX1 INVX1_770 ( .A(AES_CORE_DATAPATH_bkp_1_1__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7629_));
INVX1 INVX1_771 ( .A(AES_CORE_DATAPATH_bkp_1_1__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7634_));
INVX1 INVX1_772 ( .A(AES_CORE_DATAPATH_bkp_1_1__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7641_));
INVX1 INVX1_773 ( .A(AES_CORE_DATAPATH_bkp_1__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7644_));
INVX1 INVX1_774 ( .A(AES_CORE_DATAPATH_bkp_1_1__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7645_));
INVX1 INVX1_775 ( .A(AES_CORE_DATAPATH_bkp_1__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7650_));
INVX1 INVX1_776 ( .A(AES_CORE_DATAPATH_bkp_1__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7655_));
INVX1 INVX1_777 ( .A(AES_CORE_DATAPATH_bkp_1_1__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7656_));
INVX1 INVX1_778 ( .A(AES_CORE_DATAPATH_bkp_1__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7661_));
INVX1 INVX1_779 ( .A(AES_CORE_DATAPATH_bkp_1__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7666_));
INVX1 INVX1_78 ( .A(AES_CORE_DATAPATH_iv_2__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2650_));
INVX1 INVX1_780 ( .A(AES_CORE_DATAPATH_bkp_1_1__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7667_));
INVX1 INVX1_781 ( .A(AES_CORE_DATAPATH_bkp_1__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7672_));
INVX1 INVX1_782 ( .A(AES_CORE_DATAPATH_bkp_1_1__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7673_));
INVX1 INVX1_783 ( .A(AES_CORE_DATAPATH_bkp_1__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7678_));
INVX1 INVX1_784 ( .A(AES_CORE_DATAPATH_bkp_1_1__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7679_));
INVX1 INVX1_785 ( .A(AES_CORE_DATAPATH_bkp_1__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7684_));
INVX1 INVX1_786 ( .A(AES_CORE_DATAPATH_bkp_1__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7689_));
INVX1 INVX1_787 ( .A(AES_CORE_DATAPATH_bkp_1_1__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7690_));
INVX1 INVX1_788 ( .A(AES_CORE_DATAPATH_bkp_1__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7695_));
INVX1 INVX1_789 ( .A(AES_CORE_DATAPATH_bkp_1__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7700_));
INVX1 INVX1_79 ( .A(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2654_));
INVX1 INVX1_790 ( .A(AES_CORE_DATAPATH_bkp_1_1__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7701_));
INVX1 INVX1_791 ( .A(AES_CORE_DATAPATH_bkp_1__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7706_));
INVX1 INVX1_792 ( .A(AES_CORE_DATAPATH_bkp_1__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7711_));
INVX1 INVX1_793 ( .A(AES_CORE_DATAPATH_bkp_1_1__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7712_));
INVX1 INVX1_794 ( .A(AES_CORE_DATAPATH_bkp_1__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7717_));
INVX1 INVX1_795 ( .A(AES_CORE_DATAPATH_bkp_1__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7722_));
INVX1 INVX1_796 ( .A(AES_CORE_DATAPATH_bkp_1_1__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7723_));
INVX1 INVX1_797 ( .A(AES_CORE_DATAPATH_bkp_1__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7728_));
INVX1 INVX1_798 ( .A(AES_CORE_DATAPATH_bkp_1__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7733_));
INVX1 INVX1_799 ( .A(AES_CORE_DATAPATH_bkp_1_1__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7734_));
INVX1 INVX1_8 ( .A(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n89_));
INVX1 INVX1_80 ( .A(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2660_));
INVX1 INVX1_800 ( .A(AES_CORE_DATAPATH_bkp_1__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7739_));
INVX1 INVX1_801 ( .A(AES_CORE_DATAPATH_bkp_1__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7744_));
INVX1 INVX1_802 ( .A(AES_CORE_DATAPATH_bkp_1__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7749_));
INVX1 INVX1_803 ( .A(AES_CORE_DATAPATH_bkp_1__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7754_));
INVX1 INVX1_804 ( .A(AES_CORE_DATAPATH_bkp_1_1__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7755_));
INVX1 INVX1_805 ( .A(AES_CORE_DATAPATH_bkp_1__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7760_));
INVX1 INVX1_806 ( .A(AES_CORE_DATAPATH_bkp_1__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7765_));
INVX1 INVX1_807 ( .A(AES_CORE_DATAPATH_bkp_1_1__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7766_));
INVX1 INVX1_808 ( .A(AES_CORE_DATAPATH_bkp_1__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7771_));
INVX1 INVX1_809 ( .A(AES_CORE_DATAPATH_bkp_1__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7776_));
INVX1 INVX1_81 ( .A(AES_CORE_DATAPATH_iv_2__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2664_));
INVX1 INVX1_810 ( .A(AES_CORE_DATAPATH_bkp_1_1__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7777_));
INVX1 INVX1_811 ( .A(AES_CORE_DATAPATH_bkp_1__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7782_));
INVX1 INVX1_812 ( .A(AES_CORE_DATAPATH_bkp_1__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7787_));
INVX1 INVX1_813 ( .A(AES_CORE_DATAPATH_bkp_1__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7792_));
INVX1 INVX1_814 ( .A(AES_CORE_DATAPATH_bkp_1_1__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7793_));
INVX1 INVX1_815 ( .A(AES_CORE_DATAPATH_bkp_1__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7798_));
INVX1 INVX1_816 ( .A(AES_CORE_DATAPATH_bkp_1__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7803_));
INVX1 INVX1_817 ( .A(AES_CORE_DATAPATH_bkp_1_1__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7804_));
INVX1 INVX1_818 ( .A(AES_CORE_DATAPATH_bkp_1__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7809_));
INVX1 INVX1_819 ( .A(AES_CORE_DATAPATH_bkp_1_1__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7810_));
INVX1 INVX1_82 ( .A(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2668_));
INVX1 INVX1_820 ( .A(AES_CORE_DATAPATH_bkp_1__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7815_));
INVX1 INVX1_821 ( .A(AES_CORE_DATAPATH_iv_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7832_));
INVX1 INVX1_822 ( .A(AES_CORE_DATAPATH_iv_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7835_));
INVX1 INVX1_823 ( .A(AES_CORE_DATAPATH_iv_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7838_));
INVX1 INVX1_824 ( .A(AES_CORE_DATAPATH_iv_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7841_));
INVX1 INVX1_825 ( .A(AES_CORE_DATAPATH_iv_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7844_));
INVX1 INVX1_826 ( .A(AES_CORE_DATAPATH_iv_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7847_));
INVX1 INVX1_827 ( .A(AES_CORE_DATAPATH_bkp_0__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7955_));
INVX1 INVX1_828 ( .A(AES_CORE_DATAPATH_bkp_1_0__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7956_));
INVX1 INVX1_829 ( .A(AES_CORE_DATAPATH_bkp_0__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7961_));
INVX1 INVX1_83 ( .A(AES_CORE_DATAPATH_iv_2__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2672_));
INVX1 INVX1_830 ( .A(AES_CORE_DATAPATH_bkp_1_0__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7962_));
INVX1 INVX1_831 ( .A(AES_CORE_DATAPATH_bkp_0__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7967_));
INVX1 INVX1_832 ( .A(AES_CORE_DATAPATH_bkp_1_0__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7968_));
INVX1 INVX1_833 ( .A(AES_CORE_DATAPATH_bkp_0__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7973_));
INVX1 INVX1_834 ( .A(AES_CORE_DATAPATH_bkp_1_0__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7974_));
INVX1 INVX1_835 ( .A(AES_CORE_DATAPATH_bkp_0__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7979_));
INVX1 INVX1_836 ( .A(AES_CORE_DATAPATH_bkp_1_0__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7980_));
INVX1 INVX1_837 ( .A(AES_CORE_DATAPATH_bkp_0__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7985_));
INVX1 INVX1_838 ( .A(AES_CORE_DATAPATH_bkp_1_0__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7986_));
INVX1 INVX1_839 ( .A(AES_CORE_DATAPATH_bkp_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7991_));
INVX1 INVX1_84 ( .A(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2676_));
INVX1 INVX1_840 ( .A(AES_CORE_DATAPATH_bkp_1_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7992_));
INVX1 INVX1_841 ( .A(AES_CORE_DATAPATH_bkp_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7997_));
INVX1 INVX1_842 ( .A(AES_CORE_DATAPATH_bkp_1_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7998_));
INVX1 INVX1_843 ( .A(AES_CORE_DATAPATH_bkp_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8003_));
INVX1 INVX1_844 ( .A(AES_CORE_DATAPATH_bkp_1_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8004_));
INVX1 INVX1_845 ( .A(AES_CORE_DATAPATH_bkp_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8009_));
INVX1 INVX1_846 ( .A(AES_CORE_DATAPATH_bkp_1_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8010_));
INVX1 INVX1_847 ( .A(AES_CORE_DATAPATH_bkp_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8015_));
INVX1 INVX1_848 ( .A(AES_CORE_DATAPATH_bkp_1_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8016_));
INVX1 INVX1_849 ( .A(AES_CORE_DATAPATH_bkp_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8021_));
INVX1 INVX1_85 ( .A(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2682_));
INVX1 INVX1_850 ( .A(AES_CORE_DATAPATH_bkp_1_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8022_));
INVX1 INVX1_851 ( .A(AES_CORE_DATAPATH_bkp_0__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8027_));
INVX1 INVX1_852 ( .A(AES_CORE_DATAPATH_bkp_1_0__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8028_));
INVX1 INVX1_853 ( .A(AES_CORE_DATAPATH_bkp_0__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8033_));
INVX1 INVX1_854 ( .A(AES_CORE_DATAPATH_bkp_1_0__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8034_));
INVX1 INVX1_855 ( .A(AES_CORE_DATAPATH_bkp_0__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8039_));
INVX1 INVX1_856 ( .A(AES_CORE_DATAPATH_bkp_1_0__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8040_));
INVX1 INVX1_857 ( .A(AES_CORE_DATAPATH_bkp_0__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8045_));
INVX1 INVX1_858 ( .A(AES_CORE_DATAPATH_bkp_1_0__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8046_));
INVX1 INVX1_859 ( .A(AES_CORE_DATAPATH_bkp_0__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8051_));
INVX1 INVX1_86 ( .A(AES_CORE_DATAPATH_iv_2__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2686_));
INVX1 INVX1_860 ( .A(AES_CORE_DATAPATH_bkp_1_0__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8052_));
INVX1 INVX1_861 ( .A(AES_CORE_DATAPATH_bkp_0__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8057_));
INVX1 INVX1_862 ( .A(AES_CORE_DATAPATH_bkp_1_0__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8058_));
INVX1 INVX1_863 ( .A(AES_CORE_DATAPATH_bkp_0__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8063_));
INVX1 INVX1_864 ( .A(AES_CORE_DATAPATH_bkp_1_0__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8064_));
INVX1 INVX1_865 ( .A(AES_CORE_DATAPATH_bkp_0__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8069_));
INVX1 INVX1_866 ( .A(AES_CORE_DATAPATH_bkp_1_0__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8070_));
INVX1 INVX1_867 ( .A(AES_CORE_DATAPATH_bkp_0__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8075_));
INVX1 INVX1_868 ( .A(AES_CORE_DATAPATH_bkp_1_0__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8076_));
INVX1 INVX1_869 ( .A(AES_CORE_DATAPATH_bkp_0__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8081_));
INVX1 INVX1_87 ( .A(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2690_));
INVX1 INVX1_870 ( .A(AES_CORE_DATAPATH_bkp_1_0__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8082_));
INVX1 INVX1_871 ( .A(AES_CORE_DATAPATH_bkp_0__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8087_));
INVX1 INVX1_872 ( .A(AES_CORE_DATAPATH_bkp_1_0__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8088_));
INVX1 INVX1_873 ( .A(AES_CORE_DATAPATH_bkp_0__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8093_));
INVX1 INVX1_874 ( .A(AES_CORE_DATAPATH_bkp_1_0__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8094_));
INVX1 INVX1_875 ( .A(AES_CORE_DATAPATH_bkp_0__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8099_));
INVX1 INVX1_876 ( .A(AES_CORE_DATAPATH_bkp_1_0__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8100_));
INVX1 INVX1_877 ( .A(AES_CORE_DATAPATH_bkp_0__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8105_));
INVX1 INVX1_878 ( .A(AES_CORE_DATAPATH_bkp_1_0__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8106_));
INVX1 INVX1_879 ( .A(AES_CORE_DATAPATH_bkp_0__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8111_));
INVX1 INVX1_88 ( .A(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2696_));
INVX1 INVX1_880 ( .A(AES_CORE_DATAPATH_bkp_1_0__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8112_));
INVX1 INVX1_881 ( .A(AES_CORE_DATAPATH_bkp_0__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8117_));
INVX1 INVX1_882 ( .A(AES_CORE_DATAPATH_bkp_1_0__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8118_));
INVX1 INVX1_883 ( .A(AES_CORE_DATAPATH_bkp_0__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8123_));
INVX1 INVX1_884 ( .A(AES_CORE_DATAPATH_bkp_1_0__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8124_));
INVX1 INVX1_885 ( .A(AES_CORE_DATAPATH_bkp_0__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8129_));
INVX1 INVX1_886 ( .A(AES_CORE_DATAPATH_bkp_1_0__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8130_));
INVX1 INVX1_887 ( .A(AES_CORE_DATAPATH_bkp_0__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8135_));
INVX1 INVX1_888 ( .A(AES_CORE_DATAPATH_bkp_1_0__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8136_));
INVX1 INVX1_889 ( .A(AES_CORE_DATAPATH_bkp_0__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8141_));
INVX1 INVX1_89 ( .A(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2702_));
INVX1 INVX1_890 ( .A(AES_CORE_DATAPATH_bkp_1_0__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8142_));
INVX1 INVX1_891 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8147_));
INVX1 INVX1_892 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8150_));
INVX1 INVX1_893 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8153_));
INVX1 INVX1_894 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8156_));
INVX1 INVX1_895 ( .A(AES_CORE_CONTROL_UNIT_key_en_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8161_));
INVX1 INVX1_896 ( .A(AES_CORE_CONTROL_UNIT_key_en_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8164_));
INVX1 INVX1_897 ( .A(AES_CORE_CONTROL_UNIT_key_en_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8167_));
INVX1 INVX1_898 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2740_), .Y(\key_out[0] ));
INVX1 INVX1_899 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2764_), .Y(\key_out[2] ));
INVX1 INVX1_9 ( .A(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n102_));
INVX1 INVX1_90 ( .A(AES_CORE_DATAPATH_iv_2__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2706_));
INVX1 INVX1_900 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2774_), .Y(\key_out[3] ));
INVX1 INVX1_901 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2784_), .Y(\key_out[4] ));
INVX1 INVX1_902 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2794_), .Y(\key_out[5] ));
INVX1 INVX1_903 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2804_), .Y(\key_out[6] ));
INVX1 INVX1_904 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2840_), .Y(\key_out[9] ));
INVX1 INVX1_905 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2851_), .Y(\key_out[10] ));
INVX1 INVX1_906 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2860_), .Y(\key_out[11] ));
INVX1 INVX1_907 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2870_), .Y(\key_out[12] ));
INVX1 INVX1_908 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2880_), .Y(\key_out[13] ));
INVX1 INVX1_909 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2890_), .Y(\key_out[14] ));
INVX1 INVX1_91 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2711_));
INVX1 INVX1_910 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2900_), .Y(\key_out[15] ));
INVX1 INVX1_911 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2911_), .Y(\key_out[16] ));
INVX1 INVX1_912 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2920_), .Y(\key_out[17] ));
INVX1 INVX1_913 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2930_), .Y(\key_out[18] ));
INVX1 INVX1_914 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2940_), .Y(\key_out[19] ));
INVX1 INVX1_915 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2963_), .Y(\key_out[21] ));
INVX1 INVX1_916 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2973_), .Y(\key_out[22] ));
INVX1 INVX1_917 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3009_), .Y(\key_out[25] ));
INVX1 INVX1_918 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3019_), .Y(\key_out[26] ));
INVX1 INVX1_919 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3029_), .Y(\key_out[27] ));
INVX1 INVX1_92 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n2712_));
INVX1 INVX1_920 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3040_), .Y(\key_out[28] ));
INVX1 INVX1_921 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3050_), .Y(\key_out[29] ));
INVX1 INVX1_922 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3060_), .Y(\key_out[30] ));
INVX1 INVX1_923 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3069_), .Y(\key_out[31] ));
INVX1 INVX1_924 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n400_));
INVX1 INVX1_925 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n401_));
INVX1 INVX1_926 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_));
INVX1 INVX1_927 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_));
INVX1 INVX1_928 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n421_));
INVX1 INVX1_929 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n413_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n422_));
INVX1 INVX1_93 ( .A(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2713_));
INVX1 INVX1_930 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_));
INVX1 INVX1_931 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n431_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n432_));
INVX1 INVX1_932 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n433_));
INVX1 INVX1_933 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n406_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n439_));
INVX1 INVX1_934 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n456_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n457_));
INVX1 INVX1_935 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n458_));
INVX1 INVX1_936 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n481_));
INVX1 INVX1_937 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n475_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n489_));
INVX1 INVX1_938 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n493_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n494_));
INVX1 INVX1_939 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n495_));
INVX1 INVX1_94 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n2715_));
INVX1 INVX1_940 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n513_));
INVX1 INVX1_941 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n522_));
INVX1 INVX1_942 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n528_));
INVX1 INVX1_943 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n532_));
INVX1 INVX1_944 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n536_));
INVX1 INVX1_945 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n540_));
INVX1 INVX1_946 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n544_));
INVX1 INVX1_947 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n548_));
INVX1 INVX1_948 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n552_));
INVX1 INVX1_949 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n556_));
INVX1 INVX1_95 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n2716_));
INVX1 INVX1_950 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n560_));
INVX1 INVX1_951 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n564_));
INVX1 INVX1_952 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n568_));
INVX1 INVX1_953 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n572_));
INVX1 INVX1_954 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n576_));
INVX1 INVX1_955 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n580_));
INVX1 INVX1_956 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n584_));
INVX1 INVX1_957 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n588_));
INVX1 INVX1_958 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n592_));
INVX1 INVX1_959 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n596_));
INVX1 INVX1_96 ( .A(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2717_));
INVX1 INVX1_960 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n600_));
INVX1 INVX1_961 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n604_));
INVX1 INVX1_962 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n608_));
INVX1 INVX1_963 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n612_));
INVX1 INVX1_964 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n616_));
INVX1 INVX1_965 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n620_));
INVX1 INVX1_966 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n624_));
INVX1 INVX1_967 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n628_));
INVX1 INVX1_968 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n632_));
INVX1 INVX1_969 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n636_));
INVX1 INVX1_97 ( .A(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2722_));
INVX1 INVX1_970 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n640_));
INVX1 INVX1_971 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n644_));
INVX1 INVX1_972 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n648_));
INVX1 INVX1_973 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n652_));
INVX1 INVX1_974 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n683_));
INVX1 INVX1_975 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n689_));
INVX1 INVX1_976 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n107_));
INVX1 INVX1_977 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n114_));
INVX1 INVX1_978 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n116_));
INVX1 INVX1_979 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n128_));
INVX1 INVX1_98 ( .A(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2724_));
INVX1 INVX1_980 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n130_));
INVX1 INVX1_981 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_));
INVX1 INVX1_982 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n171_));
INVX1 INVX1_983 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n177_));
INVX1 INVX1_984 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n178_));
INVX1 INVX1_985 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n214_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n215_));
INVX1 INVX1_986 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n217_));
INVX1 INVX1_987 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n219_));
INVX1 INVX1_988 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n222_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n223_));
INVX1 INVX1_989 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n240_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n242_));
INVX1 INVX1_99 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2720_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2734_));
INVX1 INVX1_990 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n247_));
INVX1 INVX1_991 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n249_));
INVX1 INVX1_992 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n256_));
INVX1 INVX1_993 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n292_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_));
INVX1 INVX1_994 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n294_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n296_));
INVX1 INVX1_995 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n299_));
INVX1 INVX1_996 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n326_));
INVX1 INVX1_997 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n333_));
INVX1 INVX1_998 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n345_));
INVX1 INVX1_999 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n346_));
MUX2X1 MUX2X1_1 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2469_), .B(AES_CORE_DATAPATH__abc_15863_new_n2479_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2480_));
MUX2X1 MUX2X1_10 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2561_), .B(AES_CORE_DATAPATH__abc_15863_new_n2562_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2563_));
MUX2X1 MUX2X1_100 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4120_), .B(AES_CORE_DATAPATH__abc_15863_new_n2914_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__17_));
MUX2X1 MUX2X1_101 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4125_), .B(AES_CORE_DATAPATH__abc_15863_new_n2924_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__18_));
MUX2X1 MUX2X1_102 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4130_), .B(AES_CORE_DATAPATH__abc_15863_new_n2934_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__19_));
MUX2X1 MUX2X1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4135_), .B(AES_CORE_DATAPATH__abc_15863_new_n2945_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__20_));
MUX2X1 MUX2X1_104 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4140_), .B(AES_CORE_DATAPATH__abc_15863_new_n2957_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__21_));
MUX2X1 MUX2X1_105 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4145_), .B(AES_CORE_DATAPATH__abc_15863_new_n2967_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__22_));
MUX2X1 MUX2X1_106 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4150_), .B(AES_CORE_DATAPATH__abc_15863_new_n2978_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__23_));
MUX2X1 MUX2X1_107 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4155_), .B(AES_CORE_DATAPATH__abc_15863_new_n2995_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__24_));
MUX2X1 MUX2X1_108 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4160_), .B(AES_CORE_DATAPATH__abc_15863_new_n3007_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__25_));
MUX2X1 MUX2X1_109 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4165_), .B(AES_CORE_DATAPATH__abc_15863_new_n3017_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__26_));
MUX2X1 MUX2X1_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2572_), .B(AES_CORE_DATAPATH__abc_15863_new_n2568_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[12] ));
MUX2X1 MUX2X1_110 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4170_), .B(AES_CORE_DATAPATH__abc_15863_new_n3027_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__27_));
MUX2X1 MUX2X1_111 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4175_), .B(AES_CORE_DATAPATH__abc_15863_new_n3038_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__28_));
MUX2X1 MUX2X1_112 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4180_), .B(AES_CORE_DATAPATH__abc_15863_new_n3048_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__29_));
MUX2X1 MUX2X1_113 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4185_), .B(AES_CORE_DATAPATH__abc_15863_new_n3058_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__30_));
MUX2X1 MUX2X1_114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4191_), .B(AES_CORE_DATAPATH__abc_15863_new_n3063_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__31_));
MUX2X1 MUX2X1_115 ( .A(\bus_in[6] ), .B(AES_CORE_DATAPATH_key_host_2__6_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4261_));
MUX2X1 MUX2X1_116 ( .A(\bus_in[7] ), .B(AES_CORE_DATAPATH_key_host_2__7_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4264_));
MUX2X1 MUX2X1_117 ( .A(\bus_in[8] ), .B(AES_CORE_DATAPATH_key_host_2__8_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4267_));
MUX2X1 MUX2X1_118 ( .A(\bus_in[9] ), .B(AES_CORE_DATAPATH_key_host_2__9_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4270_));
MUX2X1 MUX2X1_119 ( .A(\bus_in[10] ), .B(AES_CORE_DATAPATH_key_host_2__10_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4273_));
MUX2X1 MUX2X1_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2586_), .B(AES_CORE_DATAPATH__abc_15863_new_n2582_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[14] ));
MUX2X1 MUX2X1_120 ( .A(\bus_in[11] ), .B(AES_CORE_DATAPATH_key_host_2__11_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4276_));
MUX2X1 MUX2X1_121 ( .A(\bus_in[31] ), .B(AES_CORE_DATAPATH_key_host_2__31_), .S(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4373_));
MUX2X1 MUX2X1_122 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4581_));
MUX2X1 MUX2X1_123 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4634_));
MUX2X1 MUX2X1_124 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4673_));
MUX2X1 MUX2X1_125 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4712_));
MUX2X1 MUX2X1_126 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4752_));
MUX2X1 MUX2X1_127 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4788_));
MUX2X1 MUX2X1_128 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4827_));
MUX2X1 MUX2X1_129 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4862_));
MUX2X1 MUX2X1_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2600_), .B(AES_CORE_DATAPATH__abc_15863_new_n2596_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[16] ));
MUX2X1 MUX2X1_130 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4901_));
MUX2X1 MUX2X1_131 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4936_));
MUX2X1 MUX2X1_132 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n4975_));
MUX2X1 MUX2X1_133 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5014_));
MUX2X1 MUX2X1_134 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5053_));
MUX2X1 MUX2X1_135 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5092_));
MUX2X1 MUX2X1_136 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5131_));
MUX2X1 MUX2X1_137 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5167_));
MUX2X1 MUX2X1_138 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5206_));
MUX2X1 MUX2X1_139 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5245_));
MUX2X1 MUX2X1_14 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2630_), .B(AES_CORE_DATAPATH__abc_15863_new_n2626_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[20] ));
MUX2X1 MUX2X1_140 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5284_));
MUX2X1 MUX2X1_141 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5323_));
MUX2X1 MUX2X1_142 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5362_));
MUX2X1 MUX2X1_143 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5401_));
MUX2X1 MUX2X1_144 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5440_));
MUX2X1 MUX2X1_145 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5476_));
MUX2X1 MUX2X1_146 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5515_));
MUX2X1 MUX2X1_147 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5554_));
MUX2X1 MUX2X1_148 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5593_));
MUX2X1 MUX2X1_149 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5632_));
MUX2X1 MUX2X1_15 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2644_), .B(AES_CORE_DATAPATH__abc_15863_new_n2640_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[22] ));
MUX2X1 MUX2X1_150 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5671_));
MUX2X1 MUX2X1_151 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5710_));
MUX2X1 MUX2X1_152 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5746_));
MUX2X1 MUX2X1_153 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n5785_));
MUX2X1 MUX2X1_154 ( .A(\bus_in[0] ), .B(AES_CORE_DATAPATH_key_host_3__0_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5826_));
MUX2X1 MUX2X1_155 ( .A(\bus_in[1] ), .B(AES_CORE_DATAPATH_key_host_3__1_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5831_));
MUX2X1 MUX2X1_156 ( .A(\bus_in[2] ), .B(AES_CORE_DATAPATH_key_host_3__2_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5836_));
MUX2X1 MUX2X1_157 ( .A(\bus_in[3] ), .B(AES_CORE_DATAPATH_key_host_3__3_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5841_));
MUX2X1 MUX2X1_158 ( .A(\bus_in[4] ), .B(AES_CORE_DATAPATH_key_host_3__4_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5846_));
MUX2X1 MUX2X1_159 ( .A(\bus_in[5] ), .B(AES_CORE_DATAPATH_key_host_3__5_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5851_));
MUX2X1 MUX2X1_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2658_), .B(AES_CORE_DATAPATH__abc_15863_new_n2654_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[24] ));
MUX2X1 MUX2X1_160 ( .A(\bus_in[6] ), .B(AES_CORE_DATAPATH_key_host_3__6_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5856_));
MUX2X1 MUX2X1_161 ( .A(\bus_in[7] ), .B(AES_CORE_DATAPATH_key_host_3__7_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5861_));
MUX2X1 MUX2X1_162 ( .A(\bus_in[8] ), .B(AES_CORE_DATAPATH_key_host_3__8_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5866_));
MUX2X1 MUX2X1_163 ( .A(\bus_in[9] ), .B(AES_CORE_DATAPATH_key_host_3__9_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5871_));
MUX2X1 MUX2X1_164 ( .A(\bus_in[10] ), .B(AES_CORE_DATAPATH_key_host_3__10_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5876_));
MUX2X1 MUX2X1_165 ( .A(\bus_in[11] ), .B(AES_CORE_DATAPATH_key_host_3__11_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5881_));
MUX2X1 MUX2X1_166 ( .A(\bus_in[12] ), .B(AES_CORE_DATAPATH_key_host_3__12_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5886_));
MUX2X1 MUX2X1_167 ( .A(\bus_in[13] ), .B(AES_CORE_DATAPATH_key_host_3__13_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5891_));
MUX2X1 MUX2X1_168 ( .A(\bus_in[14] ), .B(AES_CORE_DATAPATH_key_host_3__14_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5896_));
MUX2X1 MUX2X1_169 ( .A(\bus_in[15] ), .B(AES_CORE_DATAPATH_key_host_3__15_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5901_));
MUX2X1 MUX2X1_17 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2680_), .B(AES_CORE_DATAPATH__abc_15863_new_n2676_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[27] ));
MUX2X1 MUX2X1_170 ( .A(\bus_in[16] ), .B(AES_CORE_DATAPATH_key_host_3__16_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5906_));
MUX2X1 MUX2X1_171 ( .A(\bus_in[17] ), .B(AES_CORE_DATAPATH_key_host_3__17_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5911_));
MUX2X1 MUX2X1_172 ( .A(\bus_in[18] ), .B(AES_CORE_DATAPATH_key_host_3__18_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5916_));
MUX2X1 MUX2X1_173 ( .A(\bus_in[19] ), .B(AES_CORE_DATAPATH_key_host_3__19_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5921_));
MUX2X1 MUX2X1_174 ( .A(\bus_in[20] ), .B(AES_CORE_DATAPATH_key_host_3__20_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5926_));
MUX2X1 MUX2X1_175 ( .A(\bus_in[21] ), .B(AES_CORE_DATAPATH_key_host_3__21_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5931_));
MUX2X1 MUX2X1_176 ( .A(\bus_in[22] ), .B(AES_CORE_DATAPATH_key_host_3__22_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5936_));
MUX2X1 MUX2X1_177 ( .A(\bus_in[23] ), .B(AES_CORE_DATAPATH_key_host_3__23_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5941_));
MUX2X1 MUX2X1_178 ( .A(\bus_in[24] ), .B(AES_CORE_DATAPATH_key_host_3__24_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5946_));
MUX2X1 MUX2X1_179 ( .A(\bus_in[25] ), .B(AES_CORE_DATAPATH_key_host_3__25_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5951_));
MUX2X1 MUX2X1_18 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2694_), .B(AES_CORE_DATAPATH__abc_15863_new_n2690_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[29] ));
MUX2X1 MUX2X1_180 ( .A(\bus_in[26] ), .B(AES_CORE_DATAPATH_key_host_3__26_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5956_));
MUX2X1 MUX2X1_181 ( .A(\bus_in[27] ), .B(AES_CORE_DATAPATH_key_host_3__27_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5961_));
MUX2X1 MUX2X1_182 ( .A(\bus_in[28] ), .B(AES_CORE_DATAPATH_key_host_3__28_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5966_));
MUX2X1 MUX2X1_183 ( .A(\bus_in[29] ), .B(AES_CORE_DATAPATH_key_host_3__29_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5971_));
MUX2X1 MUX2X1_184 ( .A(\bus_in[30] ), .B(AES_CORE_DATAPATH_key_host_3__30_), .S(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5976_));
MUX2X1 MUX2X1_185 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6052_));
MUX2X1 MUX2X1_186 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6059_));
MUX2X1 MUX2X1_187 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6066_));
MUX2X1 MUX2X1_188 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6073_));
MUX2X1 MUX2X1_189 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6080_));
MUX2X1 MUX2X1_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2700_), .B(AES_CORE_DATAPATH__abc_15863_new_n2696_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[30] ));
MUX2X1 MUX2X1_190 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6087_));
MUX2X1 MUX2X1_191 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6094_));
MUX2X1 MUX2X1_192 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6101_));
MUX2X1 MUX2X1_193 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6108_));
MUX2X1 MUX2X1_194 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6115_));
MUX2X1 MUX2X1_195 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6122_));
MUX2X1 MUX2X1_196 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6129_));
MUX2X1 MUX2X1_197 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6136_));
MUX2X1 MUX2X1_198 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6143_));
MUX2X1 MUX2X1_199 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6150_));
MUX2X1 MUX2X1_2 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2498_), .B(AES_CORE_DATAPATH__abc_15863_new_n2494_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[2] ));
MUX2X1 MUX2X1_20 ( .A(AES_CORE_CONTROL_UNIT_key_sel), .B(AES_CORE_DATAPATH_key_sel_pp1), .S(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n3867_));
MUX2X1 MUX2X1_200 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6157_));
MUX2X1 MUX2X1_201 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6164_));
MUX2X1 MUX2X1_202 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6171_));
MUX2X1 MUX2X1_203 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6178_));
MUX2X1 MUX2X1_204 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6185_));
MUX2X1 MUX2X1_205 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6192_));
MUX2X1 MUX2X1_206 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6199_));
MUX2X1 MUX2X1_207 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6206_));
MUX2X1 MUX2X1_208 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6213_));
MUX2X1 MUX2X1_209 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6220_));
MUX2X1 MUX2X1_21 ( .A(\bus_in[0] ), .B(AES_CORE_DATAPATH_key_host_1__0_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3868_));
MUX2X1 MUX2X1_210 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6227_));
MUX2X1 MUX2X1_211 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6234_));
MUX2X1 MUX2X1_212 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6241_));
MUX2X1 MUX2X1_213 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6248_));
MUX2X1 MUX2X1_214 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6255_));
MUX2X1 MUX2X1_215 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6262_));
MUX2X1 MUX2X1_216 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6269_));
MUX2X1 MUX2X1_217 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6276_));
MUX2X1 MUX2X1_218 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6283_));
MUX2X1 MUX2X1_219 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6290_));
MUX2X1 MUX2X1_22 ( .A(\bus_in[1] ), .B(AES_CORE_DATAPATH_key_host_1__1_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3873_));
MUX2X1 MUX2X1_220 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6297_));
MUX2X1 MUX2X1_221 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6304_));
MUX2X1 MUX2X1_222 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6311_));
MUX2X1 MUX2X1_223 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6318_));
MUX2X1 MUX2X1_224 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6325_));
MUX2X1 MUX2X1_225 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6332_));
MUX2X1 MUX2X1_226 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6339_));
MUX2X1 MUX2X1_227 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6346_));
MUX2X1 MUX2X1_228 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6353_));
MUX2X1 MUX2X1_229 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6360_));
MUX2X1 MUX2X1_23 ( .A(\bus_in[2] ), .B(AES_CORE_DATAPATH_key_host_1__2_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3878_));
MUX2X1 MUX2X1_230 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6367_));
MUX2X1 MUX2X1_231 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6374_));
MUX2X1 MUX2X1_232 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6381_));
MUX2X1 MUX2X1_233 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6388_));
MUX2X1 MUX2X1_234 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6395_));
MUX2X1 MUX2X1_235 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6402_));
MUX2X1 MUX2X1_236 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6409_));
MUX2X1 MUX2X1_237 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6416_));
MUX2X1 MUX2X1_238 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6423_));
MUX2X1 MUX2X1_239 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6430_));
MUX2X1 MUX2X1_24 ( .A(\bus_in[3] ), .B(AES_CORE_DATAPATH_key_host_1__3_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3883_));
MUX2X1 MUX2X1_240 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6437_));
MUX2X1 MUX2X1_241 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6444_));
MUX2X1 MUX2X1_242 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6451_));
MUX2X1 MUX2X1_243 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6458_));
MUX2X1 MUX2X1_244 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6465_));
MUX2X1 MUX2X1_245 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6472_));
MUX2X1 MUX2X1_246 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6479_));
MUX2X1 MUX2X1_247 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6486_));
MUX2X1 MUX2X1_248 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6493_));
MUX2X1 MUX2X1_249 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6501_));
MUX2X1 MUX2X1_25 ( .A(\bus_in[4] ), .B(AES_CORE_DATAPATH_key_host_1__4_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3888_));
MUX2X1 MUX2X1_250 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6507_));
MUX2X1 MUX2X1_251 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6514_));
MUX2X1 MUX2X1_252 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6520_));
MUX2X1 MUX2X1_253 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6527_));
MUX2X1 MUX2X1_254 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6534_));
MUX2X1 MUX2X1_255 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6541_));
MUX2X1 MUX2X1_256 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6547_));
MUX2X1 MUX2X1_257 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6554_));
MUX2X1 MUX2X1_258 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6560_));
MUX2X1 MUX2X1_259 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6567_));
MUX2X1 MUX2X1_26 ( .A(\bus_in[5] ), .B(AES_CORE_DATAPATH_key_host_1__5_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3893_));
MUX2X1 MUX2X1_260 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6573_));
MUX2X1 MUX2X1_261 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6580_));
MUX2X1 MUX2X1_262 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6586_));
MUX2X1 MUX2X1_263 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6593_));
MUX2X1 MUX2X1_264 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6599_));
MUX2X1 MUX2X1_265 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6606_));
MUX2X1 MUX2X1_266 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6612_));
MUX2X1 MUX2X1_267 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6618_));
MUX2X1 MUX2X1_268 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6624_));
MUX2X1 MUX2X1_269 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6631_));
MUX2X1 MUX2X1_27 ( .A(\bus_in[6] ), .B(AES_CORE_DATAPATH_key_host_1__6_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3898_));
MUX2X1 MUX2X1_270 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6637_));
MUX2X1 MUX2X1_271 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6644_));
MUX2X1 MUX2X1_272 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6650_));
MUX2X1 MUX2X1_273 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6657_));
MUX2X1 MUX2X1_274 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6663_));
MUX2X1 MUX2X1_275 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6669_));
MUX2X1 MUX2X1_276 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6676_));
MUX2X1 MUX2X1_277 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6682_));
MUX2X1 MUX2X1_278 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6689_));
MUX2X1 MUX2X1_279 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6696_));
MUX2X1 MUX2X1_28 ( .A(\bus_in[7] ), .B(AES_CORE_DATAPATH_key_host_1__7_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3903_));
MUX2X1 MUX2X1_280 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .S(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_15863_new_n6702_));
MUX2X1 MUX2X1_29 ( .A(\bus_in[8] ), .B(AES_CORE_DATAPATH_key_host_1__8_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3908_));
MUX2X1 MUX2X1_3 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2512_), .B(AES_CORE_DATAPATH__abc_15863_new_n2508_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[4] ));
MUX2X1 MUX2X1_30 ( .A(\bus_in[9] ), .B(AES_CORE_DATAPATH_key_host_1__9_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3913_));
MUX2X1 MUX2X1_31 ( .A(\bus_in[10] ), .B(AES_CORE_DATAPATH_key_host_1__10_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3918_));
MUX2X1 MUX2X1_32 ( .A(\bus_in[11] ), .B(AES_CORE_DATAPATH_key_host_1__11_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3923_));
MUX2X1 MUX2X1_33 ( .A(\bus_in[12] ), .B(AES_CORE_DATAPATH_key_host_1__12_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3928_));
MUX2X1 MUX2X1_34 ( .A(\bus_in[13] ), .B(AES_CORE_DATAPATH_key_host_1__13_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3933_));
MUX2X1 MUX2X1_35 ( .A(\bus_in[14] ), .B(AES_CORE_DATAPATH_key_host_1__14_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3938_));
MUX2X1 MUX2X1_36 ( .A(\bus_in[15] ), .B(AES_CORE_DATAPATH_key_host_1__15_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3943_));
MUX2X1 MUX2X1_37 ( .A(\bus_in[16] ), .B(AES_CORE_DATAPATH_key_host_1__16_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3948_));
MUX2X1 MUX2X1_38 ( .A(\bus_in[17] ), .B(AES_CORE_DATAPATH_key_host_1__17_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3953_));
MUX2X1 MUX2X1_39 ( .A(\bus_in[18] ), .B(AES_CORE_DATAPATH_key_host_1__18_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3958_));
MUX2X1 MUX2X1_4 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2518_), .B(AES_CORE_DATAPATH__abc_15863_new_n2514_), .S(AES_CORE_DATAPATH__abc_15863_new_n2463_), .Y(\iv_out[5] ));
MUX2X1 MUX2X1_40 ( .A(\bus_in[19] ), .B(AES_CORE_DATAPATH_key_host_1__19_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3963_));
MUX2X1 MUX2X1_41 ( .A(\bus_in[20] ), .B(AES_CORE_DATAPATH_key_host_1__20_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3968_));
MUX2X1 MUX2X1_42 ( .A(\bus_in[21] ), .B(AES_CORE_DATAPATH_key_host_1__21_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3973_));
MUX2X1 MUX2X1_43 ( .A(\bus_in[22] ), .B(AES_CORE_DATAPATH_key_host_1__22_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3978_));
MUX2X1 MUX2X1_44 ( .A(\bus_in[23] ), .B(AES_CORE_DATAPATH_key_host_1__23_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3983_));
MUX2X1 MUX2X1_45 ( .A(\bus_in[24] ), .B(AES_CORE_DATAPATH_key_host_1__24_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3988_));
MUX2X1 MUX2X1_46 ( .A(\bus_in[25] ), .B(AES_CORE_DATAPATH_key_host_1__25_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3993_));
MUX2X1 MUX2X1_47 ( .A(\bus_in[26] ), .B(AES_CORE_DATAPATH_key_host_1__26_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n3998_));
MUX2X1 MUX2X1_48 ( .A(\bus_in[27] ), .B(AES_CORE_DATAPATH_key_host_1__27_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4003_));
MUX2X1 MUX2X1_49 ( .A(\bus_in[28] ), .B(AES_CORE_DATAPATH_key_host_1__28_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4008_));
MUX2X1 MUX2X1_5 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2521_), .B(AES_CORE_DATAPATH__abc_15863_new_n2522_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2523_));
MUX2X1 MUX2X1_50 ( .A(\bus_in[29] ), .B(AES_CORE_DATAPATH_key_host_1__29_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4013_));
MUX2X1 MUX2X1_51 ( .A(\bus_in[30] ), .B(AES_CORE_DATAPATH_key_host_1__30_), .S(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4018_));
MUX2X1 MUX2X1_52 ( .A(\bus_in[0] ), .B(AES_CORE_DATAPATH_key_host_0__0_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4035_));
MUX2X1 MUX2X1_53 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4036_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_), .S(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4037_));
MUX2X1 MUX2X1_54 ( .A(\bus_in[1] ), .B(AES_CORE_DATAPATH_key_host_0__1_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4040_));
MUX2X1 MUX2X1_55 ( .A(\bus_in[2] ), .B(AES_CORE_DATAPATH_key_host_0__2_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4045_));
MUX2X1 MUX2X1_56 ( .A(\bus_in[3] ), .B(AES_CORE_DATAPATH_key_host_0__3_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4050_));
MUX2X1 MUX2X1_57 ( .A(\bus_in[4] ), .B(AES_CORE_DATAPATH_key_host_0__4_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4055_));
MUX2X1 MUX2X1_58 ( .A(\bus_in[5] ), .B(AES_CORE_DATAPATH_key_host_0__5_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4060_));
MUX2X1 MUX2X1_59 ( .A(\bus_in[6] ), .B(AES_CORE_DATAPATH_key_host_0__6_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4065_));
MUX2X1 MUX2X1_6 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2529_), .B(AES_CORE_DATAPATH__abc_15863_new_n2530_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2531_));
MUX2X1 MUX2X1_60 ( .A(\bus_in[7] ), .B(AES_CORE_DATAPATH_key_host_0__7_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4070_));
MUX2X1 MUX2X1_61 ( .A(\bus_in[8] ), .B(AES_CORE_DATAPATH_key_host_0__8_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4075_));
MUX2X1 MUX2X1_62 ( .A(\bus_in[9] ), .B(AES_CORE_DATAPATH_key_host_0__9_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4080_));
MUX2X1 MUX2X1_63 ( .A(\bus_in[10] ), .B(AES_CORE_DATAPATH_key_host_0__10_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4085_));
MUX2X1 MUX2X1_64 ( .A(\bus_in[11] ), .B(AES_CORE_DATAPATH_key_host_0__11_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4090_));
MUX2X1 MUX2X1_65 ( .A(\bus_in[12] ), .B(AES_CORE_DATAPATH_key_host_0__12_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4095_));
MUX2X1 MUX2X1_66 ( .A(\bus_in[13] ), .B(AES_CORE_DATAPATH_key_host_0__13_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4100_));
MUX2X1 MUX2X1_67 ( .A(\bus_in[14] ), .B(AES_CORE_DATAPATH_key_host_0__14_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4105_));
MUX2X1 MUX2X1_68 ( .A(\bus_in[15] ), .B(AES_CORE_DATAPATH_key_host_0__15_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4110_));
MUX2X1 MUX2X1_69 ( .A(\bus_in[16] ), .B(AES_CORE_DATAPATH_key_host_0__16_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4115_));
MUX2X1 MUX2X1_7 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2537_), .B(AES_CORE_DATAPATH__abc_15863_new_n2538_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2539_));
MUX2X1 MUX2X1_70 ( .A(\bus_in[17] ), .B(AES_CORE_DATAPATH_key_host_0__17_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4120_));
MUX2X1 MUX2X1_71 ( .A(\bus_in[18] ), .B(AES_CORE_DATAPATH_key_host_0__18_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4125_));
MUX2X1 MUX2X1_72 ( .A(\bus_in[19] ), .B(AES_CORE_DATAPATH_key_host_0__19_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4130_));
MUX2X1 MUX2X1_73 ( .A(\bus_in[20] ), .B(AES_CORE_DATAPATH_key_host_0__20_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4135_));
MUX2X1 MUX2X1_74 ( .A(\bus_in[21] ), .B(AES_CORE_DATAPATH_key_host_0__21_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4140_));
MUX2X1 MUX2X1_75 ( .A(\bus_in[22] ), .B(AES_CORE_DATAPATH_key_host_0__22_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4145_));
MUX2X1 MUX2X1_76 ( .A(\bus_in[23] ), .B(AES_CORE_DATAPATH_key_host_0__23_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4150_));
MUX2X1 MUX2X1_77 ( .A(\bus_in[24] ), .B(AES_CORE_DATAPATH_key_host_0__24_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4155_));
MUX2X1 MUX2X1_78 ( .A(\bus_in[25] ), .B(AES_CORE_DATAPATH_key_host_0__25_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4160_));
MUX2X1 MUX2X1_79 ( .A(\bus_in[26] ), .B(AES_CORE_DATAPATH_key_host_0__26_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4165_));
MUX2X1 MUX2X1_8 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2545_), .B(AES_CORE_DATAPATH__abc_15863_new_n2546_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2547_));
MUX2X1 MUX2X1_80 ( .A(\bus_in[27] ), .B(AES_CORE_DATAPATH_key_host_0__27_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4170_));
MUX2X1 MUX2X1_81 ( .A(\bus_in[28] ), .B(AES_CORE_DATAPATH_key_host_0__28_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4175_));
MUX2X1 MUX2X1_82 ( .A(\bus_in[29] ), .B(AES_CORE_DATAPATH_key_host_0__29_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4180_));
MUX2X1 MUX2X1_83 ( .A(\bus_in[30] ), .B(AES_CORE_DATAPATH_key_host_0__30_), .S(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4185_));
MUX2X1 MUX2X1_84 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4040_), .B(AES_CORE_DATAPATH__abc_15863_new_n2749_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__1_));
MUX2X1 MUX2X1_85 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4045_), .B(AES_CORE_DATAPATH__abc_15863_new_n2762_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__2_));
MUX2X1 MUX2X1_86 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4050_), .B(AES_CORE_DATAPATH__abc_15863_new_n2768_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__3_));
MUX2X1 MUX2X1_87 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4055_), .B(AES_CORE_DATAPATH__abc_15863_new_n2778_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__4_));
MUX2X1 MUX2X1_88 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4060_), .B(AES_CORE_DATAPATH__abc_15863_new_n2792_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__5_));
MUX2X1 MUX2X1_89 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4065_), .B(AES_CORE_DATAPATH__abc_15863_new_n2798_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__6_));
MUX2X1 MUX2X1_9 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2553_), .B(AES_CORE_DATAPATH__abc_15863_new_n2554_), .S(AES_CORE_DATAPATH__abc_15863_new_n2475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2555_));
MUX2X1 MUX2X1_90 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4070_), .B(AES_CORE_DATAPATH__abc_15863_new_n2813_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__7_));
MUX2X1 MUX2X1_91 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4075_), .B(AES_CORE_DATAPATH__abc_15863_new_n2826_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__8_));
MUX2X1 MUX2X1_92 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4080_), .B(AES_CORE_DATAPATH__abc_15863_new_n2838_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__9_));
MUX2X1 MUX2X1_93 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4085_), .B(AES_CORE_DATAPATH__abc_15863_new_n2849_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__10_));
MUX2X1 MUX2X1_94 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4090_), .B(AES_CORE_DATAPATH__abc_15863_new_n2858_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__11_));
MUX2X1 MUX2X1_95 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4095_), .B(AES_CORE_DATAPATH__abc_15863_new_n2868_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__12_));
MUX2X1 MUX2X1_96 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4100_), .B(AES_CORE_DATAPATH__abc_15863_new_n2874_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__13_));
MUX2X1 MUX2X1_97 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4105_), .B(AES_CORE_DATAPATH__abc_15863_new_n2888_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__14_));
MUX2X1 MUX2X1_98 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4110_), .B(AES_CORE_DATAPATH__abc_15863_new_n2894_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__15_));
MUX2X1 MUX2X1_99 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4115_), .B(AES_CORE_DATAPATH__abc_15863_new_n2905_), .S(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__16_));
NAND2X1 NAND2X1_1 ( .A(\addr[0] ), .B(write_en), .Y(_abc_15574_new_n13_));
NAND2X1 NAND2X1_10 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n136_));
NAND2X1 NAND2X1_100 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3038_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3039_));
NAND2X1 NAND2X1_1000 ( .A(AES_CORE_DATAPATH_bkp_1_1__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7588_));
NAND2X1 NAND2X1_1001 ( .A(AES_CORE_DATAPATH_bkp_1_1__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7593_));
NAND2X1 NAND2X1_1002 ( .A(AES_CORE_DATAPATH_bkp_1_1__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7598_));
NAND2X1 NAND2X1_1003 ( .A(AES_CORE_DATAPATH_bkp_1_1__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7603_));
NAND2X1 NAND2X1_1004 ( .A(AES_CORE_DATAPATH_bkp_1_1__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7614_));
NAND2X1 NAND2X1_1005 ( .A(AES_CORE_DATAPATH_bkp_1_1__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7619_));
NAND2X1 NAND2X1_1006 ( .A(AES_CORE_DATAPATH_bkp_1_1__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7624_));
NAND2X1 NAND2X1_1007 ( .A(AES_CORE_DATAPATH_bkp_1_1__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7632_));
NAND2X1 NAND2X1_1008 ( .A(AES_CORE_DATAPATH_bkp_1_1__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7637_));
NAND2X1 NAND2X1_1009 ( .A(AES_CORE_DATAPATH_bkp_1_1__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7639_));
NAND2X1 NAND2X1_101 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3039_), .B(AES_CORE_DATAPATH__abc_15863_new_n3037_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3040_));
NAND2X1 NAND2X1_1010 ( .A(\bus_in[6] ), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7833_));
NAND2X1 NAND2X1_1011 ( .A(\bus_in[7] ), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7836_));
NAND2X1 NAND2X1_1012 ( .A(\bus_in[8] ), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7839_));
NAND2X1 NAND2X1_1013 ( .A(\bus_in[9] ), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7842_));
NAND2X1 NAND2X1_1014 ( .A(\bus_in[10] ), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7845_));
NAND2X1 NAND2X1_1015 ( .A(\bus_in[11] ), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7848_));
NAND2X1 NAND2X1_1016 ( .A(AES_CORE_DATAPATH_bkp_1_0__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7891_));
NAND2X1 NAND2X1_1017 ( .A(AES_CORE_DATAPATH_bkp_1_0__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7893_));
NAND2X1 NAND2X1_1018 ( .A(AES_CORE_DATAPATH_bkp_1_0__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7895_));
NAND2X1 NAND2X1_1019 ( .A(AES_CORE_DATAPATH_bkp_1_0__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7897_));
NAND2X1 NAND2X1_102 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3048_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3049_));
NAND2X1 NAND2X1_1020 ( .A(AES_CORE_DATAPATH_bkp_1_0__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7899_));
NAND2X1 NAND2X1_1021 ( .A(AES_CORE_DATAPATH_bkp_1_0__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7901_));
NAND2X1 NAND2X1_1022 ( .A(AES_CORE_DATAPATH_bkp_1_0__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7903_));
NAND2X1 NAND2X1_1023 ( .A(AES_CORE_DATAPATH_bkp_1_0__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7905_));
NAND2X1 NAND2X1_1024 ( .A(AES_CORE_DATAPATH_bkp_1_0__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7907_));
NAND2X1 NAND2X1_1025 ( .A(AES_CORE_DATAPATH_bkp_1_0__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7909_));
NAND2X1 NAND2X1_1026 ( .A(AES_CORE_DATAPATH_bkp_1_0__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7911_));
NAND2X1 NAND2X1_1027 ( .A(AES_CORE_DATAPATH_bkp_1_0__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7913_));
NAND2X1 NAND2X1_1028 ( .A(AES_CORE_DATAPATH_bkp_1_0__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7915_));
NAND2X1 NAND2X1_1029 ( .A(AES_CORE_DATAPATH_bkp_1_0__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7917_));
NAND2X1 NAND2X1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3049_), .B(AES_CORE_DATAPATH__abc_15863_new_n3047_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3050_));
NAND2X1 NAND2X1_1030 ( .A(AES_CORE_DATAPATH_bkp_1_0__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7919_));
NAND2X1 NAND2X1_1031 ( .A(AES_CORE_DATAPATH_bkp_1_0__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7921_));
NAND2X1 NAND2X1_1032 ( .A(AES_CORE_DATAPATH_bkp_1_0__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7923_));
NAND2X1 NAND2X1_1033 ( .A(AES_CORE_DATAPATH_bkp_1_0__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7925_));
NAND2X1 NAND2X1_1034 ( .A(AES_CORE_DATAPATH_bkp_1_0__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7927_));
NAND2X1 NAND2X1_1035 ( .A(AES_CORE_DATAPATH_bkp_1_0__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7929_));
NAND2X1 NAND2X1_1036 ( .A(AES_CORE_DATAPATH_bkp_1_0__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7931_));
NAND2X1 NAND2X1_1037 ( .A(AES_CORE_DATAPATH_bkp_1_0__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7933_));
NAND2X1 NAND2X1_1038 ( .A(AES_CORE_DATAPATH_bkp_1_0__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7935_));
NAND2X1 NAND2X1_1039 ( .A(AES_CORE_DATAPATH_bkp_1_0__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7937_));
NAND2X1 NAND2X1_104 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3058_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3059_));
NAND2X1 NAND2X1_1040 ( .A(AES_CORE_DATAPATH_bkp_1_0__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7939_));
NAND2X1 NAND2X1_1041 ( .A(AES_CORE_DATAPATH_bkp_1_0__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7941_));
NAND2X1 NAND2X1_1042 ( .A(AES_CORE_DATAPATH_bkp_1_0__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7943_));
NAND2X1 NAND2X1_1043 ( .A(AES_CORE_DATAPATH_bkp_1_0__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7945_));
NAND2X1 NAND2X1_1044 ( .A(AES_CORE_DATAPATH_bkp_1_0__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7947_));
NAND2X1 NAND2X1_1045 ( .A(AES_CORE_DATAPATH_bkp_1_0__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7949_));
NAND2X1 NAND2X1_1046 ( .A(AES_CORE_DATAPATH_bkp_1_0__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7951_));
NAND2X1 NAND2X1_1047 ( .A(AES_CORE_DATAPATH_bkp_1_0__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7953_));
NAND2X1 NAND2X1_1048 ( .A(AES_CORE_CONTROL_UNIT_col_en_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8148_));
NAND2X1 NAND2X1_1049 ( .A(AES_CORE_CONTROL_UNIT_col_en_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8151_));
NAND2X1 NAND2X1_105 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3059_), .B(AES_CORE_DATAPATH__abc_15863_new_n3057_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3060_));
NAND2X1 NAND2X1_1050 ( .A(AES_CORE_CONTROL_UNIT_col_en_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8154_));
NAND2X1 NAND2X1_1051 ( .A(AES_CORE_CONTROL_UNIT_col_en_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8157_));
NAND2X1 NAND2X1_1052 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH_key_en_pp1_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8159_));
NAND2X1 NAND2X1_1053 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH_key_en_pp1_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8162_));
NAND2X1 NAND2X1_1054 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH_key_en_pp1_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8165_));
NAND2X1 NAND2X1_1055 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH_key_en_pp1_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8168_));
NAND2X1 NAND2X1_1056 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .B(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_DATAPATH__abc_15863_new_n8170_));
NAND2X1 NAND2X1_1057 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8172_));
NAND2X1 NAND2X1_1058 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8174_));
NAND2X1 NAND2X1_1059 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8176_));
NAND2X1 NAND2X1_106 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3063_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3064_));
NAND2X1 NAND2X1_1060 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n328_));
NAND2X1 NAND2X1_1061 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n331_));
NAND2X1 NAND2X1_1062 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n334_));
NAND2X1 NAND2X1_1063 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n337_));
NAND2X1 NAND2X1_1064 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n340_));
NAND2X1 NAND2X1_1065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n343_));
NAND2X1 NAND2X1_1066 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n346_));
NAND2X1 NAND2X1_1067 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n349_));
NAND2X1 NAND2X1_1068 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n352_));
NAND2X1 NAND2X1_1069 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n355_));
NAND2X1 NAND2X1_107 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3064_), .B(AES_CORE_DATAPATH__abc_15863_new_n3068_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3069_));
NAND2X1 NAND2X1_1070 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n358_));
NAND2X1 NAND2X1_1071 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n361_));
NAND2X1 NAND2X1_1072 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n364_));
NAND2X1 NAND2X1_1073 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n367_));
NAND2X1 NAND2X1_1074 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n370_));
NAND2X1 NAND2X1_1075 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n373_));
NAND2X1 NAND2X1_1076 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n376_));
NAND2X1 NAND2X1_1077 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n379_));
NAND2X1 NAND2X1_1078 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n382_));
NAND2X1 NAND2X1_1079 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n385_));
NAND2X1 NAND2X1_108 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_rk_sel_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3075_));
NAND2X1 NAND2X1_1080 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n388_));
NAND2X1 NAND2X1_1081 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n391_));
NAND2X1 NAND2X1_1082 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n394_));
NAND2X1 NAND2X1_1083 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n397_));
NAND2X1 NAND2X1_1084 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n400_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n401_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n402_));
NAND2X1 NAND2X1_1085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n404_));
NAND2X1 NAND2X1_1086 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n406_));
NAND2X1 NAND2X1_1087 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n408_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n409_));
NAND2X1 NAND2X1_1088 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n413_));
NAND2X1 NAND2X1_1089 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n418_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n419_));
NAND2X1 NAND2X1_109 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_rk_sel_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3078_));
NAND2X1 NAND2X1_1090 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n401_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n423_));
NAND2X1 NAND2X1_1091 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n400_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_));
NAND2X1 NAND2X1_1092 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n421_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n427_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n428_));
NAND2X1 NAND2X1_1093 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n414_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n436_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n437_));
NAND2X1 NAND2X1_1094 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_));
NAND2X1 NAND2X1_1095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n447_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n448_));
NAND2X1 NAND2X1_1096 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n443_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n448_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n449_));
NAND2X1 NAND2X1_1097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n433_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n447_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n452_));
NAND2X1 NAND2X1_1098 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n431_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n453_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n454_));
NAND2X1 NAND2X1_1099 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n450_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n454_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_));
NAND2X1 NAND2X1_11 ( .A(\aes_mode[0] ), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_));
NAND2X1 NAND2X1_110 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3086_));
NAND2X1 NAND2X1_1100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_));
NAND2X1 NAND2X1_1101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n414_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n434_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n462_));
NAND2X1 NAND2X1_1102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n466_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n467_));
NAND2X1 NAND2X1_1103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n464_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n467_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n468_));
NAND2X1 NAND2X1_1104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n458_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n466_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n471_));
NAND2X1 NAND2X1_1105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n456_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n472_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n473_));
NAND2X1 NAND2X1_1106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n469_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n473_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_));
NAND2X1 NAND2X1_1107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n479_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n480_));
NAND2X1 NAND2X1_1108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n478_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n441_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n484_));
NAND2X1 NAND2X1_1109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n481_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n485_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n486_));
NAND2X1 NAND2X1_111 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3102_), .B(AES_CORE_DATAPATH__abc_15863_new_n2740_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3103_));
NAND2X1 NAND2X1_1110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n475_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n487_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n488_));
NAND2X1 NAND2X1_1111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n488_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n491_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_));
NAND2X1 NAND2X1_1112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n499_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n500_));
NAND2X1 NAND2X1_1113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n498_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n500_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n501_));
NAND2X1 NAND2X1_1114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n495_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n499_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n504_));
NAND2X1 NAND2X1_1115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n493_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n505_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n506_));
NAND2X1 NAND2X1_1116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n502_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n506_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_));
NAND2X1 NAND2X1_1117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n509_));
NAND2X1 NAND2X1_1118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n513_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n514_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n515_));
NAND2X1 NAND2X1_1119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n522_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n523_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n524_));
NAND2X1 NAND2X1_112 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3101_), .B(AES_CORE_DATAPATH__abc_15863_new_n3097_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3104_));
NAND2X1 NAND2X1_1120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n529_));
NAND2X1 NAND2X1_1121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n533_));
NAND2X1 NAND2X1_1122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n537_));
NAND2X1 NAND2X1_1123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n541_));
NAND2X1 NAND2X1_1124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n545_));
NAND2X1 NAND2X1_1125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n549_));
NAND2X1 NAND2X1_1126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n553_));
NAND2X1 NAND2X1_1127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n557_));
NAND2X1 NAND2X1_1128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n561_));
NAND2X1 NAND2X1_1129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n565_));
NAND2X1 NAND2X1_113 ( .A(AES_CORE_DATAPATH_col_3__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3113_));
NAND2X1 NAND2X1_1130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n569_));
NAND2X1 NAND2X1_1131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n573_));
NAND2X1 NAND2X1_1132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n577_));
NAND2X1 NAND2X1_1133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n581_));
NAND2X1 NAND2X1_1134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n585_));
NAND2X1 NAND2X1_1135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n589_));
NAND2X1 NAND2X1_1136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n593_));
NAND2X1 NAND2X1_1137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n597_));
NAND2X1 NAND2X1_1138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n601_));
NAND2X1 NAND2X1_1139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n605_));
NAND2X1 NAND2X1_114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3087_), .B(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3117_));
NAND2X1 NAND2X1_1140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n609_));
NAND2X1 NAND2X1_1141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n613_));
NAND2X1 NAND2X1_1142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n617_));
NAND2X1 NAND2X1_1143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n621_));
NAND2X1 NAND2X1_1144 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n625_));
NAND2X1 NAND2X1_1145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n629_));
NAND2X1 NAND2X1_1146 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n633_));
NAND2X1 NAND2X1_1147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n637_));
NAND2X1 NAND2X1_1148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n641_));
NAND2X1 NAND2X1_1149 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n645_));
NAND2X1 NAND2X1_115 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3126_), .B(AES_CORE_DATAPATH__abc_15863_new_n2751_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3127_));
NAND2X1 NAND2X1_1150 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n649_));
NAND2X1 NAND2X1_1151 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n653_));
NAND2X1 NAND2X1_1152 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n420_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n428_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n680_));
NAND2X1 NAND2X1_1153 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n683_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n449_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n684_));
NAND2X1 NAND2X1_1154 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n682_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n684_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_));
NAND2X1 NAND2X1_1155 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n689_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n501_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n690_));
NAND2X1 NAND2X1_1156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n688_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n690_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_));
NAND2X1 NAND2X1_1157 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n512_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n515_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n692_));
NAND2X1 NAND2X1_1158 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n521_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n524_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n694_));
NAND2X1 NAND2X1_1159 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n102_));
NAND2X1 NAND2X1_116 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3125_), .B(AES_CORE_DATAPATH__abc_15863_new_n3124_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3128_));
NAND2X1 NAND2X1_1160 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n102_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n101_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_));
NAND2X1 NAND2X1_1161 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n104_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n105_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n106_));
NAND2X1 NAND2X1_1162 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n113_));
NAND2X1 NAND2X1_1163 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n106_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n111_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_));
NAND2X1 NAND2X1_1164 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n119_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n113_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n120_));
NAND2X1 NAND2X1_1165 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n128_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n129_));
NAND2X1 NAND2X1_1166 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n130_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n131_));
NAND2X1 NAND2X1_1167 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n116_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n133_));
NAND2X1 NAND2X1_1168 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n114_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n134_));
NAND2X1 NAND2X1_1169 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n136_));
NAND2X1 NAND2X1_117 ( .A(AES_CORE_DATAPATH_col_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3136_));
NAND2X1 NAND2X1_1170 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n142_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n143_));
NAND2X1 NAND2X1_1171 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n133_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n134_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n144_));
NAND2X1 NAND2X1_1172 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n145_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n146_));
NAND2X1 NAND2X1_1173 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n154_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n157_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_));
NAND2X1 NAND2X1_1174 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n136_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n135_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n163_));
NAND2X1 NAND2X1_1175 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n129_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n131_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n166_));
NAND2X1 NAND2X1_1176 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n171_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n172_));
NAND2X1 NAND2X1_1177 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n173_));
NAND2X1 NAND2X1_1178 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n173_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n172_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n174_));
NAND2X1 NAND2X1_1179 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n177_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n178_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n179_));
NAND2X1 NAND2X1_118 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3139_));
NAND2X1 NAND2X1_1180 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n180_));
NAND2X1 NAND2X1_1181 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n180_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n179_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_));
NAND2X1 NAND2X1_1182 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n187_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n193_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n194_));
NAND2X1 NAND2X1_1183 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n214_));
NAND2X1 NAND2X1_1184 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n216_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n221_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n222_));
NAND2X1 NAND2X1_1185 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n228_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n231_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_));
NAND2X1 NAND2X1_1186 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n239_));
NAND2X1 NAND2X1_1187 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n239_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n238_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n240_));
NAND2X1 NAND2X1_1188 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n241_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n243_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n244_));
NAND2X1 NAND2X1_1189 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n255_));
NAND2X1 NAND2X1_119 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3148_), .B(AES_CORE_DATAPATH__abc_15863_new_n2764_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3149_));
NAND2X1 NAND2X1_1190 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n257_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n253_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n259_));
NAND2X1 NAND2X1_1191 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n217_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n219_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n262_));
NAND2X1 NAND2X1_1192 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n214_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n262_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n264_));
NAND2X1 NAND2X1_1193 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n249_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n267_));
NAND2X1 NAND2X1_1194 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n247_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n268_));
NAND2X1 NAND2X1_1195 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n171_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n269_));
NAND2X1 NAND2X1_1196 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n270_));
NAND2X1 NAND2X1_1197 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n247_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n249_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n272_));
NAND2X1 NAND2X1_1198 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n274_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n222_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n275_));
NAND2X1 NAND2X1_1199 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n278_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n279_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n280_));
NAND2X1 NAND2X1_12 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n154_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n157_));
NAND2X1 NAND2X1_120 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3147_), .B(AES_CORE_DATAPATH__abc_15863_new_n3146_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3150_));
NAND2X1 NAND2X1_1200 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n284_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n288_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_));
NAND2X1 NAND2X1_1201 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n294_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n166_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n295_));
NAND2X1 NAND2X1_1202 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n163_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n296_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n297_));
NAND2X1 NAND2X1_1203 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n295_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n297_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n298_));
NAND2X1 NAND2X1_1204 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n166_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n296_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n311_));
NAND2X1 NAND2X1_1205 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n163_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n294_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n312_));
NAND2X1 NAND2X1_1206 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n312_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n311_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n313_));
NAND2X1 NAND2X1_1207 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n317_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n320_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_));
NAND2X1 NAND2X1_1208 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n328_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n298_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n329_));
NAND2X1 NAND2X1_1209 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n330_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n313_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n331_));
NAND2X1 NAND2X1_121 ( .A(AES_CORE_DATAPATH_col_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3158_));
NAND2X1 NAND2X1_1210 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n328_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n313_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n334_));
NAND2X1 NAND2X1_1211 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n330_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n298_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n335_));
NAND2X1 NAND2X1_1212 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n340_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n337_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_));
NAND2X1 NAND2X1_1213 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n345_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n346_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n347_));
NAND2X1 NAND2X1_1214 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n348_));
NAND2X1 NAND2X1_1215 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n348_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n347_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n349_));
NAND2X1 NAND2X1_1216 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n367_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n369_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_));
NAND2X1 NAND2X1_1217 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n375_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n377_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n378_));
NAND2X1 NAND2X1_1218 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n391_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n388_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_));
NAND2X1 NAND2X1_1219 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n300_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n301_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n398_));
NAND2X1 NAND2X1_122 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3170_), .B(AES_CORE_DATAPATH__abc_15863_new_n3169_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3173_));
NAND2X1 NAND2X1_1220 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n402_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n405_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_));
NAND2X1 NAND2X1_1221 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n414_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n417_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_));
NAND2X1 NAND2X1_1222 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n446_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n447_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_));
NAND2X1 NAND2X1_1223 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n457_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n458_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_));
NAND2X1 NAND2X1_1224 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n464_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n466_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_));
NAND2X1 NAND2X1_1225 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n471_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n472_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_));
NAND2X1 NAND2X1_1226 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n478_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n479_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_));
NAND2X1 NAND2X1_1227 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n493_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n494_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_));
NAND2X1 NAND2X1_1228 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n504_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n505_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_));
NAND2X1 NAND2X1_1229 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n511_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n512_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_));
NAND2X1 NAND2X1_123 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3173_), .B(AES_CORE_DATAPATH__abc_15863_new_n2774_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3174_));
NAND2X1 NAND2X1_1230 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n518_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n519_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_));
NAND2X1 NAND2X1_1231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n52_));
NAND2X1 NAND2X1_1232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n51_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_));
NAND2X1 NAND2X1_1233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n58_));
NAND2X1 NAND2X1_1234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n60_));
NAND2X1 NAND2X1_1235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n63_));
NAND2X1 NAND2X1_1236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n64_));
NAND2X1 NAND2X1_1237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n70_));
NAND2X1 NAND2X1_1238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n71_));
NAND2X1 NAND2X1_1239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n72_));
NAND2X1 NAND2X1_124 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3179_), .B(AES_CORE_DATAPATH__abc_15863_new_n3175_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3180_));
NAND2X1 NAND2X1_1240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n73_));
NAND2X1 NAND2X1_1241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n74_));
NAND2X1 NAND2X1_1242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n75_));
NAND2X1 NAND2X1_1243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n74_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n76_));
NAND2X1 NAND2X1_1244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n76_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n77_));
NAND2X1 NAND2X1_1245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n64_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n84_));
NAND2X1 NAND2X1_1246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n85_));
NAND2X1 NAND2X1_1247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n87_));
NAND2X1 NAND2X1_1248 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n88_));
NAND2X1 NAND2X1_1249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n97_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n98_));
NAND2X1 NAND2X1_125 ( .A(AES_CORE_DATAPATH_col_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3181_));
NAND2X1 NAND2X1_1250 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n101_));
NAND2X1 NAND2X1_1251 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n98_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n101_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n102_));
NAND2X1 NAND2X1_1252 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n104_));
NAND2X1 NAND2X1_1253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n104_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n103_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n105_));
NAND2X1 NAND2X1_1254 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n110_));
NAND2X1 NAND2X1_1255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n111_));
NAND2X1 NAND2X1_1256 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_));
NAND2X1 NAND2X1_1257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n125_));
NAND2X1 NAND2X1_1258 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n130_));
NAND2X1 NAND2X1_1259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n132_));
NAND2X1 NAND2X1_126 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3184_));
NAND2X1 NAND2X1_1260 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n139_));
NAND2X1 NAND2X1_1261 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n144_));
NAND2X1 NAND2X1_1262 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n151_));
NAND2X1 NAND2X1_1263 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n154_));
NAND2X1 NAND2X1_1264 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n155_));
NAND2X1 NAND2X1_1265 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n155_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n156_));
NAND2X1 NAND2X1_1266 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n160_));
NAND2X1 NAND2X1_1267 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n161_));
NAND2X1 NAND2X1_1268 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n162_));
NAND2X1 NAND2X1_1269 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n163_));
NAND2X1 NAND2X1_127 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3193_), .B(AES_CORE_DATAPATH__abc_15863_new_n2784_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3194_));
NAND2X1 NAND2X1_1270 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n164_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n165_));
NAND2X1 NAND2X1_1271 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n168_));
NAND2X1 NAND2X1_1272 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_));
NAND2X1 NAND2X1_1273 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n174_));
NAND2X1 NAND2X1_1274 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n179_));
NAND2X1 NAND2X1_1275 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n180_));
NAND2X1 NAND2X1_1276 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_));
NAND2X1 NAND2X1_1277 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n179_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n189_));
NAND2X1 NAND2X1_1278 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n191_));
NAND2X1 NAND2X1_1279 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n192_));
NAND2X1 NAND2X1_128 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3192_), .B(AES_CORE_DATAPATH__abc_15863_new_n3191_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3195_));
NAND2X1 NAND2X1_1280 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n191_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n193_));
NAND2X1 NAND2X1_1281 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n190_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n194_));
NAND2X1 NAND2X1_1282 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n197_));
NAND2X1 NAND2X1_1283 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n201_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n202_));
NAND2X1 NAND2X1_1284 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n202_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_));
NAND2X1 NAND2X1_1285 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n207_));
NAND2X1 NAND2X1_1286 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n212_));
NAND2X1 NAND2X1_1287 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n215_));
NAND2X1 NAND2X1_1288 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n217_));
NAND2X1 NAND2X1_1289 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n215_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n217_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n218_));
NAND2X1 NAND2X1_129 ( .A(AES_CORE_DATAPATH_col_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3203_));
NAND2X1 NAND2X1_1290 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n222_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_));
NAND2X1 NAND2X1_1291 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n228_));
NAND2X1 NAND2X1_1292 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n229_));
NAND2X1 NAND2X1_1293 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n229_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n228_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n230_));
NAND2X1 NAND2X1_1294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n233_));
NAND2X1 NAND2X1_1295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n233_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n234_));
NAND2X1 NAND2X1_1296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n237_));
NAND2X1 NAND2X1_1297 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n239_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n241_));
NAND2X1 NAND2X1_1298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n237_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n241_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n242_));
NAND2X1 NAND2X1_1299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n243_));
NAND2X1 NAND2X1_13 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n163_));
NAND2X1 NAND2X1_130 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3206_));
NAND2X1 NAND2X1_1300 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n244_));
NAND2X1 NAND2X1_1301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n245_));
NAND2X1 NAND2X1_1302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n246_));
NAND2X1 NAND2X1_1303 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n247_));
NAND2X1 NAND2X1_1304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n248_));
NAND2X1 NAND2X1_1305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n249_));
NAND2X1 NAND2X1_1306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n251_));
NAND2X1 NAND2X1_1307 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n252_));
NAND2X1 NAND2X1_1308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n254_));
NAND2X1 NAND2X1_1309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n258_));
NAND2X1 NAND2X1_131 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3215_), .B(AES_CORE_DATAPATH__abc_15863_new_n2794_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3216_));
NAND2X1 NAND2X1_1310 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n259_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n262_));
NAND2X1 NAND2X1_1311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n253_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n264_));
NAND2X1 NAND2X1_1312 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n257_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n265_));
NAND2X1 NAND2X1_1313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n263_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n268_));
NAND2X1 NAND2X1_1314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n274_));
NAND2X1 NAND2X1_1315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n275_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n269_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_));
NAND2X1 NAND2X1_1316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n258_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n277_));
NAND2X1 NAND2X1_1317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n280_));
NAND2X1 NAND2X1_1318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n281_));
NAND2X1 NAND2X1_1319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n284_));
NAND2X1 NAND2X1_132 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3214_), .B(AES_CORE_DATAPATH__abc_15863_new_n3213_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3217_));
NAND2X1 NAND2X1_1320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n287_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n288_));
NAND2X1 NAND2X1_1321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n295_));
NAND2X1 NAND2X1_1322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n303_));
NAND2X1 NAND2X1_1323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_));
NAND2X1 NAND2X1_1324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n315_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n317_));
NAND2X1 NAND2X1_1325 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n320_));
NAND2X1 NAND2X1_1326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n323_));
NAND2X1 NAND2X1_1327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n321_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n324_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_));
NAND2X1 NAND2X1_1328 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n328_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n329_));
NAND2X1 NAND2X1_1329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n334_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_));
NAND2X1 NAND2X1_133 ( .A(AES_CORE_DATAPATH_col_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3225_));
NAND2X1 NAND2X1_1330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n340_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_));
NAND2X1 NAND2X1_1331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n348_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_));
NAND2X1 NAND2X1_1332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_));
NAND2X1 NAND2X1_1333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_));
NAND2X1 NAND2X1_1334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n370_));
NAND2X1 NAND2X1_1335 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n374_));
NAND2X1 NAND2X1_1336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n375_));
NAND2X1 NAND2X1_1337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n376_));
NAND2X1 NAND2X1_1338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n376_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n382_));
NAND2X1 NAND2X1_1339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n383_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_));
NAND2X1 NAND2X1_134 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3228_));
NAND2X1 NAND2X1_1340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n393_));
NAND2X1 NAND2X1_1341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n405_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n404_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n406_));
NAND2X1 NAND2X1_1342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n408_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n410_));
NAND2X1 NAND2X1_1343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_));
NAND2X1 NAND2X1_1344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n421_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n417_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_));
NAND2X1 NAND2X1_1345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n397_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n396_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n427_));
NAND2X1 NAND2X1_1346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n429_));
NAND2X1 NAND2X1_1347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n435_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n436_));
NAND2X1 NAND2X1_1348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n442_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n444_));
NAND2X1 NAND2X1_1349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n438_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n450_));
NAND2X1 NAND2X1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3237_), .B(AES_CORE_DATAPATH__abc_15863_new_n2804_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3238_));
NAND2X1 NAND2X1_1350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_));
NAND2X1 NAND2X1_1351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n456_));
NAND2X1 NAND2X1_1352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n434_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n466_));
NAND2X1 NAND2X1_1353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n467_));
NAND2X1 NAND2X1_1354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n463_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n469_));
NAND2X1 NAND2X1_1355 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n471_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_));
NAND2X1 NAND2X1_1356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n489_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n486_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_));
NAND2X1 NAND2X1_1357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_));
NAND2X1 NAND2X1_1358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n377_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_));
NAND2X1 NAND2X1_1359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n52_));
NAND2X1 NAND2X1_136 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3236_), .B(AES_CORE_DATAPATH__abc_15863_new_n3235_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3239_));
NAND2X1 NAND2X1_1360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n51_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_));
NAND2X1 NAND2X1_1361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n58_));
NAND2X1 NAND2X1_1362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n60_));
NAND2X1 NAND2X1_1363 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n63_));
NAND2X1 NAND2X1_1364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n64_));
NAND2X1 NAND2X1_1365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n70_));
NAND2X1 NAND2X1_1366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n71_));
NAND2X1 NAND2X1_1367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n72_));
NAND2X1 NAND2X1_1368 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n73_));
NAND2X1 NAND2X1_1369 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n74_));
NAND2X1 NAND2X1_137 ( .A(AES_CORE_DATAPATH_col_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3247_));
NAND2X1 NAND2X1_1370 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n75_));
NAND2X1 NAND2X1_1371 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n74_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n76_));
NAND2X1 NAND2X1_1372 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n76_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n77_));
NAND2X1 NAND2X1_1373 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n64_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n84_));
NAND2X1 NAND2X1_1374 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n85_));
NAND2X1 NAND2X1_1375 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n87_));
NAND2X1 NAND2X1_1376 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n88_));
NAND2X1 NAND2X1_1377 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n97_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n98_));
NAND2X1 NAND2X1_1378 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n101_));
NAND2X1 NAND2X1_1379 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n98_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n101_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n102_));
NAND2X1 NAND2X1_138 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3259_), .B(AES_CORE_DATAPATH__abc_15863_new_n2815_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3260_));
NAND2X1 NAND2X1_1380 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n104_));
NAND2X1 NAND2X1_1381 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n104_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n103_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n105_));
NAND2X1 NAND2X1_1382 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n110_));
NAND2X1 NAND2X1_1383 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n111_));
NAND2X1 NAND2X1_1384 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_));
NAND2X1 NAND2X1_1385 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n125_));
NAND2X1 NAND2X1_1386 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n130_));
NAND2X1 NAND2X1_1387 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n132_));
NAND2X1 NAND2X1_1388 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n139_));
NAND2X1 NAND2X1_1389 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n144_));
NAND2X1 NAND2X1_139 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3258_), .B(AES_CORE_DATAPATH__abc_15863_new_n3257_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3261_));
NAND2X1 NAND2X1_1390 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n151_));
NAND2X1 NAND2X1_1391 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n154_));
NAND2X1 NAND2X1_1392 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n155_));
NAND2X1 NAND2X1_1393 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n155_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n156_));
NAND2X1 NAND2X1_1394 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n160_));
NAND2X1 NAND2X1_1395 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n161_));
NAND2X1 NAND2X1_1396 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n162_));
NAND2X1 NAND2X1_1397 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n163_));
NAND2X1 NAND2X1_1398 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n164_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n165_));
NAND2X1 NAND2X1_1399 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n168_));
NAND2X1 NAND2X1_14 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n168_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n169_));
NAND2X1 NAND2X1_140 ( .A(AES_CORE_DATAPATH_col_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3269_));
NAND2X1 NAND2X1_1400 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_));
NAND2X1 NAND2X1_1401 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n174_));
NAND2X1 NAND2X1_1402 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n179_));
NAND2X1 NAND2X1_1403 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n180_));
NAND2X1 NAND2X1_1404 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_));
NAND2X1 NAND2X1_1405 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n179_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n189_));
NAND2X1 NAND2X1_1406 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n191_));
NAND2X1 NAND2X1_1407 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n192_));
NAND2X1 NAND2X1_1408 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n191_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n193_));
NAND2X1 NAND2X1_1409 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n190_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n194_));
NAND2X1 NAND2X1_141 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3272_));
NAND2X1 NAND2X1_1410 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n197_));
NAND2X1 NAND2X1_1411 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n201_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n202_));
NAND2X1 NAND2X1_1412 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n202_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_));
NAND2X1 NAND2X1_1413 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n207_));
NAND2X1 NAND2X1_1414 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n212_));
NAND2X1 NAND2X1_1415 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n215_));
NAND2X1 NAND2X1_1416 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n217_));
NAND2X1 NAND2X1_1417 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n215_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n217_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n218_));
NAND2X1 NAND2X1_1418 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n222_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_));
NAND2X1 NAND2X1_1419 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n228_));
NAND2X1 NAND2X1_142 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3281_), .B(AES_CORE_DATAPATH__abc_15863_new_n2828_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3282_));
NAND2X1 NAND2X1_1420 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n229_));
NAND2X1 NAND2X1_1421 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n229_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n228_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n230_));
NAND2X1 NAND2X1_1422 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n233_));
NAND2X1 NAND2X1_1423 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n233_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n234_));
NAND2X1 NAND2X1_1424 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n237_));
NAND2X1 NAND2X1_1425 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n239_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n241_));
NAND2X1 NAND2X1_1426 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n237_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n241_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n242_));
NAND2X1 NAND2X1_1427 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n243_));
NAND2X1 NAND2X1_1428 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n244_));
NAND2X1 NAND2X1_1429 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n245_));
NAND2X1 NAND2X1_143 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3280_), .B(AES_CORE_DATAPATH__abc_15863_new_n3279_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3283_));
NAND2X1 NAND2X1_1430 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n246_));
NAND2X1 NAND2X1_1431 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n247_));
NAND2X1 NAND2X1_1432 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n248_));
NAND2X1 NAND2X1_1433 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n249_));
NAND2X1 NAND2X1_1434 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n251_));
NAND2X1 NAND2X1_1435 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n252_));
NAND2X1 NAND2X1_1436 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n254_));
NAND2X1 NAND2X1_1437 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n258_));
NAND2X1 NAND2X1_1438 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n259_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n262_));
NAND2X1 NAND2X1_1439 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n253_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n264_));
NAND2X1 NAND2X1_144 ( .A(AES_CORE_DATAPATH_col_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3291_));
NAND2X1 NAND2X1_1440 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n257_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n265_));
NAND2X1 NAND2X1_1441 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n263_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n268_));
NAND2X1 NAND2X1_1442 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n274_));
NAND2X1 NAND2X1_1443 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n275_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n269_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_));
NAND2X1 NAND2X1_1444 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n258_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n277_));
NAND2X1 NAND2X1_1445 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n280_));
NAND2X1 NAND2X1_1446 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n281_));
NAND2X1 NAND2X1_1447 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n284_));
NAND2X1 NAND2X1_1448 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n287_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n288_));
NAND2X1 NAND2X1_1449 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n295_));
NAND2X1 NAND2X1_145 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3302_), .B(AES_CORE_DATAPATH__abc_15863_new_n3301_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3305_));
NAND2X1 NAND2X1_1450 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n303_));
NAND2X1 NAND2X1_1451 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_));
NAND2X1 NAND2X1_1452 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n315_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n317_));
NAND2X1 NAND2X1_1453 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n320_));
NAND2X1 NAND2X1_1454 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n323_));
NAND2X1 NAND2X1_1455 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n321_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n324_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_));
NAND2X1 NAND2X1_1456 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n328_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n329_));
NAND2X1 NAND2X1_1457 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n334_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_));
NAND2X1 NAND2X1_1458 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n340_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_));
NAND2X1 NAND2X1_1459 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n348_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_));
NAND2X1 NAND2X1_146 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3305_), .B(AES_CORE_DATAPATH__abc_15863_new_n2840_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3306_));
NAND2X1 NAND2X1_1460 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_));
NAND2X1 NAND2X1_1461 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_));
NAND2X1 NAND2X1_1462 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n370_));
NAND2X1 NAND2X1_1463 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n374_));
NAND2X1 NAND2X1_1464 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n375_));
NAND2X1 NAND2X1_1465 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n376_));
NAND2X1 NAND2X1_1466 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n376_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n382_));
NAND2X1 NAND2X1_1467 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n383_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_));
NAND2X1 NAND2X1_1468 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n393_));
NAND2X1 NAND2X1_1469 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n405_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n404_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n406_));
NAND2X1 NAND2X1_147 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3311_), .B(AES_CORE_DATAPATH__abc_15863_new_n3307_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3312_));
NAND2X1 NAND2X1_1470 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n408_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n410_));
NAND2X1 NAND2X1_1471 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_));
NAND2X1 NAND2X1_1472 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n421_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n417_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_));
NAND2X1 NAND2X1_1473 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n397_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n396_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n427_));
NAND2X1 NAND2X1_1474 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n429_));
NAND2X1 NAND2X1_1475 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n435_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n436_));
NAND2X1 NAND2X1_1476 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n442_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n444_));
NAND2X1 NAND2X1_1477 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n438_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n450_));
NAND2X1 NAND2X1_1478 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_));
NAND2X1 NAND2X1_1479 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n456_));
NAND2X1 NAND2X1_148 ( .A(AES_CORE_DATAPATH_col_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3313_));
NAND2X1 NAND2X1_1480 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n434_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n466_));
NAND2X1 NAND2X1_1481 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n467_));
NAND2X1 NAND2X1_1482 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n463_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n469_));
NAND2X1 NAND2X1_1483 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n471_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_));
NAND2X1 NAND2X1_1484 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n489_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n486_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_));
NAND2X1 NAND2X1_1485 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_));
NAND2X1 NAND2X1_1486 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n377_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_));
NAND2X1 NAND2X1_1487 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n52_));
NAND2X1 NAND2X1_1488 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n51_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_));
NAND2X1 NAND2X1_1489 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n58_));
NAND2X1 NAND2X1_149 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3316_));
NAND2X1 NAND2X1_1490 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n60_));
NAND2X1 NAND2X1_1491 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n63_));
NAND2X1 NAND2X1_1492 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n64_));
NAND2X1 NAND2X1_1493 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n70_));
NAND2X1 NAND2X1_1494 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n71_));
NAND2X1 NAND2X1_1495 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n72_));
NAND2X1 NAND2X1_1496 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n73_));
NAND2X1 NAND2X1_1497 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n74_));
NAND2X1 NAND2X1_1498 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n75_));
NAND2X1 NAND2X1_1499 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n74_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n76_));
NAND2X1 NAND2X1_15 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n188_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n186_), .Y(AES_CORE_CONTROL_UNIT_col_sel_0_));
NAND2X1 NAND2X1_150 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3325_), .B(AES_CORE_DATAPATH__abc_15863_new_n2851_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3326_));
NAND2X1 NAND2X1_1500 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n76_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n77_));
NAND2X1 NAND2X1_1501 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n64_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n84_));
NAND2X1 NAND2X1_1502 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n85_));
NAND2X1 NAND2X1_1503 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n87_));
NAND2X1 NAND2X1_1504 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n88_));
NAND2X1 NAND2X1_1505 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n97_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n98_));
NAND2X1 NAND2X1_1506 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n101_));
NAND2X1 NAND2X1_1507 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n98_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n101_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n102_));
NAND2X1 NAND2X1_1508 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n104_));
NAND2X1 NAND2X1_1509 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n104_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n103_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n105_));
NAND2X1 NAND2X1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3324_), .B(AES_CORE_DATAPATH__abc_15863_new_n3323_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3327_));
NAND2X1 NAND2X1_1510 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n110_));
NAND2X1 NAND2X1_1511 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n111_));
NAND2X1 NAND2X1_1512 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_));
NAND2X1 NAND2X1_1513 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n125_));
NAND2X1 NAND2X1_1514 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n130_));
NAND2X1 NAND2X1_1515 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n132_));
NAND2X1 NAND2X1_1516 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n139_));
NAND2X1 NAND2X1_1517 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n144_));
NAND2X1 NAND2X1_1518 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n151_));
NAND2X1 NAND2X1_1519 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n154_));
NAND2X1 NAND2X1_152 ( .A(AES_CORE_DATAPATH_col_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3335_));
NAND2X1 NAND2X1_1520 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n155_));
NAND2X1 NAND2X1_1521 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n155_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n156_));
NAND2X1 NAND2X1_1522 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n160_));
NAND2X1 NAND2X1_1523 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n161_));
NAND2X1 NAND2X1_1524 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n162_));
NAND2X1 NAND2X1_1525 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n163_));
NAND2X1 NAND2X1_1526 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n164_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n165_));
NAND2X1 NAND2X1_1527 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n168_));
NAND2X1 NAND2X1_1528 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_));
NAND2X1 NAND2X1_1529 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n174_));
NAND2X1 NAND2X1_153 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3346_), .B(AES_CORE_DATAPATH__abc_15863_new_n3345_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3349_));
NAND2X1 NAND2X1_1530 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n179_));
NAND2X1 NAND2X1_1531 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n180_));
NAND2X1 NAND2X1_1532 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_));
NAND2X1 NAND2X1_1533 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n179_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n189_));
NAND2X1 NAND2X1_1534 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n191_));
NAND2X1 NAND2X1_1535 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n192_));
NAND2X1 NAND2X1_1536 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n191_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n193_));
NAND2X1 NAND2X1_1537 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n190_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n194_));
NAND2X1 NAND2X1_1538 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n197_));
NAND2X1 NAND2X1_1539 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n201_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n202_));
NAND2X1 NAND2X1_154 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3349_), .B(AES_CORE_DATAPATH__abc_15863_new_n2860_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3350_));
NAND2X1 NAND2X1_1540 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n202_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_));
NAND2X1 NAND2X1_1541 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n207_));
NAND2X1 NAND2X1_1542 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n212_));
NAND2X1 NAND2X1_1543 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n215_));
NAND2X1 NAND2X1_1544 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n217_));
NAND2X1 NAND2X1_1545 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n215_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n217_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n218_));
NAND2X1 NAND2X1_1546 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n222_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_));
NAND2X1 NAND2X1_1547 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n228_));
NAND2X1 NAND2X1_1548 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n229_));
NAND2X1 NAND2X1_1549 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n229_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n228_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n230_));
NAND2X1 NAND2X1_155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3355_), .B(AES_CORE_DATAPATH__abc_15863_new_n3351_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3356_));
NAND2X1 NAND2X1_1550 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n233_));
NAND2X1 NAND2X1_1551 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n233_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n234_));
NAND2X1 NAND2X1_1552 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n237_));
NAND2X1 NAND2X1_1553 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n239_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n241_));
NAND2X1 NAND2X1_1554 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n237_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n241_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n242_));
NAND2X1 NAND2X1_1555 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n243_));
NAND2X1 NAND2X1_1556 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n244_));
NAND2X1 NAND2X1_1557 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n245_));
NAND2X1 NAND2X1_1558 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n246_));
NAND2X1 NAND2X1_1559 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n247_));
NAND2X1 NAND2X1_156 ( .A(AES_CORE_DATAPATH_col_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3357_));
NAND2X1 NAND2X1_1560 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n248_));
NAND2X1 NAND2X1_1561 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n249_));
NAND2X1 NAND2X1_1562 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n251_));
NAND2X1 NAND2X1_1563 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n252_));
NAND2X1 NAND2X1_1564 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n254_));
NAND2X1 NAND2X1_1565 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n258_));
NAND2X1 NAND2X1_1566 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n259_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n262_));
NAND2X1 NAND2X1_1567 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n253_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n264_));
NAND2X1 NAND2X1_1568 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n257_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n265_));
NAND2X1 NAND2X1_1569 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n263_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n268_));
NAND2X1 NAND2X1_157 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3360_));
NAND2X1 NAND2X1_1570 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n274_));
NAND2X1 NAND2X1_1571 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n275_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n269_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_));
NAND2X1 NAND2X1_1572 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n258_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n277_));
NAND2X1 NAND2X1_1573 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n280_));
NAND2X1 NAND2X1_1574 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n281_));
NAND2X1 NAND2X1_1575 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n284_));
NAND2X1 NAND2X1_1576 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n287_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n288_));
NAND2X1 NAND2X1_1577 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n295_));
NAND2X1 NAND2X1_1578 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n303_));
NAND2X1 NAND2X1_1579 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_));
NAND2X1 NAND2X1_158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3369_), .B(AES_CORE_DATAPATH__abc_15863_new_n2870_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3370_));
NAND2X1 NAND2X1_1580 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n315_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n317_));
NAND2X1 NAND2X1_1581 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n320_));
NAND2X1 NAND2X1_1582 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n323_));
NAND2X1 NAND2X1_1583 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n321_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n324_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_));
NAND2X1 NAND2X1_1584 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n328_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n329_));
NAND2X1 NAND2X1_1585 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n334_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_));
NAND2X1 NAND2X1_1586 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n340_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_));
NAND2X1 NAND2X1_1587 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n348_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_));
NAND2X1 NAND2X1_1588 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_));
NAND2X1 NAND2X1_1589 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_));
NAND2X1 NAND2X1_159 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3368_), .B(AES_CORE_DATAPATH__abc_15863_new_n3367_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3371_));
NAND2X1 NAND2X1_1590 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n370_));
NAND2X1 NAND2X1_1591 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n374_));
NAND2X1 NAND2X1_1592 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n375_));
NAND2X1 NAND2X1_1593 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n376_));
NAND2X1 NAND2X1_1594 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n376_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n382_));
NAND2X1 NAND2X1_1595 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n383_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_));
NAND2X1 NAND2X1_1596 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n393_));
NAND2X1 NAND2X1_1597 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n405_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n404_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n406_));
NAND2X1 NAND2X1_1598 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n408_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n410_));
NAND2X1 NAND2X1_1599 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_));
NAND2X1 NAND2X1_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT_key_out_sel_0_));
NAND2X1 NAND2X1_160 ( .A(AES_CORE_DATAPATH_col_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3379_));
NAND2X1 NAND2X1_1600 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n421_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n417_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_));
NAND2X1 NAND2X1_1601 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n397_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n396_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n427_));
NAND2X1 NAND2X1_1602 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n429_));
NAND2X1 NAND2X1_1603 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n435_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n436_));
NAND2X1 NAND2X1_1604 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n442_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n444_));
NAND2X1 NAND2X1_1605 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n438_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n450_));
NAND2X1 NAND2X1_1606 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_));
NAND2X1 NAND2X1_1607 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n456_));
NAND2X1 NAND2X1_1608 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n434_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n466_));
NAND2X1 NAND2X1_1609 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n467_));
NAND2X1 NAND2X1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3390_), .B(AES_CORE_DATAPATH__abc_15863_new_n3389_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3393_));
NAND2X1 NAND2X1_1610 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n463_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n469_));
NAND2X1 NAND2X1_1611 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n471_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_));
NAND2X1 NAND2X1_1612 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n489_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n486_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_));
NAND2X1 NAND2X1_1613 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_));
NAND2X1 NAND2X1_1614 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n377_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_));
NAND2X1 NAND2X1_1615 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n52_));
NAND2X1 NAND2X1_1616 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n51_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_));
NAND2X1 NAND2X1_1617 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n58_));
NAND2X1 NAND2X1_1618 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n60_));
NAND2X1 NAND2X1_1619 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n63_));
NAND2X1 NAND2X1_162 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3393_), .B(AES_CORE_DATAPATH__abc_15863_new_n2880_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3394_));
NAND2X1 NAND2X1_1620 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n64_));
NAND2X1 NAND2X1_1621 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n70_));
NAND2X1 NAND2X1_1622 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n71_));
NAND2X1 NAND2X1_1623 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n72_));
NAND2X1 NAND2X1_1624 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n73_));
NAND2X1 NAND2X1_1625 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n74_));
NAND2X1 NAND2X1_1626 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n75_));
NAND2X1 NAND2X1_1627 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n74_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n76_));
NAND2X1 NAND2X1_1628 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n76_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n77_));
NAND2X1 NAND2X1_1629 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n64_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n84_));
NAND2X1 NAND2X1_163 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3399_), .B(AES_CORE_DATAPATH__abc_15863_new_n3395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3400_));
NAND2X1 NAND2X1_1630 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n85_));
NAND2X1 NAND2X1_1631 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n87_));
NAND2X1 NAND2X1_1632 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n88_));
NAND2X1 NAND2X1_1633 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n97_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n98_));
NAND2X1 NAND2X1_1634 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n101_));
NAND2X1 NAND2X1_1635 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n98_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n101_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n102_));
NAND2X1 NAND2X1_1636 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n104_));
NAND2X1 NAND2X1_1637 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n104_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n103_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n105_));
NAND2X1 NAND2X1_1638 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n110_));
NAND2X1 NAND2X1_1639 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n69_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n87_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n111_));
NAND2X1 NAND2X1_164 ( .A(AES_CORE_DATAPATH_col_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3401_));
NAND2X1 NAND2X1_1640 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_));
NAND2X1 NAND2X1_1641 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n125_));
NAND2X1 NAND2X1_1642 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n130_));
NAND2X1 NAND2X1_1643 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n132_));
NAND2X1 NAND2X1_1644 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n139_));
NAND2X1 NAND2X1_1645 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n144_));
NAND2X1 NAND2X1_1646 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n151_));
NAND2X1 NAND2X1_1647 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n154_));
NAND2X1 NAND2X1_1648 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n155_));
NAND2X1 NAND2X1_1649 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n155_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n156_));
NAND2X1 NAND2X1_165 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3404_));
NAND2X1 NAND2X1_1650 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n160_));
NAND2X1 NAND2X1_1651 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n161_));
NAND2X1 NAND2X1_1652 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n162_));
NAND2X1 NAND2X1_1653 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n163_));
NAND2X1 NAND2X1_1654 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n164_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n165_));
NAND2X1 NAND2X1_1655 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n166_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n168_));
NAND2X1 NAND2X1_1656 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_));
NAND2X1 NAND2X1_1657 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n174_));
NAND2X1 NAND2X1_1658 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n179_));
NAND2X1 NAND2X1_1659 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n180_));
NAND2X1 NAND2X1_166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3413_), .B(AES_CORE_DATAPATH__abc_15863_new_n2890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3414_));
NAND2X1 NAND2X1_1660 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_));
NAND2X1 NAND2X1_1661 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n179_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n189_));
NAND2X1 NAND2X1_1662 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n191_));
NAND2X1 NAND2X1_1663 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n192_));
NAND2X1 NAND2X1_1664 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n191_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n193_));
NAND2X1 NAND2X1_1665 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n190_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n194_));
NAND2X1 NAND2X1_1666 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n197_));
NAND2X1 NAND2X1_1667 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n201_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n202_));
NAND2X1 NAND2X1_1668 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n202_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_));
NAND2X1 NAND2X1_1669 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n207_));
NAND2X1 NAND2X1_167 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3412_), .B(AES_CORE_DATAPATH__abc_15863_new_n3411_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3415_));
NAND2X1 NAND2X1_1670 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n212_));
NAND2X1 NAND2X1_1671 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n215_));
NAND2X1 NAND2X1_1672 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n217_));
NAND2X1 NAND2X1_1673 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n215_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n217_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n218_));
NAND2X1 NAND2X1_1674 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n222_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_));
NAND2X1 NAND2X1_1675 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n228_));
NAND2X1 NAND2X1_1676 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n229_));
NAND2X1 NAND2X1_1677 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n229_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n228_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n230_));
NAND2X1 NAND2X1_1678 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n233_));
NAND2X1 NAND2X1_1679 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n233_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n234_));
NAND2X1 NAND2X1_168 ( .A(AES_CORE_DATAPATH_col_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3423_));
NAND2X1 NAND2X1_1680 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n237_));
NAND2X1 NAND2X1_1681 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n239_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n241_));
NAND2X1 NAND2X1_1682 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n237_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n241_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n242_));
NAND2X1 NAND2X1_1683 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n243_));
NAND2X1 NAND2X1_1684 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n240_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n244_));
NAND2X1 NAND2X1_1685 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n236_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n245_));
NAND2X1 NAND2X1_1686 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n246_));
NAND2X1 NAND2X1_1687 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n247_));
NAND2X1 NAND2X1_1688 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n248_));
NAND2X1 NAND2X1_1689 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n249_));
NAND2X1 NAND2X1_169 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3434_), .B(AES_CORE_DATAPATH__abc_15863_new_n3433_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3437_));
NAND2X1 NAND2X1_1690 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n251_));
NAND2X1 NAND2X1_1691 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n252_));
NAND2X1 NAND2X1_1692 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n254_));
NAND2X1 NAND2X1_1693 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n258_));
NAND2X1 NAND2X1_1694 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n259_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n262_));
NAND2X1 NAND2X1_1695 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n253_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n264_));
NAND2X1 NAND2X1_1696 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n257_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n250_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n265_));
NAND2X1 NAND2X1_1697 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n263_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n268_));
NAND2X1 NAND2X1_1698 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n274_));
NAND2X1 NAND2X1_1699 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n275_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n269_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_));
NAND2X1 NAND2X1_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n176_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT_key_out_sel_1_));
NAND2X1 NAND2X1_170 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3437_), .B(AES_CORE_DATAPATH__abc_15863_new_n2900_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3438_));
NAND2X1 NAND2X1_1700 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n258_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n277_));
NAND2X1 NAND2X1_1701 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n280_));
NAND2X1 NAND2X1_1702 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n281_));
NAND2X1 NAND2X1_1703 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n157_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n284_));
NAND2X1 NAND2X1_1704 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n287_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n288_));
NAND2X1 NAND2X1_1705 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n295_));
NAND2X1 NAND2X1_1706 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n303_));
NAND2X1 NAND2X1_1707 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_));
NAND2X1 NAND2X1_1708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n315_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n317_));
NAND2X1 NAND2X1_1709 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n320_));
NAND2X1 NAND2X1_171 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3443_), .B(AES_CORE_DATAPATH__abc_15863_new_n3439_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3444_));
NAND2X1 NAND2X1_1710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n323_));
NAND2X1 NAND2X1_1711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n321_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n324_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_));
NAND2X1 NAND2X1_1712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n328_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n329_));
NAND2X1 NAND2X1_1713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n334_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_));
NAND2X1 NAND2X1_1714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n340_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_));
NAND2X1 NAND2X1_1715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n348_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_));
NAND2X1 NAND2X1_1716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_));
NAND2X1 NAND2X1_1717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_));
NAND2X1 NAND2X1_1718 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n370_));
NAND2X1 NAND2X1_1719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n374_));
NAND2X1 NAND2X1_172 ( .A(AES_CORE_DATAPATH_col_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3445_));
NAND2X1 NAND2X1_1720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n375_));
NAND2X1 NAND2X1_1721 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n376_));
NAND2X1 NAND2X1_1722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n376_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n382_));
NAND2X1 NAND2X1_1723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n383_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_));
NAND2X1 NAND2X1_1724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n393_));
NAND2X1 NAND2X1_1725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n405_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n404_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n406_));
NAND2X1 NAND2X1_1726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n408_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n410_));
NAND2X1 NAND2X1_1727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_));
NAND2X1 NAND2X1_1728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n421_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n417_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_));
NAND2X1 NAND2X1_1729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n397_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n396_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n427_));
NAND2X1 NAND2X1_173 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3448_));
NAND2X1 NAND2X1_1730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n429_));
NAND2X1 NAND2X1_1731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n431_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n435_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n436_));
NAND2X1 NAND2X1_1732 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n442_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n444_));
NAND2X1 NAND2X1_1733 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n438_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n450_));
NAND2X1 NAND2X1_1734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_));
NAND2X1 NAND2X1_1735 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n456_));
NAND2X1 NAND2X1_1736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n434_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n466_));
NAND2X1 NAND2X1_1737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n467_));
NAND2X1 NAND2X1_1738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n463_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n469_));
NAND2X1 NAND2X1_1739 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n471_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_));
NAND2X1 NAND2X1_174 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3457_), .B(AES_CORE_DATAPATH__abc_15863_new_n2911_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3458_));
NAND2X1 NAND2X1_1740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n489_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n486_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_));
NAND2X1 NAND2X1_1741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_));
NAND2X1 NAND2X1_1742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n377_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_));
NAND2X1 NAND2X1_175 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3456_), .B(AES_CORE_DATAPATH__abc_15863_new_n3455_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3459_));
NAND2X1 NAND2X1_176 ( .A(AES_CORE_DATAPATH_col_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3467_));
NAND2X1 NAND2X1_177 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3478_), .B(AES_CORE_DATAPATH__abc_15863_new_n3477_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3481_));
NAND2X1 NAND2X1_178 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3481_), .B(AES_CORE_DATAPATH__abc_15863_new_n2920_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3482_));
NAND2X1 NAND2X1_179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3487_), .B(AES_CORE_DATAPATH__abc_15863_new_n3483_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3488_));
NAND2X1 NAND2X1_18 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n212_));
NAND2X1 NAND2X1_180 ( .A(AES_CORE_DATAPATH_col_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3489_));
NAND2X1 NAND2X1_181 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3500_), .B(AES_CORE_DATAPATH__abc_15863_new_n3499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3501_));
NAND2X1 NAND2X1_182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3501_), .B(AES_CORE_DATAPATH__abc_15863_new_n2930_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3502_));
NAND2X1 NAND2X1_183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3509_), .B(AES_CORE_DATAPATH__abc_15863_new_n3505_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3510_));
NAND2X1 NAND2X1_184 ( .A(AES_CORE_DATAPATH_col_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3511_));
NAND2X1 NAND2X1_185 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3522_), .B(AES_CORE_DATAPATH__abc_15863_new_n3521_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3525_));
NAND2X1 NAND2X1_186 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3525_), .B(AES_CORE_DATAPATH__abc_15863_new_n2940_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3526_));
NAND2X1 NAND2X1_187 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3531_), .B(AES_CORE_DATAPATH__abc_15863_new_n3527_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3532_));
NAND2X1 NAND2X1_188 ( .A(AES_CORE_DATAPATH_col_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3533_));
NAND2X1 NAND2X1_189 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3536_));
NAND2X1 NAND2X1_19 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_0_));
NAND2X1 NAND2X1_190 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3545_), .B(AES_CORE_DATAPATH__abc_15863_new_n2951_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3546_));
NAND2X1 NAND2X1_191 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3544_), .B(AES_CORE_DATAPATH__abc_15863_new_n3543_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3547_));
NAND2X1 NAND2X1_192 ( .A(AES_CORE_DATAPATH_col_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3555_));
NAND2X1 NAND2X1_193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3566_), .B(AES_CORE_DATAPATH__abc_15863_new_n3565_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3569_));
NAND2X1 NAND2X1_194 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3569_), .B(AES_CORE_DATAPATH__abc_15863_new_n2963_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3570_));
NAND2X1 NAND2X1_195 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3575_), .B(AES_CORE_DATAPATH__abc_15863_new_n3571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3576_));
NAND2X1 NAND2X1_196 ( .A(AES_CORE_DATAPATH_col_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3577_));
NAND2X1 NAND2X1_197 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3580_));
NAND2X1 NAND2X1_198 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3589_), .B(AES_CORE_DATAPATH__abc_15863_new_n2973_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3590_));
NAND2X1 NAND2X1_199 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3588_), .B(AES_CORE_DATAPATH__abc_15863_new_n3587_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3591_));
NAND2X1 NAND2X1_2 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n77_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n80_), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt));
NAND2X1 NAND2X1_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n176_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_1_));
NAND2X1 NAND2X1_200 ( .A(AES_CORE_DATAPATH_col_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3599_));
NAND2X1 NAND2X1_201 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3611_), .B(AES_CORE_DATAPATH__abc_15863_new_n2984_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3612_));
NAND2X1 NAND2X1_202 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3610_), .B(AES_CORE_DATAPATH__abc_15863_new_n3609_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3613_));
NAND2X1 NAND2X1_203 ( .A(AES_CORE_DATAPATH_col_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3621_));
NAND2X1 NAND2X1_204 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3624_));
NAND2X1 NAND2X1_205 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3633_), .B(AES_CORE_DATAPATH__abc_15863_new_n2997_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3634_));
NAND2X1 NAND2X1_206 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3632_), .B(AES_CORE_DATAPATH__abc_15863_new_n3631_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3635_));
NAND2X1 NAND2X1_207 ( .A(AES_CORE_DATAPATH_col_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3643_));
NAND2X1 NAND2X1_208 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3654_), .B(AES_CORE_DATAPATH__abc_15863_new_n3653_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3657_));
NAND2X1 NAND2X1_209 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3657_), .B(AES_CORE_DATAPATH__abc_15863_new_n3009_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3658_));
NAND2X1 NAND2X1_21 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2459_));
NAND2X1 NAND2X1_210 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3663_), .B(AES_CORE_DATAPATH__abc_15863_new_n3659_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3664_));
NAND2X1 NAND2X1_211 ( .A(AES_CORE_DATAPATH_col_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3665_));
NAND2X1 NAND2X1_212 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3676_), .B(AES_CORE_DATAPATH__abc_15863_new_n3675_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3677_));
NAND2X1 NAND2X1_213 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3677_), .B(AES_CORE_DATAPATH__abc_15863_new_n3019_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3678_));
NAND2X1 NAND2X1_214 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3685_), .B(AES_CORE_DATAPATH__abc_15863_new_n3681_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3686_));
NAND2X1 NAND2X1_215 ( .A(AES_CORE_DATAPATH_col_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3687_));
NAND2X1 NAND2X1_216 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3690_));
NAND2X1 NAND2X1_217 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3699_), .B(AES_CORE_DATAPATH__abc_15863_new_n3029_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3700_));
NAND2X1 NAND2X1_218 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3698_), .B(AES_CORE_DATAPATH__abc_15863_new_n3697_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3701_));
NAND2X1 NAND2X1_219 ( .A(AES_CORE_DATAPATH_col_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3709_));
NAND2X1 NAND2X1_22 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2464_));
NAND2X1 NAND2X1_220 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3720_), .B(AES_CORE_DATAPATH__abc_15863_new_n3719_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3723_));
NAND2X1 NAND2X1_221 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3723_), .B(AES_CORE_DATAPATH__abc_15863_new_n3040_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3724_));
NAND2X1 NAND2X1_222 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3729_), .B(AES_CORE_DATAPATH__abc_15863_new_n3725_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3730_));
NAND2X1 NAND2X1_223 ( .A(AES_CORE_DATAPATH_col_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3731_));
NAND2X1 NAND2X1_224 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3734_));
NAND2X1 NAND2X1_225 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3743_), .B(AES_CORE_DATAPATH__abc_15863_new_n3050_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3744_));
NAND2X1 NAND2X1_226 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3742_), .B(AES_CORE_DATAPATH__abc_15863_new_n3741_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3745_));
NAND2X1 NAND2X1_227 ( .A(AES_CORE_DATAPATH_col_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3753_));
NAND2X1 NAND2X1_228 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .B(AES_CORE_DATAPATH__abc_15863_new_n3085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3756_));
NAND2X1 NAND2X1_229 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3765_), .B(AES_CORE_DATAPATH__abc_15863_new_n3060_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3766_));
NAND2X1 NAND2X1_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2465_), .B(AES_CORE_DATAPATH__abc_15863_new_n2464_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2466_));
NAND2X1 NAND2X1_230 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3764_), .B(AES_CORE_DATAPATH__abc_15863_new_n3763_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3767_));
NAND2X1 NAND2X1_231 ( .A(AES_CORE_DATAPATH_col_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3775_));
NAND2X1 NAND2X1_232 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3786_), .B(AES_CORE_DATAPATH__abc_15863_new_n3785_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3789_));
NAND2X1 NAND2X1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3789_), .B(AES_CORE_DATAPATH__abc_15863_new_n3069_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3790_));
NAND2X1 NAND2X1_234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3795_), .B(AES_CORE_DATAPATH__abc_15863_new_n3791_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3796_));
NAND2X1 NAND2X1_235 ( .A(AES_CORE_DATAPATH_col_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3797_));
NAND2X1 NAND2X1_236 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3799_));
NAND2X1 NAND2X1_237 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3801_));
NAND2X1 NAND2X1_238 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3803_));
NAND2X1 NAND2X1_239 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3805_));
NAND2X1 NAND2X1_24 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2471_));
NAND2X1 NAND2X1_240 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3807_));
NAND2X1 NAND2X1_241 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3809_));
NAND2X1 NAND2X1_242 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3811_));
NAND2X1 NAND2X1_243 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3813_));
NAND2X1 NAND2X1_244 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3815_));
NAND2X1 NAND2X1_245 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3817_));
NAND2X1 NAND2X1_246 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3819_));
NAND2X1 NAND2X1_247 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3821_));
NAND2X1 NAND2X1_248 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3823_));
NAND2X1 NAND2X1_249 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3825_));
NAND2X1 NAND2X1_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2472_), .B(AES_CORE_DATAPATH__abc_15863_new_n2471_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2473_));
NAND2X1 NAND2X1_250 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3827_));
NAND2X1 NAND2X1_251 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3829_));
NAND2X1 NAND2X1_252 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3831_));
NAND2X1 NAND2X1_253 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3833_));
NAND2X1 NAND2X1_254 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3835_));
NAND2X1 NAND2X1_255 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3837_));
NAND2X1 NAND2X1_256 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3839_));
NAND2X1 NAND2X1_257 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3841_));
NAND2X1 NAND2X1_258 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3843_));
NAND2X1 NAND2X1_259 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3845_));
NAND2X1 NAND2X1_26 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2470_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2475_));
NAND2X1 NAND2X1_260 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3847_));
NAND2X1 NAND2X1_261 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3849_));
NAND2X1 NAND2X1_262 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3851_));
NAND2X1 NAND2X1_263 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3853_));
NAND2X1 NAND2X1_264 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3855_));
NAND2X1 NAND2X1_265 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3857_));
NAND2X1 NAND2X1_266 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3859_));
NAND2X1 NAND2X1_267 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3861_));
NAND2X1 NAND2X1_268 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH_rk_out_sel));
NAND2X1 NAND2X1_269 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3868_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3869_));
NAND2X1 NAND2X1_27 ( .A(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2476_));
NAND2X1 NAND2X1_270 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3871_));
NAND2X1 NAND2X1_271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3873_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3874_));
NAND2X1 NAND2X1_272 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3876_));
NAND2X1 NAND2X1_273 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3878_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3879_));
NAND2X1 NAND2X1_274 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3881_));
NAND2X1 NAND2X1_275 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3883_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3884_));
NAND2X1 NAND2X1_276 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3886_));
NAND2X1 NAND2X1_277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3888_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3889_));
NAND2X1 NAND2X1_278 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3891_));
NAND2X1 NAND2X1_279 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3893_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3894_));
NAND2X1 NAND2X1_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2477_), .B(AES_CORE_DATAPATH__abc_15863_new_n2476_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2478_));
NAND2X1 NAND2X1_280 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3896_));
NAND2X1 NAND2X1_281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3898_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3899_));
NAND2X1 NAND2X1_282 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3901_));
NAND2X1 NAND2X1_283 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3903_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3904_));
NAND2X1 NAND2X1_284 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3906_));
NAND2X1 NAND2X1_285 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3908_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3909_));
NAND2X1 NAND2X1_286 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3911_));
NAND2X1 NAND2X1_287 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3913_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3914_));
NAND2X1 NAND2X1_288 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3916_));
NAND2X1 NAND2X1_289 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3918_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3919_));
NAND2X1 NAND2X1_29 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2489_), .B(AES_CORE_DATAPATH__abc_15863_new_n2491_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2492_));
NAND2X1 NAND2X1_290 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3921_));
NAND2X1 NAND2X1_291 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3923_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3924_));
NAND2X1 NAND2X1_292 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3926_));
NAND2X1 NAND2X1_293 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3928_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3929_));
NAND2X1 NAND2X1_294 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3931_));
NAND2X1 NAND2X1_295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3933_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3934_));
NAND2X1 NAND2X1_296 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3936_));
NAND2X1 NAND2X1_297 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3938_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3939_));
NAND2X1 NAND2X1_298 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3941_));
NAND2X1 NAND2X1_299 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3943_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3944_));
NAND2X1 NAND2X1_3 ( .A(AES_CORE_CONTROL_UNIT_rd_count_1_), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n83_));
NAND2X1 NAND2X1_30 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2503_), .B(AES_CORE_DATAPATH__abc_15863_new_n2505_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2506_));
NAND2X1 NAND2X1_300 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3946_));
NAND2X1 NAND2X1_301 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3948_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3949_));
NAND2X1 NAND2X1_302 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3951_));
NAND2X1 NAND2X1_303 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3953_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3954_));
NAND2X1 NAND2X1_304 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3956_));
NAND2X1 NAND2X1_305 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3958_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3959_));
NAND2X1 NAND2X1_306 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3961_));
NAND2X1 NAND2X1_307 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3963_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3964_));
NAND2X1 NAND2X1_308 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3966_));
NAND2X1 NAND2X1_309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3968_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3969_));
NAND2X1 NAND2X1_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2577_), .B(AES_CORE_DATAPATH__abc_15863_new_n2579_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2580_));
NAND2X1 NAND2X1_310 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3971_));
NAND2X1 NAND2X1_311 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3973_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3974_));
NAND2X1 NAND2X1_312 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3976_));
NAND2X1 NAND2X1_313 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3978_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3979_));
NAND2X1 NAND2X1_314 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3981_));
NAND2X1 NAND2X1_315 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3983_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3984_));
NAND2X1 NAND2X1_316 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3986_));
NAND2X1 NAND2X1_317 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3988_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3989_));
NAND2X1 NAND2X1_318 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3991_));
NAND2X1 NAND2X1_319 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3993_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3994_));
NAND2X1 NAND2X1_32 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2591_), .B(AES_CORE_DATAPATH__abc_15863_new_n2593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2594_));
NAND2X1 NAND2X1_320 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3996_));
NAND2X1 NAND2X1_321 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3998_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3999_));
NAND2X1 NAND2X1_322 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4001_));
NAND2X1 NAND2X1_323 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4003_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4004_));
NAND2X1 NAND2X1_324 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4006_));
NAND2X1 NAND2X1_325 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4008_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4009_));
NAND2X1 NAND2X1_326 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4011_));
NAND2X1 NAND2X1_327 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4013_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4014_));
NAND2X1 NAND2X1_328 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4016_));
NAND2X1 NAND2X1_329 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4018_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4019_));
NAND2X1 NAND2X1_33 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2605_), .B(AES_CORE_DATAPATH__abc_15863_new_n2607_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2608_));
NAND2X1 NAND2X1_330 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4021_));
NAND2X1 NAND2X1_331 ( .A(\key_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4023_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4024_));
NAND2X1 NAND2X1_332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4025_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4026_));
NAND2X1 NAND2X1_333 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n3866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4028_));
NAND2X1 NAND2X1_334 ( .A(AES_CORE_DATAPATH_key_en_pp1_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2712_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4031_));
NAND2X1 NAND2X1_335 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4038_));
NAND2X1 NAND2X1_336 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4040_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4041_));
NAND2X1 NAND2X1_337 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4043_));
NAND2X1 NAND2X1_338 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4045_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4046_));
NAND2X1 NAND2X1_339 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4048_));
NAND2X1 NAND2X1_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2613_), .B(AES_CORE_DATAPATH__abc_15863_new_n2615_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2616_));
NAND2X1 NAND2X1_340 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4050_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4051_));
NAND2X1 NAND2X1_341 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4053_));
NAND2X1 NAND2X1_342 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4055_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4056_));
NAND2X1 NAND2X1_343 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4058_));
NAND2X1 NAND2X1_344 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4060_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4061_));
NAND2X1 NAND2X1_345 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4063_));
NAND2X1 NAND2X1_346 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4065_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4066_));
NAND2X1 NAND2X1_347 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4068_));
NAND2X1 NAND2X1_348 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4070_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4071_));
NAND2X1 NAND2X1_349 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4073_));
NAND2X1 NAND2X1_35 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2621_), .B(AES_CORE_DATAPATH__abc_15863_new_n2623_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2624_));
NAND2X1 NAND2X1_350 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4075_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4076_));
NAND2X1 NAND2X1_351 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4078_));
NAND2X1 NAND2X1_352 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4080_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4081_));
NAND2X1 NAND2X1_353 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4083_));
NAND2X1 NAND2X1_354 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4085_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4086_));
NAND2X1 NAND2X1_355 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4088_));
NAND2X1 NAND2X1_356 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4090_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4091_));
NAND2X1 NAND2X1_357 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4093_));
NAND2X1 NAND2X1_358 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4095_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4096_));
NAND2X1 NAND2X1_359 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4098_));
NAND2X1 NAND2X1_36 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2635_), .B(AES_CORE_DATAPATH__abc_15863_new_n2637_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2638_));
NAND2X1 NAND2X1_360 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4100_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4101_));
NAND2X1 NAND2X1_361 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4103_));
NAND2X1 NAND2X1_362 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4105_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4106_));
NAND2X1 NAND2X1_363 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4108_));
NAND2X1 NAND2X1_364 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4110_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4111_));
NAND2X1 NAND2X1_365 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4113_));
NAND2X1 NAND2X1_366 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4115_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4116_));
NAND2X1 NAND2X1_367 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4118_));
NAND2X1 NAND2X1_368 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4120_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4121_));
NAND2X1 NAND2X1_369 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4123_));
NAND2X1 NAND2X1_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2649_), .B(AES_CORE_DATAPATH__abc_15863_new_n2651_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2652_));
NAND2X1 NAND2X1_370 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4125_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4126_));
NAND2X1 NAND2X1_371 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4128_));
NAND2X1 NAND2X1_372 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4130_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4131_));
NAND2X1 NAND2X1_373 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4133_));
NAND2X1 NAND2X1_374 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4135_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4136_));
NAND2X1 NAND2X1_375 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4138_));
NAND2X1 NAND2X1_376 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4140_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4141_));
NAND2X1 NAND2X1_377 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4143_));
NAND2X1 NAND2X1_378 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4145_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4146_));
NAND2X1 NAND2X1_379 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4148_));
NAND2X1 NAND2X1_38 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2663_), .B(AES_CORE_DATAPATH__abc_15863_new_n2665_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2666_));
NAND2X1 NAND2X1_380 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4150_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4151_));
NAND2X1 NAND2X1_381 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4153_));
NAND2X1 NAND2X1_382 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4155_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4156_));
NAND2X1 NAND2X1_383 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4158_));
NAND2X1 NAND2X1_384 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4160_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4161_));
NAND2X1 NAND2X1_385 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4163_));
NAND2X1 NAND2X1_386 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4165_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4166_));
NAND2X1 NAND2X1_387 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4168_));
NAND2X1 NAND2X1_388 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4170_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4171_));
NAND2X1 NAND2X1_389 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4173_));
NAND2X1 NAND2X1_39 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2671_), .B(AES_CORE_DATAPATH__abc_15863_new_n2673_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2674_));
NAND2X1 NAND2X1_390 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4175_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4176_));
NAND2X1 NAND2X1_391 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4178_));
NAND2X1 NAND2X1_392 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4180_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4181_));
NAND2X1 NAND2X1_393 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4183_));
NAND2X1 NAND2X1_394 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4185_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4186_));
NAND2X1 NAND2X1_395 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4188_));
NAND2X1 NAND2X1_396 ( .A(\key_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4023_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4190_));
NAND2X1 NAND2X1_397 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4191_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4192_));
NAND2X1 NAND2X1_398 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4194_));
NAND2X1 NAND2X1_399 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n4196_));
NAND2X1 NAND2X1_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n85_));
NAND2X1 NAND2X1_40 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2685_), .B(AES_CORE_DATAPATH__abc_15863_new_n2687_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2688_));
NAND2X1 NAND2X1_400 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n4230_));
NAND2X1 NAND2X1_401 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4231_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4232_));
NAND2X1 NAND2X1_402 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4236_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4237_));
NAND2X1 NAND2X1_403 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4241_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4242_));
NAND2X1 NAND2X1_404 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4246_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4247_));
NAND2X1 NAND2X1_405 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4251_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4252_));
NAND2X1 NAND2X1_406 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4256_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4257_));
NAND2X1 NAND2X1_407 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4279_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4280_));
NAND2X1 NAND2X1_408 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4284_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4285_));
NAND2X1 NAND2X1_409 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4289_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4290_));
NAND2X1 NAND2X1_41 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2705_), .B(AES_CORE_DATAPATH__abc_15863_new_n2707_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2708_));
NAND2X1 NAND2X1_410 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4294_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4295_));
NAND2X1 NAND2X1_411 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4299_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4300_));
NAND2X1 NAND2X1_412 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4304_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4305_));
NAND2X1 NAND2X1_413 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4309_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4310_));
NAND2X1 NAND2X1_414 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4314_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4315_));
NAND2X1 NAND2X1_415 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4319_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4320_));
NAND2X1 NAND2X1_416 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4324_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4325_));
NAND2X1 NAND2X1_417 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4329_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4330_));
NAND2X1 NAND2X1_418 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4334_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4335_));
NAND2X1 NAND2X1_419 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4339_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4340_));
NAND2X1 NAND2X1_42 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2720_), .B(AES_CORE_DATAPATH__abc_15863_new_n2719_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2721_));
NAND2X1 NAND2X1_420 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4344_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4345_));
NAND2X1 NAND2X1_421 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4349_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4350_));
NAND2X1 NAND2X1_422 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4354_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4355_));
NAND2X1 NAND2X1_423 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4359_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4360_));
NAND2X1 NAND2X1_424 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4364_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4365_));
NAND2X1 NAND2X1_425 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4369_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4370_));
NAND2X1 NAND2X1_426 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n4376_));
NAND2X1 NAND2X1_427 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4233_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4443_));
NAND2X1 NAND2X1_428 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4445_));
NAND2X1 NAND2X1_429 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4238_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4447_));
NAND2X1 NAND2X1_43 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2727_), .B(AES_CORE_DATAPATH__abc_15863_new_n2726_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2728_));
NAND2X1 NAND2X1_430 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4449_));
NAND2X1 NAND2X1_431 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4243_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4451_));
NAND2X1 NAND2X1_432 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4453_));
NAND2X1 NAND2X1_433 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4248_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4455_));
NAND2X1 NAND2X1_434 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4457_));
NAND2X1 NAND2X1_435 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4253_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4459_));
NAND2X1 NAND2X1_436 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4461_));
NAND2X1 NAND2X1_437 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4258_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4463_));
NAND2X1 NAND2X1_438 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4465_));
NAND2X1 NAND2X1_439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4261_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4467_));
NAND2X1 NAND2X1_44 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2711_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2730_));
NAND2X1 NAND2X1_440 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4469_));
NAND2X1 NAND2X1_441 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4264_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4471_));
NAND2X1 NAND2X1_442 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4473_));
NAND2X1 NAND2X1_443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4267_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4475_));
NAND2X1 NAND2X1_444 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4477_));
NAND2X1 NAND2X1_445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4270_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4479_));
NAND2X1 NAND2X1_446 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4481_));
NAND2X1 NAND2X1_447 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4273_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4483_));
NAND2X1 NAND2X1_448 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4485_));
NAND2X1 NAND2X1_449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4276_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4487_));
NAND2X1 NAND2X1_45 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2730_), .B(AES_CORE_DATAPATH__abc_15863_new_n2739_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2740_));
NAND2X1 NAND2X1_450 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4489_));
NAND2X1 NAND2X1_451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4281_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4491_));
NAND2X1 NAND2X1_452 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4493_));
NAND2X1 NAND2X1_453 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4286_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4495_));
NAND2X1 NAND2X1_454 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4497_));
NAND2X1 NAND2X1_455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4291_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4499_));
NAND2X1 NAND2X1_456 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4501_));
NAND2X1 NAND2X1_457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4296_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4503_));
NAND2X1 NAND2X1_458 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4505_));
NAND2X1 NAND2X1_459 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4301_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4507_));
NAND2X1 NAND2X1_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2749_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2750_));
NAND2X1 NAND2X1_460 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4509_));
NAND2X1 NAND2X1_461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4306_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4511_));
NAND2X1 NAND2X1_462 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4513_));
NAND2X1 NAND2X1_463 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4311_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4515_));
NAND2X1 NAND2X1_464 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4517_));
NAND2X1 NAND2X1_465 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4316_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4519_));
NAND2X1 NAND2X1_466 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4521_));
NAND2X1 NAND2X1_467 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4321_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4523_));
NAND2X1 NAND2X1_468 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4525_));
NAND2X1 NAND2X1_469 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4326_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4527_));
NAND2X1 NAND2X1_47 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2750_), .B(AES_CORE_DATAPATH__abc_15863_new_n2748_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2751_));
NAND2X1 NAND2X1_470 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4529_));
NAND2X1 NAND2X1_471 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4331_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4531_));
NAND2X1 NAND2X1_472 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4533_));
NAND2X1 NAND2X1_473 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4336_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4535_));
NAND2X1 NAND2X1_474 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4537_));
NAND2X1 NAND2X1_475 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4341_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4539_));
NAND2X1 NAND2X1_476 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4541_));
NAND2X1 NAND2X1_477 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4346_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4543_));
NAND2X1 NAND2X1_478 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4545_));
NAND2X1 NAND2X1_479 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4351_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4547_));
NAND2X1 NAND2X1_48 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2762_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2763_));
NAND2X1 NAND2X1_480 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4549_));
NAND2X1 NAND2X1_481 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4356_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4551_));
NAND2X1 NAND2X1_482 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4553_));
NAND2X1 NAND2X1_483 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4361_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4555_));
NAND2X1 NAND2X1_484 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4557_));
NAND2X1 NAND2X1_485 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4366_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4559_));
NAND2X1 NAND2X1_486 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4561_));
NAND2X1 NAND2X1_487 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4371_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4563_));
NAND2X1 NAND2X1_488 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4565_));
NAND2X1 NAND2X1_489 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4373_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4567_));
NAND2X1 NAND2X1_49 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2763_), .B(AES_CORE_DATAPATH__abc_15863_new_n2761_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2764_));
NAND2X1 NAND2X1_490 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4442_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4569_));
NAND2X1 NAND2X1_491 ( .A(AES_CORE_DATAPATH_col_0__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4572_));
NAND2X1 NAND2X1_492 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_sel_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4574_));
NAND2X1 NAND2X1_493 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_sel_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4577_));
NAND2X1 NAND2X1_494 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3111_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4586_));
NAND2X1 NAND2X1_495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4575_), .B(AES_CORE_DATAPATH__abc_15863_new_n4584_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4587_));
NAND2X1 NAND2X1_496 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4595_));
NAND2X1 NAND2X1_497 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4602_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4603_));
NAND2X1 NAND2X1_498 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4612_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4613_));
NAND2X1 NAND2X1_499 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4614_));
NAND2X1 NAND2X1_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n78_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n79_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_));
NAND2X1 NAND2X1_50 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2768_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2769_));
NAND2X1 NAND2X1_500 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4610_), .B(AES_CORE_DATAPATH__abc_15863_new_n4616_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4617_));
NAND2X1 NAND2X1_501 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4627_));
NAND2X1 NAND2X1_502 ( .A(AES_CORE_DATAPATH_col_0__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4633_));
NAND2X1 NAND2X1_503 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4643_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4644_));
NAND2X1 NAND2X1_504 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4649_));
NAND2X1 NAND2X1_505 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3128_), .B(AES_CORE_DATAPATH__abc_15863_new_n2751_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4653_));
NAND2X1 NAND2X1_506 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4651_), .B(AES_CORE_DATAPATH__abc_15863_new_n4659_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4660_));
NAND2X1 NAND2X1_507 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4665_));
NAND2X1 NAND2X1_508 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3134_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4668_));
NAND2X1 NAND2X1_509 ( .A(AES_CORE_DATAPATH_col_0__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4672_));
NAND2X1 NAND2X1_51 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2769_), .B(AES_CORE_DATAPATH__abc_15863_new_n2773_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2774_));
NAND2X1 NAND2X1_510 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4680_));
NAND2X1 NAND2X1_511 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4684_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4685_));
NAND2X1 NAND2X1_512 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4694_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4695_));
NAND2X1 NAND2X1_513 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4696_));
NAND2X1 NAND2X1_514 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4692_), .B(AES_CORE_DATAPATH__abc_15863_new_n4698_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4699_));
NAND2X1 NAND2X1_515 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4704_));
NAND2X1 NAND2X1_516 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3156_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4707_));
NAND2X1 NAND2X1_517 ( .A(AES_CORE_DATAPATH_col_0__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4711_));
NAND2X1 NAND2X1_518 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3171_), .B(AES_CORE_DATAPATH__abc_15863_new_n2774_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4715_));
NAND2X1 NAND2X1_519 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4724_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4725_));
NAND2X1 NAND2X1_52 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2778_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2779_));
NAND2X1 NAND2X1_520 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4730_));
NAND2X1 NAND2X1_521 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4732_), .B(AES_CORE_DATAPATH__abc_15863_new_n4736_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4737_));
NAND2X1 NAND2X1_522 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4742_));
NAND2X1 NAND2X1_523 ( .A(AES_CORE_DATAPATH_col_0__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4751_));
NAND2X1 NAND2X1_524 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4759_));
NAND2X1 NAND2X1_525 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4770_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4771_));
NAND2X1 NAND2X1_526 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[4] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4772_));
NAND2X1 NAND2X1_527 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4768_), .B(AES_CORE_DATAPATH__abc_15863_new_n4774_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4775_));
NAND2X1 NAND2X1_528 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4780_));
NAND2X1 NAND2X1_529 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3201_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4783_));
NAND2X1 NAND2X1_53 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2779_), .B(AES_CORE_DATAPATH__abc_15863_new_n2783_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2784_));
NAND2X1 NAND2X1_530 ( .A(AES_CORE_DATAPATH_col_0__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4787_));
NAND2X1 NAND2X1_531 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4795_));
NAND2X1 NAND2X1_532 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4799_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4800_));
NAND2X1 NAND2X1_533 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4809_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4810_));
NAND2X1 NAND2X1_534 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[5] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4811_));
NAND2X1 NAND2X1_535 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4807_), .B(AES_CORE_DATAPATH__abc_15863_new_n4813_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4814_));
NAND2X1 NAND2X1_536 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4819_));
NAND2X1 NAND2X1_537 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3223_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4822_));
NAND2X1 NAND2X1_538 ( .A(AES_CORE_DATAPATH_col_0__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4826_));
NAND2X1 NAND2X1_539 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4834_));
NAND2X1 NAND2X1_54 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2792_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2793_));
NAND2X1 NAND2X1_540 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4845_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4846_));
NAND2X1 NAND2X1_541 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4843_), .B(AES_CORE_DATAPATH__abc_15863_new_n4848_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4849_));
NAND2X1 NAND2X1_542 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4854_));
NAND2X1 NAND2X1_543 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3245_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4857_));
NAND2X1 NAND2X1_544 ( .A(AES_CORE_DATAPATH_col_0__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4861_));
NAND2X1 NAND2X1_545 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4871_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4872_));
NAND2X1 NAND2X1_546 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[7] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4877_));
NAND2X1 NAND2X1_547 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3261_), .B(AES_CORE_DATAPATH__abc_15863_new_n2815_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4881_));
NAND2X1 NAND2X1_548 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4879_), .B(AES_CORE_DATAPATH__abc_15863_new_n4887_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4888_));
NAND2X1 NAND2X1_549 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4893_));
NAND2X1 NAND2X1_55 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2793_), .B(AES_CORE_DATAPATH__abc_15863_new_n2791_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2794_));
NAND2X1 NAND2X1_550 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3267_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4896_));
NAND2X1 NAND2X1_551 ( .A(AES_CORE_DATAPATH_col_0__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4900_));
NAND2X1 NAND2X1_552 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4908_));
NAND2X1 NAND2X1_553 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4919_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4920_));
NAND2X1 NAND2X1_554 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4917_), .B(AES_CORE_DATAPATH__abc_15863_new_n4922_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4923_));
NAND2X1 NAND2X1_555 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4928_));
NAND2X1 NAND2X1_556 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3289_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4931_));
NAND2X1 NAND2X1_557 ( .A(AES_CORE_DATAPATH_col_0__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4935_));
NAND2X1 NAND2X1_558 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3303_), .B(AES_CORE_DATAPATH__abc_15863_new_n2840_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4939_));
NAND2X1 NAND2X1_559 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4948_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4949_));
NAND2X1 NAND2X1_56 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2798_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2799_));
NAND2X1 NAND2X1_560 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[9] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4954_));
NAND2X1 NAND2X1_561 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4956_), .B(AES_CORE_DATAPATH__abc_15863_new_n4960_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4961_));
NAND2X1 NAND2X1_562 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4966_));
NAND2X1 NAND2X1_563 ( .A(AES_CORE_DATAPATH_col_0__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4974_));
NAND2X1 NAND2X1_564 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4982_));
NAND2X1 NAND2X1_565 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n4986_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4987_));
NAND2X1 NAND2X1_566 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4996_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4997_));
NAND2X1 NAND2X1_567 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[10] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n4998_));
NAND2X1 NAND2X1_568 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4994_), .B(AES_CORE_DATAPATH__abc_15863_new_n5000_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5001_));
NAND2X1 NAND2X1_569 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5006_));
NAND2X1 NAND2X1_57 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2799_), .B(AES_CORE_DATAPATH__abc_15863_new_n2803_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2804_));
NAND2X1 NAND2X1_570 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3333_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5009_));
NAND2X1 NAND2X1_571 ( .A(AES_CORE_DATAPATH_col_0__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5013_));
NAND2X1 NAND2X1_572 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3347_), .B(AES_CORE_DATAPATH__abc_15863_new_n2860_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5017_));
NAND2X1 NAND2X1_573 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5026_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5027_));
NAND2X1 NAND2X1_574 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[11] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5032_));
NAND2X1 NAND2X1_575 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5034_), .B(AES_CORE_DATAPATH__abc_15863_new_n5038_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5039_));
NAND2X1 NAND2X1_576 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5044_));
NAND2X1 NAND2X1_577 ( .A(AES_CORE_DATAPATH_col_0__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5052_));
NAND2X1 NAND2X1_578 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5060_));
NAND2X1 NAND2X1_579 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5064_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5065_));
NAND2X1 NAND2X1_58 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2813_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2814_));
NAND2X1 NAND2X1_580 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5074_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5075_));
NAND2X1 NAND2X1_581 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[12] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5076_));
NAND2X1 NAND2X1_582 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5072_), .B(AES_CORE_DATAPATH__abc_15863_new_n5078_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5079_));
NAND2X1 NAND2X1_583 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5084_));
NAND2X1 NAND2X1_584 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3377_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5087_));
NAND2X1 NAND2X1_585 ( .A(AES_CORE_DATAPATH_col_0__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5091_));
NAND2X1 NAND2X1_586 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3391_), .B(AES_CORE_DATAPATH__abc_15863_new_n2880_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5095_));
NAND2X1 NAND2X1_587 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5104_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5105_));
NAND2X1 NAND2X1_588 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[13] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5110_));
NAND2X1 NAND2X1_589 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5112_), .B(AES_CORE_DATAPATH__abc_15863_new_n5116_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5117_));
NAND2X1 NAND2X1_59 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2814_), .B(AES_CORE_DATAPATH__abc_15863_new_n2812_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2815_));
NAND2X1 NAND2X1_590 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5122_));
NAND2X1 NAND2X1_591 ( .A(AES_CORE_DATAPATH_col_0__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5130_));
NAND2X1 NAND2X1_592 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5138_));
NAND2X1 NAND2X1_593 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5149_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5150_));
NAND2X1 NAND2X1_594 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[14] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5151_));
NAND2X1 NAND2X1_595 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5147_), .B(AES_CORE_DATAPATH__abc_15863_new_n5153_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5154_));
NAND2X1 NAND2X1_596 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5159_));
NAND2X1 NAND2X1_597 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3421_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5162_));
NAND2X1 NAND2X1_598 ( .A(AES_CORE_DATAPATH_col_0__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5166_));
NAND2X1 NAND2X1_599 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3435_), .B(AES_CORE_DATAPATH__abc_15863_new_n2900_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5170_));
NAND2X1 NAND2X1_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n98_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n99_));
NAND2X1 NAND2X1_60 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2826_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2827_));
NAND2X1 NAND2X1_600 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5179_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5180_));
NAND2X1 NAND2X1_601 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[15] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5185_));
NAND2X1 NAND2X1_602 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5187_), .B(AES_CORE_DATAPATH__abc_15863_new_n5191_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5192_));
NAND2X1 NAND2X1_603 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5197_));
NAND2X1 NAND2X1_604 ( .A(AES_CORE_DATAPATH_col_0__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5205_));
NAND2X1 NAND2X1_605 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5213_));
NAND2X1 NAND2X1_606 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5217_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5218_));
NAND2X1 NAND2X1_607 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5227_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5228_));
NAND2X1 NAND2X1_608 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[16] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5229_));
NAND2X1 NAND2X1_609 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5225_), .B(AES_CORE_DATAPATH__abc_15863_new_n5231_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5232_));
NAND2X1 NAND2X1_61 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2827_), .B(AES_CORE_DATAPATH__abc_15863_new_n2825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2828_));
NAND2X1 NAND2X1_610 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5237_));
NAND2X1 NAND2X1_611 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3465_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5240_));
NAND2X1 NAND2X1_612 ( .A(AES_CORE_DATAPATH_col_0__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5244_));
NAND2X1 NAND2X1_613 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3479_), .B(AES_CORE_DATAPATH__abc_15863_new_n2920_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5248_));
NAND2X1 NAND2X1_614 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5257_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5258_));
NAND2X1 NAND2X1_615 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[17] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5263_));
NAND2X1 NAND2X1_616 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5265_), .B(AES_CORE_DATAPATH__abc_15863_new_n5269_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5270_));
NAND2X1 NAND2X1_617 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5275_));
NAND2X1 NAND2X1_618 ( .A(AES_CORE_DATAPATH_col_0__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5283_));
NAND2X1 NAND2X1_619 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3503_), .B(AES_CORE_DATAPATH__abc_15863_new_n2930_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5287_));
NAND2X1 NAND2X1_62 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2838_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2839_));
NAND2X1 NAND2X1_620 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5296_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5297_));
NAND2X1 NAND2X1_621 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[18] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5302_));
NAND2X1 NAND2X1_622 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5304_), .B(AES_CORE_DATAPATH__abc_15863_new_n5308_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5309_));
NAND2X1 NAND2X1_623 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5314_));
NAND2X1 NAND2X1_624 ( .A(AES_CORE_DATAPATH_col_0__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5322_));
NAND2X1 NAND2X1_625 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3523_), .B(AES_CORE_DATAPATH__abc_15863_new_n2940_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5326_));
NAND2X1 NAND2X1_626 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5335_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5336_));
NAND2X1 NAND2X1_627 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[19] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5341_));
NAND2X1 NAND2X1_628 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5343_), .B(AES_CORE_DATAPATH__abc_15863_new_n5347_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5348_));
NAND2X1 NAND2X1_629 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5353_));
NAND2X1 NAND2X1_63 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2839_), .B(AES_CORE_DATAPATH__abc_15863_new_n2837_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2840_));
NAND2X1 NAND2X1_630 ( .A(AES_CORE_DATAPATH_col_0__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5361_));
NAND2X1 NAND2X1_631 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5369_));
NAND2X1 NAND2X1_632 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5373_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5374_));
NAND2X1 NAND2X1_633 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5383_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5384_));
NAND2X1 NAND2X1_634 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[20] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5385_));
NAND2X1 NAND2X1_635 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5381_), .B(AES_CORE_DATAPATH__abc_15863_new_n5387_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5388_));
NAND2X1 NAND2X1_636 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5393_));
NAND2X1 NAND2X1_637 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3553_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5396_));
NAND2X1 NAND2X1_638 ( .A(AES_CORE_DATAPATH_col_0__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5400_));
NAND2X1 NAND2X1_639 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3567_), .B(AES_CORE_DATAPATH__abc_15863_new_n2963_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5404_));
NAND2X1 NAND2X1_64 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2849_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2850_));
NAND2X1 NAND2X1_640 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5413_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5414_));
NAND2X1 NAND2X1_641 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[21] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5419_));
NAND2X1 NAND2X1_642 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5421_), .B(AES_CORE_DATAPATH__abc_15863_new_n5425_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5426_));
NAND2X1 NAND2X1_643 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5431_));
NAND2X1 NAND2X1_644 ( .A(AES_CORE_DATAPATH_col_0__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5439_));
NAND2X1 NAND2X1_645 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5447_));
NAND2X1 NAND2X1_646 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5458_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5459_));
NAND2X1 NAND2X1_647 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[22] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5460_));
NAND2X1 NAND2X1_648 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5456_), .B(AES_CORE_DATAPATH__abc_15863_new_n5462_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5463_));
NAND2X1 NAND2X1_649 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5468_));
NAND2X1 NAND2X1_65 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2850_), .B(AES_CORE_DATAPATH__abc_15863_new_n2848_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2851_));
NAND2X1 NAND2X1_650 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3597_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5471_));
NAND2X1 NAND2X1_651 ( .A(AES_CORE_DATAPATH_col_0__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5475_));
NAND2X1 NAND2X1_652 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5485_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5486_));
NAND2X1 NAND2X1_653 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[23] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5491_));
NAND2X1 NAND2X1_654 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3613_), .B(AES_CORE_DATAPATH__abc_15863_new_n2984_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5495_));
NAND2X1 NAND2X1_655 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5493_), .B(AES_CORE_DATAPATH__abc_15863_new_n5501_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5502_));
NAND2X1 NAND2X1_656 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5507_));
NAND2X1 NAND2X1_657 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3619_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5510_));
NAND2X1 NAND2X1_658 ( .A(AES_CORE_DATAPATH_col_0__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5514_));
NAND2X1 NAND2X1_659 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5522_));
NAND2X1 NAND2X1_66 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2858_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2859_));
NAND2X1 NAND2X1_660 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5526_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5527_));
NAND2X1 NAND2X1_661 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5536_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5537_));
NAND2X1 NAND2X1_662 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[24] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5538_));
NAND2X1 NAND2X1_663 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5534_), .B(AES_CORE_DATAPATH__abc_15863_new_n5540_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5541_));
NAND2X1 NAND2X1_664 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5546_));
NAND2X1 NAND2X1_665 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3641_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5549_));
NAND2X1 NAND2X1_666 ( .A(AES_CORE_DATAPATH_col_0__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5553_));
NAND2X1 NAND2X1_667 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3655_), .B(AES_CORE_DATAPATH__abc_15863_new_n3009_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5557_));
NAND2X1 NAND2X1_668 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5566_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5567_));
NAND2X1 NAND2X1_669 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[25] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5572_));
NAND2X1 NAND2X1_67 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2859_), .B(AES_CORE_DATAPATH__abc_15863_new_n2857_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2860_));
NAND2X1 NAND2X1_670 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5574_), .B(AES_CORE_DATAPATH__abc_15863_new_n5578_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5579_));
NAND2X1 NAND2X1_671 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5584_));
NAND2X1 NAND2X1_672 ( .A(AES_CORE_DATAPATH_col_0__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5592_));
NAND2X1 NAND2X1_673 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3679_), .B(AES_CORE_DATAPATH__abc_15863_new_n3019_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5596_));
NAND2X1 NAND2X1_674 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5605_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5606_));
NAND2X1 NAND2X1_675 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[26] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5611_));
NAND2X1 NAND2X1_676 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5613_), .B(AES_CORE_DATAPATH__abc_15863_new_n5617_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5618_));
NAND2X1 NAND2X1_677 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5623_));
NAND2X1 NAND2X1_678 ( .A(AES_CORE_DATAPATH_col_0__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5631_));
NAND2X1 NAND2X1_679 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5639_));
NAND2X1 NAND2X1_68 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2868_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2869_));
NAND2X1 NAND2X1_680 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5643_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5644_));
NAND2X1 NAND2X1_681 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5653_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5654_));
NAND2X1 NAND2X1_682 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[27] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5655_));
NAND2X1 NAND2X1_683 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5651_), .B(AES_CORE_DATAPATH__abc_15863_new_n5657_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5658_));
NAND2X1 NAND2X1_684 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5663_));
NAND2X1 NAND2X1_685 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3707_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5666_));
NAND2X1 NAND2X1_686 ( .A(AES_CORE_DATAPATH_col_0__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5670_));
NAND2X1 NAND2X1_687 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3721_), .B(AES_CORE_DATAPATH__abc_15863_new_n3040_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5674_));
NAND2X1 NAND2X1_688 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5683_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5684_));
NAND2X1 NAND2X1_689 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[28] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5689_));
NAND2X1 NAND2X1_69 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2869_), .B(AES_CORE_DATAPATH__abc_15863_new_n2867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2870_));
NAND2X1 NAND2X1_690 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5691_), .B(AES_CORE_DATAPATH__abc_15863_new_n5695_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5696_));
NAND2X1 NAND2X1_691 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5701_));
NAND2X1 NAND2X1_692 ( .A(AES_CORE_DATAPATH_col_0__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5709_));
NAND2X1 NAND2X1_693 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5717_));
NAND2X1 NAND2X1_694 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5728_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5729_));
NAND2X1 NAND2X1_695 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[29] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5730_));
NAND2X1 NAND2X1_696 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5726_), .B(AES_CORE_DATAPATH__abc_15863_new_n5732_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5733_));
NAND2X1 NAND2X1_697 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5738_));
NAND2X1 NAND2X1_698 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3751_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5741_));
NAND2X1 NAND2X1_699 ( .A(AES_CORE_DATAPATH_col_0__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5745_));
NAND2X1 NAND2X1_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_));
NAND2X1 NAND2X1_70 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2874_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2875_));
NAND2X1 NAND2X1_700 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5753_));
NAND2X1 NAND2X1_701 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5757_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5758_));
NAND2X1 NAND2X1_702 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5767_), .B(AES_CORE_DATAPATH__abc_15863_new_n4592_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5768_));
NAND2X1 NAND2X1_703 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[30] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5769_));
NAND2X1 NAND2X1_704 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5765_), .B(AES_CORE_DATAPATH__abc_15863_new_n5771_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5772_));
NAND2X1 NAND2X1_705 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5777_));
NAND2X1 NAND2X1_706 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3773_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5780_));
NAND2X1 NAND2X1_707 ( .A(AES_CORE_DATAPATH_col_0__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5784_));
NAND2X1 NAND2X1_708 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3787_), .B(AES_CORE_DATAPATH__abc_15863_new_n3069_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5788_));
NAND2X1 NAND2X1_709 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5797_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5798_));
NAND2X1 NAND2X1_71 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2875_), .B(AES_CORE_DATAPATH__abc_15863_new_n2879_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2880_));
NAND2X1 NAND2X1_710 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(\iv_out[31] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n5803_));
NAND2X1 NAND2X1_711 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5805_), .B(AES_CORE_DATAPATH__abc_15863_new_n5809_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5810_));
NAND2X1 NAND2X1_712 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4626_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5815_));
NAND2X1 NAND2X1_713 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5826_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5827_));
NAND2X1 NAND2X1_714 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5829_));
NAND2X1 NAND2X1_715 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5831_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5832_));
NAND2X1 NAND2X1_716 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5834_));
NAND2X1 NAND2X1_717 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5836_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5837_));
NAND2X1 NAND2X1_718 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5839_));
NAND2X1 NAND2X1_719 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5841_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5842_));
NAND2X1 NAND2X1_72 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2888_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2889_));
NAND2X1 NAND2X1_720 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5844_));
NAND2X1 NAND2X1_721 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5846_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5847_));
NAND2X1 NAND2X1_722 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5849_));
NAND2X1 NAND2X1_723 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5851_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5852_));
NAND2X1 NAND2X1_724 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5854_));
NAND2X1 NAND2X1_725 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5856_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5857_));
NAND2X1 NAND2X1_726 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5859_));
NAND2X1 NAND2X1_727 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5861_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5862_));
NAND2X1 NAND2X1_728 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5864_));
NAND2X1 NAND2X1_729 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5867_));
NAND2X1 NAND2X1_73 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2889_), .B(AES_CORE_DATAPATH__abc_15863_new_n2887_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2890_));
NAND2X1 NAND2X1_730 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5869_));
NAND2X1 NAND2X1_731 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5871_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5872_));
NAND2X1 NAND2X1_732 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5874_));
NAND2X1 NAND2X1_733 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5876_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5877_));
NAND2X1 NAND2X1_734 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5879_));
NAND2X1 NAND2X1_735 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5881_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5882_));
NAND2X1 NAND2X1_736 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5884_));
NAND2X1 NAND2X1_737 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5886_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5887_));
NAND2X1 NAND2X1_738 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5889_));
NAND2X1 NAND2X1_739 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5891_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5892_));
NAND2X1 NAND2X1_74 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2894_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2895_));
NAND2X1 NAND2X1_740 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5894_));
NAND2X1 NAND2X1_741 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5896_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5897_));
NAND2X1 NAND2X1_742 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5899_));
NAND2X1 NAND2X1_743 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5901_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5902_));
NAND2X1 NAND2X1_744 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5904_));
NAND2X1 NAND2X1_745 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5906_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5907_));
NAND2X1 NAND2X1_746 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5909_));
NAND2X1 NAND2X1_747 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5911_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5912_));
NAND2X1 NAND2X1_748 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5914_));
NAND2X1 NAND2X1_749 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5916_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5917_));
NAND2X1 NAND2X1_75 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2895_), .B(AES_CORE_DATAPATH__abc_15863_new_n2899_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2900_));
NAND2X1 NAND2X1_750 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5919_));
NAND2X1 NAND2X1_751 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5921_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5922_));
NAND2X1 NAND2X1_752 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5924_));
NAND2X1 NAND2X1_753 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5926_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5927_));
NAND2X1 NAND2X1_754 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5929_));
NAND2X1 NAND2X1_755 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5931_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5932_));
NAND2X1 NAND2X1_756 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5934_));
NAND2X1 NAND2X1_757 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5936_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5937_));
NAND2X1 NAND2X1_758 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5939_));
NAND2X1 NAND2X1_759 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5941_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5942_));
NAND2X1 NAND2X1_76 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2905_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2906_));
NAND2X1 NAND2X1_760 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5944_));
NAND2X1 NAND2X1_761 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5946_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5947_));
NAND2X1 NAND2X1_762 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5949_));
NAND2X1 NAND2X1_763 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5951_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5952_));
NAND2X1 NAND2X1_764 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5954_));
NAND2X1 NAND2X1_765 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5956_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5957_));
NAND2X1 NAND2X1_766 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5959_));
NAND2X1 NAND2X1_767 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5961_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5962_));
NAND2X1 NAND2X1_768 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5964_));
NAND2X1 NAND2X1_769 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5966_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5967_));
NAND2X1 NAND2X1_77 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2906_), .B(AES_CORE_DATAPATH__abc_15863_new_n2910_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2911_));
NAND2X1 NAND2X1_770 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5969_));
NAND2X1 NAND2X1_771 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5971_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5972_));
NAND2X1 NAND2X1_772 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5974_));
NAND2X1 NAND2X1_773 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5976_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5977_));
NAND2X1 NAND2X1_774 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5979_));
NAND2X1 NAND2X1_775 ( .A(\key_en[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4023_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5981_));
NAND2X1 NAND2X1_776 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3867_), .B(AES_CORE_DATAPATH__abc_15863_new_n5982_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5983_));
NAND2X1 NAND2X1_777 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n5825_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5985_));
NAND2X1 NAND2X1_778 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n5987_));
NAND2X1 NAND2X1_779 ( .A(AES_CORE_DATAPATH_col_3__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6051_));
NAND2X1 NAND2X1_78 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2914_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2915_));
NAND2X1 NAND2X1_780 ( .A(AES_CORE_DATAPATH_col_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6058_));
NAND2X1 NAND2X1_781 ( .A(AES_CORE_DATAPATH_col_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6065_));
NAND2X1 NAND2X1_782 ( .A(AES_CORE_DATAPATH_col_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6072_));
NAND2X1 NAND2X1_783 ( .A(AES_CORE_DATAPATH_col_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6079_));
NAND2X1 NAND2X1_784 ( .A(AES_CORE_DATAPATH_col_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6086_));
NAND2X1 NAND2X1_785 ( .A(AES_CORE_DATAPATH_col_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6093_));
NAND2X1 NAND2X1_786 ( .A(AES_CORE_DATAPATH_col_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6100_));
NAND2X1 NAND2X1_787 ( .A(AES_CORE_DATAPATH_col_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6107_));
NAND2X1 NAND2X1_788 ( .A(AES_CORE_DATAPATH_col_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6114_));
NAND2X1 NAND2X1_789 ( .A(AES_CORE_DATAPATH_col_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6121_));
NAND2X1 NAND2X1_79 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2915_), .B(AES_CORE_DATAPATH__abc_15863_new_n2919_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2920_));
NAND2X1 NAND2X1_790 ( .A(AES_CORE_DATAPATH_col_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6128_));
NAND2X1 NAND2X1_791 ( .A(AES_CORE_DATAPATH_col_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6135_));
NAND2X1 NAND2X1_792 ( .A(AES_CORE_DATAPATH_col_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6142_));
NAND2X1 NAND2X1_793 ( .A(AES_CORE_DATAPATH_col_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6149_));
NAND2X1 NAND2X1_794 ( .A(AES_CORE_DATAPATH_col_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6156_));
NAND2X1 NAND2X1_795 ( .A(AES_CORE_DATAPATH_col_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6163_));
NAND2X1 NAND2X1_796 ( .A(AES_CORE_DATAPATH_col_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6170_));
NAND2X1 NAND2X1_797 ( .A(AES_CORE_DATAPATH_col_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6177_));
NAND2X1 NAND2X1_798 ( .A(AES_CORE_DATAPATH_col_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6184_));
NAND2X1 NAND2X1_799 ( .A(AES_CORE_DATAPATH_col_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6191_));
NAND2X1 NAND2X1_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n124_), .Y(AES_CORE_CONTROL_UNIT_bypass_rk));
NAND2X1 NAND2X1_80 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2924_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2925_));
NAND2X1 NAND2X1_800 ( .A(AES_CORE_DATAPATH_col_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6198_));
NAND2X1 NAND2X1_801 ( .A(AES_CORE_DATAPATH_col_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6205_));
NAND2X1 NAND2X1_802 ( .A(AES_CORE_DATAPATH_col_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6212_));
NAND2X1 NAND2X1_803 ( .A(AES_CORE_DATAPATH_col_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6219_));
NAND2X1 NAND2X1_804 ( .A(AES_CORE_DATAPATH_col_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6226_));
NAND2X1 NAND2X1_805 ( .A(AES_CORE_DATAPATH_col_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6233_));
NAND2X1 NAND2X1_806 ( .A(AES_CORE_DATAPATH_col_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6240_));
NAND2X1 NAND2X1_807 ( .A(AES_CORE_DATAPATH_col_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6247_));
NAND2X1 NAND2X1_808 ( .A(AES_CORE_DATAPATH_col_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6254_));
NAND2X1 NAND2X1_809 ( .A(AES_CORE_DATAPATH_col_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6261_));
NAND2X1 NAND2X1_81 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2925_), .B(AES_CORE_DATAPATH__abc_15863_new_n2929_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2930_));
NAND2X1 NAND2X1_810 ( .A(AES_CORE_DATAPATH_col_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n2461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6268_));
NAND2X1 NAND2X1_811 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6275_));
NAND2X1 NAND2X1_812 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6282_));
NAND2X1 NAND2X1_813 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6289_));
NAND2X1 NAND2X1_814 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6296_));
NAND2X1 NAND2X1_815 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6303_));
NAND2X1 NAND2X1_816 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6310_));
NAND2X1 NAND2X1_817 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6317_));
NAND2X1 NAND2X1_818 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6324_));
NAND2X1 NAND2X1_819 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6331_));
NAND2X1 NAND2X1_82 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2934_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2935_));
NAND2X1 NAND2X1_820 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6338_));
NAND2X1 NAND2X1_821 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6345_));
NAND2X1 NAND2X1_822 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6352_));
NAND2X1 NAND2X1_823 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6359_));
NAND2X1 NAND2X1_824 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6366_));
NAND2X1 NAND2X1_825 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6373_));
NAND2X1 NAND2X1_826 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6380_));
NAND2X1 NAND2X1_827 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6387_));
NAND2X1 NAND2X1_828 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6394_));
NAND2X1 NAND2X1_829 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6401_));
NAND2X1 NAND2X1_83 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2935_), .B(AES_CORE_DATAPATH__abc_15863_new_n2939_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2940_));
NAND2X1 NAND2X1_830 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6408_));
NAND2X1 NAND2X1_831 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6415_));
NAND2X1 NAND2X1_832 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6422_));
NAND2X1 NAND2X1_833 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6429_));
NAND2X1 NAND2X1_834 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6436_));
NAND2X1 NAND2X1_835 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6443_));
NAND2X1 NAND2X1_836 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6450_));
NAND2X1 NAND2X1_837 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6457_));
NAND2X1 NAND2X1_838 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6464_));
NAND2X1 NAND2X1_839 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6471_));
NAND2X1 NAND2X1_84 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2945_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2946_));
NAND2X1 NAND2X1_840 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6478_));
NAND2X1 NAND2X1_841 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6485_));
NAND2X1 NAND2X1_842 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .B(AES_CORE_DATAPATH__abc_15863_new_n2474_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6492_));
NAND2X1 NAND2X1_843 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6500_));
NAND2X1 NAND2X1_844 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6510_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6511_));
NAND2X1 NAND2X1_845 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6513_));
NAND2X1 NAND2X1_846 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6523_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6524_));
NAND2X1 NAND2X1_847 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6526_));
NAND2X1 NAND2X1_848 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6533_));
NAND2X1 NAND2X1_849 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6540_));
NAND2X1 NAND2X1_85 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2946_), .B(AES_CORE_DATAPATH__abc_15863_new_n2950_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2951_));
NAND2X1 NAND2X1_850 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6550_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6551_));
NAND2X1 NAND2X1_851 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6553_));
NAND2X1 NAND2X1_852 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6564_));
NAND2X1 NAND2X1_853 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6566_));
NAND2X1 NAND2X1_854 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6576_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6577_));
NAND2X1 NAND2X1_855 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6579_));
NAND2X1 NAND2X1_856 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6589_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6590_));
NAND2X1 NAND2X1_857 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6592_));
NAND2X1 NAND2X1_858 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6602_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6603_));
NAND2X1 NAND2X1_859 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6605_));
NAND2X1 NAND2X1_86 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2957_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2958_));
NAND2X1 NAND2X1_860 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6615_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6616_));
NAND2X1 NAND2X1_861 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6621_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6622_));
NAND2X1 NAND2X1_862 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6627_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6628_));
NAND2X1 NAND2X1_863 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6630_));
NAND2X1 NAND2X1_864 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6640_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6641_));
NAND2X1 NAND2X1_865 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6643_));
NAND2X1 NAND2X1_866 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6653_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6654_));
NAND2X1 NAND2X1_867 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6656_));
NAND2X1 NAND2X1_868 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6666_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6667_));
NAND2X1 NAND2X1_869 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6672_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6673_));
NAND2X1 NAND2X1_87 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2958_), .B(AES_CORE_DATAPATH__abc_15863_new_n2962_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2963_));
NAND2X1 NAND2X1_870 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6675_));
NAND2X1 NAND2X1_871 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6685_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6686_));
NAND2X1 NAND2X1_872 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6688_));
NAND2X1 NAND2X1_873 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .B(AES_CORE_DATAPATH__abc_15863_new_n6499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6695_));
NAND2X1 NAND2X1_874 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2466_), .B(AES_CORE_DATAPATH__abc_15863_new_n6705_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6706_));
NAND2X1 NAND2X1_875 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_DATAPATH__abc_15863_new_n6710_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6711_));
NAND2X1 NAND2X1_876 ( .A(AES_CORE_DATAPATH_bkp_1_3__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6714_));
NAND2X1 NAND2X1_877 ( .A(AES_CORE_DATAPATH_bkp_1_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6716_));
NAND2X1 NAND2X1_878 ( .A(AES_CORE_DATAPATH_bkp_1_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6718_));
NAND2X1 NAND2X1_879 ( .A(AES_CORE_DATAPATH_bkp_1_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6720_));
NAND2X1 NAND2X1_88 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2967_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2968_));
NAND2X1 NAND2X1_880 ( .A(AES_CORE_DATAPATH_bkp_1_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6722_));
NAND2X1 NAND2X1_881 ( .A(AES_CORE_DATAPATH_bkp_1_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6724_));
NAND2X1 NAND2X1_882 ( .A(AES_CORE_DATAPATH_bkp_1_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6726_));
NAND2X1 NAND2X1_883 ( .A(AES_CORE_DATAPATH_bkp_1_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6728_));
NAND2X1 NAND2X1_884 ( .A(AES_CORE_DATAPATH_bkp_1_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6730_));
NAND2X1 NAND2X1_885 ( .A(AES_CORE_DATAPATH_bkp_1_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6732_));
NAND2X1 NAND2X1_886 ( .A(AES_CORE_DATAPATH_bkp_1_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6734_));
NAND2X1 NAND2X1_887 ( .A(AES_CORE_DATAPATH_bkp_1_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6736_));
NAND2X1 NAND2X1_888 ( .A(AES_CORE_DATAPATH_bkp_1_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6738_));
NAND2X1 NAND2X1_889 ( .A(AES_CORE_DATAPATH_bkp_1_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6740_));
NAND2X1 NAND2X1_89 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2968_), .B(AES_CORE_DATAPATH__abc_15863_new_n2972_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2973_));
NAND2X1 NAND2X1_890 ( .A(AES_CORE_DATAPATH_bkp_1_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6742_));
NAND2X1 NAND2X1_891 ( .A(AES_CORE_DATAPATH_bkp_1_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6744_));
NAND2X1 NAND2X1_892 ( .A(AES_CORE_DATAPATH_bkp_1_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6746_));
NAND2X1 NAND2X1_893 ( .A(AES_CORE_DATAPATH_bkp_1_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6748_));
NAND2X1 NAND2X1_894 ( .A(AES_CORE_DATAPATH_bkp_1_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6750_));
NAND2X1 NAND2X1_895 ( .A(AES_CORE_DATAPATH_bkp_1_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6752_));
NAND2X1 NAND2X1_896 ( .A(AES_CORE_DATAPATH_bkp_1_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6754_));
NAND2X1 NAND2X1_897 ( .A(AES_CORE_DATAPATH_bkp_1_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6756_));
NAND2X1 NAND2X1_898 ( .A(AES_CORE_DATAPATH_bkp_1_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6758_));
NAND2X1 NAND2X1_899 ( .A(AES_CORE_DATAPATH_bkp_1_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6760_));
NAND2X1 NAND2X1_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n78_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n133_));
NAND2X1 NAND2X1_90 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2978_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2979_));
NAND2X1 NAND2X1_900 ( .A(AES_CORE_DATAPATH_bkp_1_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6762_));
NAND2X1 NAND2X1_901 ( .A(AES_CORE_DATAPATH_bkp_1_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6764_));
NAND2X1 NAND2X1_902 ( .A(AES_CORE_DATAPATH_bkp_1_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6766_));
NAND2X1 NAND2X1_903 ( .A(AES_CORE_DATAPATH_bkp_1_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6768_));
NAND2X1 NAND2X1_904 ( .A(AES_CORE_DATAPATH_bkp_1_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6770_));
NAND2X1 NAND2X1_905 ( .A(AES_CORE_DATAPATH_bkp_1_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6772_));
NAND2X1 NAND2X1_906 ( .A(AES_CORE_DATAPATH_bkp_1_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6774_));
NAND2X1 NAND2X1_907 ( .A(AES_CORE_DATAPATH_bkp_1_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6776_));
NAND2X1 NAND2X1_908 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4236_), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6985_));
NAND2X1 NAND2X1_909 ( .A(AES_CORE_DATAPATH_iv_3__0_), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6986_));
NAND2X1 NAND2X1_91 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2979_), .B(AES_CORE_DATAPATH__abc_15863_new_n2983_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2984_));
NAND2X1 NAND2X1_910 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n6987_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6988_));
NAND2X1 NAND2X1_911 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(AES_CORE_DATAPATH__abc_15863_new_n6995_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6996_));
NAND2X1 NAND2X1_912 ( .A(AES_CORE_DATAPATH_iv_3__2_), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7000_));
NAND2X1 NAND2X1_913 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(AES_CORE_DATAPATH__abc_15863_new_n7003_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7004_));
NAND2X1 NAND2X1_914 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(AES_CORE_DATAPATH__abc_15863_new_n7009_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7010_));
NAND2X1 NAND2X1_915 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7014_), .B(AES_CORE_DATAPATH__abc_15863_new_n7001_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7026_));
NAND2X1 NAND2X1_916 ( .A(AES_CORE_DATAPATH_iv_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n7027_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7028_));
NAND2X1 NAND2X1_917 ( .A(AES_CORE_DATAPATH_iv_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7040_));
NAND2X1 NAND2X1_918 ( .A(AES_CORE_DATAPATH_iv_3__8_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7041_));
NAND2X1 NAND2X1_919 ( .A(AES_CORE_DATAPATH_iv_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7047_));
NAND2X1 NAND2X1_92 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2995_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2996_));
NAND2X1 NAND2X1_920 ( .A(AES_CORE_DATAPATH_iv_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n7042_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7048_));
NAND2X1 NAND2X1_921 ( .A(AES_CORE_DATAPATH_iv_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n7039_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7054_));
NAND2X1 NAND2X1_922 ( .A(AES_CORE_DATAPATH_iv_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n7055_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7060_));
NAND2X1 NAND2X1_923 ( .A(AES_CORE_DATAPATH_iv_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n7078_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7084_));
NAND2X1 NAND2X1_924 ( .A(AES_CORE_DATAPATH_iv_3__10_), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7107_));
NAND2X1 NAND2X1_925 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7115_), .B(AES_CORE_DATAPATH__abc_15863_new_n7112_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7117_));
NAND2X1 NAND2X1_926 ( .A(AES_CORE_DATAPATH_iv_3__20_), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7130_));
NAND2X1 NAND2X1_927 ( .A(AES_CORE_DATAPATH_iv_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n7131_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7139_));
NAND2X1 NAND2X1_928 ( .A(AES_CORE_DATAPATH_iv_3__22_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7145_));
NAND2X1 NAND2X1_929 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7147_), .B(AES_CORE_DATAPATH__abc_15863_new_n7112_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7148_));
NAND2X1 NAND2X1_93 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2996_), .B(AES_CORE_DATAPATH__abc_15863_new_n2994_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2997_));
NAND2X1 NAND2X1_930 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7163_), .B(AES_CORE_DATAPATH__abc_15863_new_n7149_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7164_));
NAND2X1 NAND2X1_931 ( .A(AES_CORE_DATAPATH_iv_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n7165_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7173_));
NAND2X1 NAND2X1_932 ( .A(AES_CORE_DATAPATH_iv_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n7180_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7189_));
NAND2X1 NAND2X1_933 ( .A(AES_CORE_DATAPATH_iv_3__28_), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7195_));
NAND2X1 NAND2X1_934 ( .A(AES_CORE_DATAPATH_iv_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n7196_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7204_));
NAND2X1 NAND2X1_935 ( .A(\bus_in[0] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7210_));
NAND2X1 NAND2X1_936 ( .A(\bus_in[1] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7212_));
NAND2X1 NAND2X1_937 ( .A(\bus_in[3] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7216_));
NAND2X1 NAND2X1_938 ( .A(\bus_in[6] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7222_));
NAND2X1 NAND2X1_939 ( .A(\bus_in[7] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7224_));
NAND2X1 NAND2X1_94 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3007_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3008_));
NAND2X1 NAND2X1_940 ( .A(\bus_in[8] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7226_));
NAND2X1 NAND2X1_941 ( .A(\bus_in[9] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7228_));
NAND2X1 NAND2X1_942 ( .A(\bus_in[10] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7230_));
NAND2X1 NAND2X1_943 ( .A(\bus_in[11] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7232_));
NAND2X1 NAND2X1_944 ( .A(\bus_in[13] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7236_));
NAND2X1 NAND2X1_945 ( .A(\bus_in[15] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7240_));
NAND2X1 NAND2X1_946 ( .A(\bus_in[17] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7244_));
NAND2X1 NAND2X1_947 ( .A(\bus_in[18] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7246_));
NAND2X1 NAND2X1_948 ( .A(\bus_in[19] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7248_));
NAND2X1 NAND2X1_949 ( .A(\bus_in[21] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7252_));
NAND2X1 NAND2X1_95 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3008_), .B(AES_CORE_DATAPATH__abc_15863_new_n3006_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3009_));
NAND2X1 NAND2X1_950 ( .A(\bus_in[23] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7256_));
NAND2X1 NAND2X1_951 ( .A(\bus_in[25] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7260_));
NAND2X1 NAND2X1_952 ( .A(\bus_in[26] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7262_));
NAND2X1 NAND2X1_953 ( .A(\bus_in[28] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7266_));
NAND2X1 NAND2X1_954 ( .A(\bus_in[31] ), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7272_));
NAND2X1 NAND2X1_955 ( .A(AES_CORE_DATAPATH_bkp_1_2__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7275_));
NAND2X1 NAND2X1_956 ( .A(AES_CORE_DATAPATH_bkp_1_2__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7277_));
NAND2X1 NAND2X1_957 ( .A(AES_CORE_DATAPATH_bkp_1_2__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7279_));
NAND2X1 NAND2X1_958 ( .A(AES_CORE_DATAPATH_bkp_1_2__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7281_));
NAND2X1 NAND2X1_959 ( .A(AES_CORE_DATAPATH_bkp_1_2__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7283_));
NAND2X1 NAND2X1_96 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3017_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3018_));
NAND2X1 NAND2X1_960 ( .A(AES_CORE_DATAPATH_bkp_1_2__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7285_));
NAND2X1 NAND2X1_961 ( .A(AES_CORE_DATAPATH_bkp_1_2__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7287_));
NAND2X1 NAND2X1_962 ( .A(AES_CORE_DATAPATH_bkp_1_2__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7289_));
NAND2X1 NAND2X1_963 ( .A(AES_CORE_DATAPATH_bkp_1_2__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7291_));
NAND2X1 NAND2X1_964 ( .A(AES_CORE_DATAPATH_bkp_1_2__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7293_));
NAND2X1 NAND2X1_965 ( .A(AES_CORE_DATAPATH_bkp_1_2__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7295_));
NAND2X1 NAND2X1_966 ( .A(AES_CORE_DATAPATH_bkp_1_2__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7297_));
NAND2X1 NAND2X1_967 ( .A(AES_CORE_DATAPATH_bkp_1_2__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7299_));
NAND2X1 NAND2X1_968 ( .A(AES_CORE_DATAPATH_bkp_1_2__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7301_));
NAND2X1 NAND2X1_969 ( .A(AES_CORE_DATAPATH_bkp_1_2__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7303_));
NAND2X1 NAND2X1_97 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3018_), .B(AES_CORE_DATAPATH__abc_15863_new_n3016_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3019_));
NAND2X1 NAND2X1_970 ( .A(AES_CORE_DATAPATH_bkp_1_2__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7305_));
NAND2X1 NAND2X1_971 ( .A(AES_CORE_DATAPATH_bkp_1_2__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7307_));
NAND2X1 NAND2X1_972 ( .A(AES_CORE_DATAPATH_bkp_1_2__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7309_));
NAND2X1 NAND2X1_973 ( .A(AES_CORE_DATAPATH_bkp_1_2__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7311_));
NAND2X1 NAND2X1_974 ( .A(AES_CORE_DATAPATH_bkp_1_2__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7313_));
NAND2X1 NAND2X1_975 ( .A(AES_CORE_DATAPATH_bkp_1_2__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7315_));
NAND2X1 NAND2X1_976 ( .A(AES_CORE_DATAPATH_bkp_1_2__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7317_));
NAND2X1 NAND2X1_977 ( .A(AES_CORE_DATAPATH_bkp_1_2__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7319_));
NAND2X1 NAND2X1_978 ( .A(AES_CORE_DATAPATH_bkp_1_2__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7321_));
NAND2X1 NAND2X1_979 ( .A(AES_CORE_DATAPATH_bkp_1_2__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7323_));
NAND2X1 NAND2X1_98 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3027_), .B(AES_CORE_DATAPATH__abc_15863_new_n2729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3028_));
NAND2X1 NAND2X1_980 ( .A(AES_CORE_DATAPATH_bkp_1_2__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7325_));
NAND2X1 NAND2X1_981 ( .A(AES_CORE_DATAPATH_bkp_1_2__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7327_));
NAND2X1 NAND2X1_982 ( .A(AES_CORE_DATAPATH_bkp_1_2__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7329_));
NAND2X1 NAND2X1_983 ( .A(AES_CORE_DATAPATH_bkp_1_2__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7331_));
NAND2X1 NAND2X1_984 ( .A(AES_CORE_DATAPATH_bkp_1_2__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7333_));
NAND2X1 NAND2X1_985 ( .A(AES_CORE_DATAPATH_bkp_1_2__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7335_));
NAND2X1 NAND2X1_986 ( .A(AES_CORE_DATAPATH_bkp_1_2__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7337_));
NAND2X1 NAND2X1_987 ( .A(\bus_in[0] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7499_));
NAND2X1 NAND2X1_988 ( .A(\bus_in[6] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7511_));
NAND2X1 NAND2X1_989 ( .A(\bus_in[7] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7513_));
NAND2X1 NAND2X1_99 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3028_), .B(AES_CORE_DATAPATH__abc_15863_new_n3026_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3029_));
NAND2X1 NAND2X1_990 ( .A(\bus_in[8] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7515_));
NAND2X1 NAND2X1_991 ( .A(\bus_in[9] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7517_));
NAND2X1 NAND2X1_992 ( .A(\bus_in[10] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7519_));
NAND2X1 NAND2X1_993 ( .A(\bus_in[11] ), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7521_));
NAND2X1 NAND2X1_994 ( .A(AES_CORE_DATAPATH_bkp_1_1__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7564_));
NAND2X1 NAND2X1_995 ( .A(AES_CORE_DATAPATH_bkp_1_1__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7569_));
NAND2X1 NAND2X1_996 ( .A(AES_CORE_DATAPATH_bkp_1_1__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7574_));
NAND2X1 NAND2X1_997 ( .A(AES_CORE_DATAPATH_bkp_1_1__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7576_));
NAND2X1 NAND2X1_998 ( .A(AES_CORE_DATAPATH_bkp_1_1__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7578_));
NAND2X1 NAND2X1_999 ( .A(AES_CORE_DATAPATH_bkp_1_1__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7583_));
NAND3X1 NAND3X1_1 ( .A(\addr[1] ), .B(\addr[0] ), .C(write_en), .Y(_abc_15574_new_n17_));
NAND3X1 NAND3X1_10 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n2717_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2718_));
NAND3X1 NAND3X1_100 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3034_), .B(AES_CORE_DATAPATH__abc_15863_new_n3035_), .C(AES_CORE_DATAPATH__abc_15863_new_n3036_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3037_));
NAND3X1 NAND3X1_1000 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n91_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n92_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n93_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_));
NAND3X1 NAND3X1_1001 ( .A(\data_type[0] ), .B(\bus_in[22] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n95_));
NAND3X1 NAND3X1_1002 ( .A(\data_type[1] ), .B(\bus_in[30] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n96_));
NAND3X1 NAND3X1_1003 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n95_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n96_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n97_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_));
NAND3X1 NAND3X1_1004 ( .A(\data_type[0] ), .B(\bus_in[23] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n99_));
NAND3X1 NAND3X1_1005 ( .A(\data_type[1] ), .B(\bus_in[31] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n100_));
NAND3X1 NAND3X1_1006 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n99_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n100_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n101_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_));
NAND3X1 NAND3X1_1007 ( .A(\data_type[0] ), .B(\bus_in[24] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n103_));
NAND3X1 NAND3X1_1008 ( .A(\data_type[1] ), .B(\bus_in[16] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n104_));
NAND3X1 NAND3X1_1009 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n103_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n104_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n105_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_));
NAND3X1 NAND3X1_101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3044_));
NAND3X1 NAND3X1_1010 ( .A(\data_type[0] ), .B(\bus_in[25] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n107_));
NAND3X1 NAND3X1_1011 ( .A(\data_type[1] ), .B(\bus_in[17] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n108_));
NAND3X1 NAND3X1_1012 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n107_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n108_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n109_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_));
NAND3X1 NAND3X1_1013 ( .A(\data_type[0] ), .B(\bus_in[26] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n111_));
NAND3X1 NAND3X1_1014 ( .A(\data_type[1] ), .B(\bus_in[18] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n112_));
NAND3X1 NAND3X1_1015 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n111_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n112_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n113_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_));
NAND3X1 NAND3X1_1016 ( .A(\data_type[0] ), .B(\bus_in[27] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n115_));
NAND3X1 NAND3X1_1017 ( .A(\data_type[1] ), .B(\bus_in[19] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n116_));
NAND3X1 NAND3X1_1018 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n115_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n116_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n117_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_));
NAND3X1 NAND3X1_1019 ( .A(\data_type[0] ), .B(\bus_in[28] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n119_));
NAND3X1 NAND3X1_102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3045_));
NAND3X1 NAND3X1_1020 ( .A(\data_type[1] ), .B(\bus_in[20] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n120_));
NAND3X1 NAND3X1_1021 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n119_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n120_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n121_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_));
NAND3X1 NAND3X1_1022 ( .A(\data_type[0] ), .B(\bus_in[29] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n123_));
NAND3X1 NAND3X1_1023 ( .A(\data_type[1] ), .B(\bus_in[21] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n124_));
NAND3X1 NAND3X1_1024 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n123_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n124_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n125_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_));
NAND3X1 NAND3X1_1025 ( .A(\data_type[0] ), .B(\bus_in[30] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n127_));
NAND3X1 NAND3X1_1026 ( .A(\data_type[1] ), .B(\bus_in[22] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n128_));
NAND3X1 NAND3X1_1027 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n127_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n128_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n129_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_));
NAND3X1 NAND3X1_1028 ( .A(\data_type[0] ), .B(\bus_in[31] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n131_));
NAND3X1 NAND3X1_1029 ( .A(\data_type[1] ), .B(\bus_in[23] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n132_));
NAND3X1 NAND3X1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3044_), .B(AES_CORE_DATAPATH__abc_15863_new_n3045_), .C(AES_CORE_DATAPATH__abc_15863_new_n3046_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3047_));
NAND3X1 NAND3X1_1030 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n131_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n132_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n133_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_));
NAND3X1 NAND3X1_1031 ( .A(\data_type[0] ), .B(\bus_in[0] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n135_));
NAND3X1 NAND3X1_1032 ( .A(\data_type[1] ), .B(\bus_in[8] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n136_));
NAND3X1 NAND3X1_1033 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n135_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n136_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n137_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_));
NAND3X1 NAND3X1_1034 ( .A(\data_type[0] ), .B(\bus_in[1] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n139_));
NAND3X1 NAND3X1_1035 ( .A(\data_type[1] ), .B(\bus_in[9] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n140_));
NAND3X1 NAND3X1_1036 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n139_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n140_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n141_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_));
NAND3X1 NAND3X1_1037 ( .A(\data_type[0] ), .B(\bus_in[2] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n143_));
NAND3X1 NAND3X1_1038 ( .A(\data_type[1] ), .B(\bus_in[10] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n144_));
NAND3X1 NAND3X1_1039 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n143_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n144_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n145_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_));
NAND3X1 NAND3X1_104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3054_));
NAND3X1 NAND3X1_1040 ( .A(\data_type[0] ), .B(\bus_in[3] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n147_));
NAND3X1 NAND3X1_1041 ( .A(\data_type[1] ), .B(\bus_in[11] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n148_));
NAND3X1 NAND3X1_1042 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n147_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n148_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n149_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_));
NAND3X1 NAND3X1_1043 ( .A(\data_type[0] ), .B(\bus_in[4] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n151_));
NAND3X1 NAND3X1_1044 ( .A(\data_type[1] ), .B(\bus_in[12] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n152_));
NAND3X1 NAND3X1_1045 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n151_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n152_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n153_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_));
NAND3X1 NAND3X1_1046 ( .A(\data_type[0] ), .B(\bus_in[5] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n155_));
NAND3X1 NAND3X1_1047 ( .A(\data_type[1] ), .B(\bus_in[13] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n156_));
NAND3X1 NAND3X1_1048 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n155_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n156_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n157_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_));
NAND3X1 NAND3X1_1049 ( .A(\data_type[0] ), .B(\bus_in[6] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n159_));
NAND3X1 NAND3X1_105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3055_));
NAND3X1 NAND3X1_1050 ( .A(\data_type[1] ), .B(\bus_in[14] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n160_));
NAND3X1 NAND3X1_1051 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n159_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n160_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n161_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_));
NAND3X1 NAND3X1_1052 ( .A(\data_type[0] ), .B(\bus_in[7] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n163_));
NAND3X1 NAND3X1_1053 ( .A(\data_type[1] ), .B(\bus_in[15] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n164_));
NAND3X1 NAND3X1_1054 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n163_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n164_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n165_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_));
NAND3X1 NAND3X1_1055 ( .A(\data_type[0] ), .B(\bus_in[8] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n167_));
NAND3X1 NAND3X1_1056 ( .A(\data_type[1] ), .B(\bus_in[0] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n168_));
NAND3X1 NAND3X1_1057 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n167_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n168_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n169_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_));
NAND3X1 NAND3X1_1058 ( .A(\data_type[0] ), .B(\bus_in[9] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n171_));
NAND3X1 NAND3X1_1059 ( .A(\data_type[1] ), .B(\bus_in[1] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n172_));
NAND3X1 NAND3X1_106 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3054_), .B(AES_CORE_DATAPATH__abc_15863_new_n3055_), .C(AES_CORE_DATAPATH__abc_15863_new_n3056_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3057_));
NAND3X1 NAND3X1_1060 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n171_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n172_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n173_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_));
NAND3X1 NAND3X1_1061 ( .A(\data_type[0] ), .B(\bus_in[10] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n175_));
NAND3X1 NAND3X1_1062 ( .A(\data_type[1] ), .B(\bus_in[2] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n176_));
NAND3X1 NAND3X1_1063 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n175_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n176_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n177_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_));
NAND3X1 NAND3X1_1064 ( .A(\data_type[0] ), .B(\bus_in[11] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n179_));
NAND3X1 NAND3X1_1065 ( .A(\data_type[1] ), .B(\bus_in[3] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n180_));
NAND3X1 NAND3X1_1066 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n179_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n180_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n181_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_));
NAND3X1 NAND3X1_1067 ( .A(\data_type[0] ), .B(\bus_in[12] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n183_));
NAND3X1 NAND3X1_1068 ( .A(\data_type[1] ), .B(\bus_in[4] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n184_));
NAND3X1 NAND3X1_1069 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n183_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n184_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n185_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_));
NAND3X1 NAND3X1_107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3065_));
NAND3X1 NAND3X1_1070 ( .A(\data_type[0] ), .B(\bus_in[13] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n187_));
NAND3X1 NAND3X1_1071 ( .A(\data_type[1] ), .B(\bus_in[5] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n188_));
NAND3X1 NAND3X1_1072 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n187_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n188_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n189_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_));
NAND3X1 NAND3X1_1073 ( .A(\data_type[0] ), .B(\bus_in[14] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n191_));
NAND3X1 NAND3X1_1074 ( .A(\data_type[1] ), .B(\bus_in[6] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n192_));
NAND3X1 NAND3X1_1075 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n191_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n192_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n193_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_));
NAND3X1 NAND3X1_1076 ( .A(\data_type[0] ), .B(\bus_in[15] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n195_));
NAND3X1 NAND3X1_1077 ( .A(\data_type[1] ), .B(\bus_in[7] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n196_));
NAND3X1 NAND3X1_1078 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n195_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n196_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n197_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_));
NAND3X1 NAND3X1_1079 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n68_));
NAND3X1 NAND3X1_108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3066_));
NAND3X1 NAND3X1_1080 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n70_));
NAND3X1 NAND3X1_1081 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n68_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n70_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n73_), .Y(\col_out[0] ));
NAND3X1 NAND3X1_1082 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n75_));
NAND3X1 NAND3X1_1083 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n76_));
NAND3X1 NAND3X1_1084 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n75_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n76_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n77_), .Y(\col_out[1] ));
NAND3X1 NAND3X1_1085 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n79_));
NAND3X1 NAND3X1_1086 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n80_));
NAND3X1 NAND3X1_1087 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n79_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n80_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n81_), .Y(\col_out[2] ));
NAND3X1 NAND3X1_1088 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n83_));
NAND3X1 NAND3X1_1089 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n84_));
NAND3X1 NAND3X1_109 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3065_), .B(AES_CORE_DATAPATH__abc_15863_new_n3066_), .C(AES_CORE_DATAPATH__abc_15863_new_n3067_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3068_));
NAND3X1 NAND3X1_1090 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n83_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n84_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n85_), .Y(\col_out[3] ));
NAND3X1 NAND3X1_1091 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n87_));
NAND3X1 NAND3X1_1092 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n88_));
NAND3X1 NAND3X1_1093 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n87_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n88_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n89_), .Y(\col_out[4] ));
NAND3X1 NAND3X1_1094 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n91_));
NAND3X1 NAND3X1_1095 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n92_));
NAND3X1 NAND3X1_1096 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n91_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n92_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n93_), .Y(\col_out[5] ));
NAND3X1 NAND3X1_1097 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n95_));
NAND3X1 NAND3X1_1098 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n96_));
NAND3X1 NAND3X1_1099 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n95_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n96_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n97_), .Y(\col_out[6] ));
NAND3X1 NAND3X1_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2712_), .B(AES_CORE_DATAPATH__abc_15863_new_n2714_), .C(AES_CORE_DATAPATH__abc_15863_new_n2718_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2719_));
NAND3X1 NAND3X1_110 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3088_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3089_));
NAND3X1 NAND3X1_1100 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n99_));
NAND3X1 NAND3X1_1101 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n100_));
NAND3X1 NAND3X1_1102 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n99_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n100_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n101_), .Y(\col_out[7] ));
NAND3X1 NAND3X1_1103 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n103_));
NAND3X1 NAND3X1_1104 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n104_));
NAND3X1 NAND3X1_1105 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n103_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n104_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n105_), .Y(\col_out[8] ));
NAND3X1 NAND3X1_1106 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n107_));
NAND3X1 NAND3X1_1107 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n108_));
NAND3X1 NAND3X1_1108 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n107_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n108_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n109_), .Y(\col_out[9] ));
NAND3X1 NAND3X1_1109 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n111_));
NAND3X1 NAND3X1_111 ( .A(AES_CORE_DATAPATH_col_0__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3092_));
NAND3X1 NAND3X1_1110 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n112_));
NAND3X1 NAND3X1_1111 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n111_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n112_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n113_), .Y(\col_out[10] ));
NAND3X1 NAND3X1_1112 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n115_));
NAND3X1 NAND3X1_1113 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n116_));
NAND3X1 NAND3X1_1114 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n115_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n116_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n117_), .Y(\col_out[11] ));
NAND3X1 NAND3X1_1115 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n119_));
NAND3X1 NAND3X1_1116 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n120_));
NAND3X1 NAND3X1_1117 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n119_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n120_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n121_), .Y(\col_out[12] ));
NAND3X1 NAND3X1_1118 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n123_));
NAND3X1 NAND3X1_1119 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n124_));
NAND3X1 NAND3X1_112 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3093_));
NAND3X1 NAND3X1_1120 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n123_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n124_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n125_), .Y(\col_out[13] ));
NAND3X1 NAND3X1_1121 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n127_));
NAND3X1 NAND3X1_1122 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n128_));
NAND3X1 NAND3X1_1123 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n127_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n128_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n129_), .Y(\col_out[14] ));
NAND3X1 NAND3X1_1124 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n131_));
NAND3X1 NAND3X1_1125 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n132_));
NAND3X1 NAND3X1_1126 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n131_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n132_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n133_), .Y(\col_out[15] ));
NAND3X1 NAND3X1_1127 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n135_));
NAND3X1 NAND3X1_1128 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n136_));
NAND3X1 NAND3X1_1129 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n135_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n136_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n137_), .Y(\col_out[16] ));
NAND3X1 NAND3X1_113 ( .A(AES_CORE_DATAPATH_col_3__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3095_));
NAND3X1 NAND3X1_1130 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n139_));
NAND3X1 NAND3X1_1131 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n140_));
NAND3X1 NAND3X1_1132 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n139_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n140_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n141_), .Y(\col_out[17] ));
NAND3X1 NAND3X1_1133 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n143_));
NAND3X1 NAND3X1_1134 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n144_));
NAND3X1 NAND3X1_1135 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n143_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n144_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n145_), .Y(\col_out[18] ));
NAND3X1 NAND3X1_1136 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n147_));
NAND3X1 NAND3X1_1137 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n148_));
NAND3X1 NAND3X1_1138 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n147_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n148_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n149_), .Y(\col_out[19] ));
NAND3X1 NAND3X1_1139 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n151_));
NAND3X1 NAND3X1_114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3092_), .B(AES_CORE_DATAPATH__abc_15863_new_n3093_), .C(AES_CORE_DATAPATH__abc_15863_new_n3095_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3096_));
NAND3X1 NAND3X1_1140 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n152_));
NAND3X1 NAND3X1_1141 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n151_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n152_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n153_), .Y(\col_out[20] ));
NAND3X1 NAND3X1_1142 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n155_));
NAND3X1 NAND3X1_1143 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n156_));
NAND3X1 NAND3X1_1144 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n155_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n156_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n157_), .Y(\col_out[21] ));
NAND3X1 NAND3X1_1145 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n159_));
NAND3X1 NAND3X1_1146 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n160_));
NAND3X1 NAND3X1_1147 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n159_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n160_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n161_), .Y(\col_out[22] ));
NAND3X1 NAND3X1_1148 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n163_));
NAND3X1 NAND3X1_1149 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n164_));
NAND3X1 NAND3X1_115 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2730_), .B(AES_CORE_DATAPATH__abc_15863_new_n2739_), .C(AES_CORE_DATAPATH__abc_15863_new_n3104_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3105_));
NAND3X1 NAND3X1_1150 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n163_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n164_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n165_), .Y(\col_out[23] ));
NAND3X1 NAND3X1_1151 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n167_));
NAND3X1 NAND3X1_1152 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n168_));
NAND3X1 NAND3X1_1153 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n167_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n168_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n169_), .Y(\col_out[24] ));
NAND3X1 NAND3X1_1154 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n171_));
NAND3X1 NAND3X1_1155 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n172_));
NAND3X1 NAND3X1_1156 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n171_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n172_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n173_), .Y(\col_out[25] ));
NAND3X1 NAND3X1_1157 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n175_));
NAND3X1 NAND3X1_1158 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n176_));
NAND3X1 NAND3X1_1159 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n175_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n176_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n177_), .Y(\col_out[26] ));
NAND3X1 NAND3X1_116 ( .A(AES_CORE_DATAPATH_col_0__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3119_));
NAND3X1 NAND3X1_1160 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n179_));
NAND3X1 NAND3X1_1161 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n180_));
NAND3X1 NAND3X1_1162 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n179_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n180_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n181_), .Y(\col_out[27] ));
NAND3X1 NAND3X1_1163 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n183_));
NAND3X1 NAND3X1_1164 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n184_));
NAND3X1 NAND3X1_1165 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n183_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n184_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n185_), .Y(\col_out[28] ));
NAND3X1 NAND3X1_1166 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n187_));
NAND3X1 NAND3X1_1167 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n188_));
NAND3X1 NAND3X1_1168 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n187_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n188_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n189_), .Y(\col_out[29] ));
NAND3X1 NAND3X1_1169 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n191_));
NAND3X1 NAND3X1_117 ( .A(AES_CORE_DATAPATH_col_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3120_));
NAND3X1 NAND3X1_1170 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n192_));
NAND3X1 NAND3X1_1171 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n191_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n192_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n193_), .Y(\col_out[30] ));
NAND3X1 NAND3X1_1172 ( .A(\data_type[0] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n195_));
NAND3X1 NAND3X1_1173 ( .A(\data_type[1] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n196_));
NAND3X1 NAND3X1_1174 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n195_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n196_), .C(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n197_), .Y(\col_out[31] ));
NAND3X1 NAND3X1_118 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3121_));
NAND3X1 NAND3X1_119 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3119_), .B(AES_CORE_DATAPATH__abc_15863_new_n3121_), .C(AES_CORE_DATAPATH__abc_15863_new_n3120_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3122_));
NAND3X1 NAND3X1_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_DATAPATH__abc_15863_new_n2724_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2725_));
NAND3X1 NAND3X1_120 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2748_), .B(AES_CORE_DATAPATH__abc_15863_new_n2750_), .C(AES_CORE_DATAPATH__abc_15863_new_n3128_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3129_));
NAND3X1 NAND3X1_121 ( .A(AES_CORE_DATAPATH_col_0__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3141_));
NAND3X1 NAND3X1_122 ( .A(AES_CORE_DATAPATH_col_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3142_));
NAND3X1 NAND3X1_123 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3143_));
NAND3X1 NAND3X1_124 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3141_), .B(AES_CORE_DATAPATH__abc_15863_new_n3143_), .C(AES_CORE_DATAPATH__abc_15863_new_n3142_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3144_));
NAND3X1 NAND3X1_125 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2761_), .B(AES_CORE_DATAPATH__abc_15863_new_n2763_), .C(AES_CORE_DATAPATH__abc_15863_new_n3150_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3151_));
NAND3X1 NAND3X1_126 ( .A(AES_CORE_DATAPATH_col_0__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3163_));
NAND3X1 NAND3X1_127 ( .A(AES_CORE_DATAPATH_col_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3164_));
NAND3X1 NAND3X1_128 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3165_));
NAND3X1 NAND3X1_129 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3163_), .B(AES_CORE_DATAPATH__abc_15863_new_n3165_), .C(AES_CORE_DATAPATH__abc_15863_new_n3164_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3166_));
NAND3X1 NAND3X1_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2712_), .B(AES_CORE_DATAPATH__abc_15863_new_n2723_), .C(AES_CORE_DATAPATH__abc_15863_new_n2725_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2726_));
NAND3X1 NAND3X1_130 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2769_), .B(AES_CORE_DATAPATH__abc_15863_new_n2773_), .C(AES_CORE_DATAPATH__abc_15863_new_n3171_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3172_));
NAND3X1 NAND3X1_131 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3172_), .C(AES_CORE_DATAPATH__abc_15863_new_n3174_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3175_));
NAND3X1 NAND3X1_132 ( .A(AES_CORE_DATAPATH_col_0__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3186_));
NAND3X1 NAND3X1_133 ( .A(AES_CORE_DATAPATH_col_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3187_));
NAND3X1 NAND3X1_134 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3188_));
NAND3X1 NAND3X1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3186_), .B(AES_CORE_DATAPATH__abc_15863_new_n3188_), .C(AES_CORE_DATAPATH__abc_15863_new_n3187_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3189_));
NAND3X1 NAND3X1_136 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2779_), .B(AES_CORE_DATAPATH__abc_15863_new_n2783_), .C(AES_CORE_DATAPATH__abc_15863_new_n3195_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3196_));
NAND3X1 NAND3X1_137 ( .A(AES_CORE_DATAPATH_col_0__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3208_));
NAND3X1 NAND3X1_138 ( .A(AES_CORE_DATAPATH_col_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3209_));
NAND3X1 NAND3X1_139 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3210_));
NAND3X1 NAND3X1_14 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2731_));
NAND3X1 NAND3X1_140 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3208_), .B(AES_CORE_DATAPATH__abc_15863_new_n3210_), .C(AES_CORE_DATAPATH__abc_15863_new_n3209_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3211_));
NAND3X1 NAND3X1_141 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2791_), .B(AES_CORE_DATAPATH__abc_15863_new_n2793_), .C(AES_CORE_DATAPATH__abc_15863_new_n3217_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3218_));
NAND3X1 NAND3X1_142 ( .A(AES_CORE_DATAPATH_col_0__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3230_));
NAND3X1 NAND3X1_143 ( .A(AES_CORE_DATAPATH_col_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3231_));
NAND3X1 NAND3X1_144 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3232_));
NAND3X1 NAND3X1_145 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3230_), .B(AES_CORE_DATAPATH__abc_15863_new_n3232_), .C(AES_CORE_DATAPATH__abc_15863_new_n3231_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3233_));
NAND3X1 NAND3X1_146 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2799_), .B(AES_CORE_DATAPATH__abc_15863_new_n2803_), .C(AES_CORE_DATAPATH__abc_15863_new_n3239_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3240_));
NAND3X1 NAND3X1_147 ( .A(AES_CORE_DATAPATH_col_0__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3252_));
NAND3X1 NAND3X1_148 ( .A(AES_CORE_DATAPATH_col_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3253_));
NAND3X1 NAND3X1_149 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3254_));
NAND3X1 NAND3X1_15 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2736_));
NAND3X1 NAND3X1_150 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3252_), .B(AES_CORE_DATAPATH__abc_15863_new_n3254_), .C(AES_CORE_DATAPATH__abc_15863_new_n3253_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3255_));
NAND3X1 NAND3X1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2812_), .B(AES_CORE_DATAPATH__abc_15863_new_n2814_), .C(AES_CORE_DATAPATH__abc_15863_new_n3261_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3262_));
NAND3X1 NAND3X1_152 ( .A(AES_CORE_DATAPATH_col_0__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3274_));
NAND3X1 NAND3X1_153 ( .A(AES_CORE_DATAPATH_col_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3275_));
NAND3X1 NAND3X1_154 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3276_));
NAND3X1 NAND3X1_155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3274_), .B(AES_CORE_DATAPATH__abc_15863_new_n3276_), .C(AES_CORE_DATAPATH__abc_15863_new_n3275_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3277_));
NAND3X1 NAND3X1_156 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2825_), .B(AES_CORE_DATAPATH__abc_15863_new_n2827_), .C(AES_CORE_DATAPATH__abc_15863_new_n3283_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3284_));
NAND3X1 NAND3X1_157 ( .A(AES_CORE_DATAPATH_col_0__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3296_));
NAND3X1 NAND3X1_158 ( .A(AES_CORE_DATAPATH_col_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3297_));
NAND3X1 NAND3X1_159 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3298_));
NAND3X1 NAND3X1_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2731_), .B(AES_CORE_DATAPATH__abc_15863_new_n2736_), .C(AES_CORE_DATAPATH__abc_15863_new_n2738_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2739_));
NAND3X1 NAND3X1_160 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3296_), .B(AES_CORE_DATAPATH__abc_15863_new_n3298_), .C(AES_CORE_DATAPATH__abc_15863_new_n3297_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3299_));
NAND3X1 NAND3X1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2837_), .B(AES_CORE_DATAPATH__abc_15863_new_n2839_), .C(AES_CORE_DATAPATH__abc_15863_new_n3303_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3304_));
NAND3X1 NAND3X1_162 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3304_), .C(AES_CORE_DATAPATH__abc_15863_new_n3306_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3307_));
NAND3X1 NAND3X1_163 ( .A(AES_CORE_DATAPATH_col_0__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3318_));
NAND3X1 NAND3X1_164 ( .A(AES_CORE_DATAPATH_col_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3319_));
NAND3X1 NAND3X1_165 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3320_));
NAND3X1 NAND3X1_166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3318_), .B(AES_CORE_DATAPATH__abc_15863_new_n3320_), .C(AES_CORE_DATAPATH__abc_15863_new_n3319_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3321_));
NAND3X1 NAND3X1_167 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2848_), .B(AES_CORE_DATAPATH__abc_15863_new_n2850_), .C(AES_CORE_DATAPATH__abc_15863_new_n3327_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3328_));
NAND3X1 NAND3X1_168 ( .A(AES_CORE_DATAPATH_col_0__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3340_));
NAND3X1 NAND3X1_169 ( .A(AES_CORE_DATAPATH_col_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3341_));
NAND3X1 NAND3X1_17 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2745_));
NAND3X1 NAND3X1_170 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3342_));
NAND3X1 NAND3X1_171 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3340_), .B(AES_CORE_DATAPATH__abc_15863_new_n3342_), .C(AES_CORE_DATAPATH__abc_15863_new_n3341_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3343_));
NAND3X1 NAND3X1_172 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2857_), .B(AES_CORE_DATAPATH__abc_15863_new_n2859_), .C(AES_CORE_DATAPATH__abc_15863_new_n3347_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3348_));
NAND3X1 NAND3X1_173 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3348_), .C(AES_CORE_DATAPATH__abc_15863_new_n3350_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3351_));
NAND3X1 NAND3X1_174 ( .A(AES_CORE_DATAPATH_col_0__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3362_));
NAND3X1 NAND3X1_175 ( .A(AES_CORE_DATAPATH_col_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3363_));
NAND3X1 NAND3X1_176 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3364_));
NAND3X1 NAND3X1_177 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3362_), .B(AES_CORE_DATAPATH__abc_15863_new_n3364_), .C(AES_CORE_DATAPATH__abc_15863_new_n3363_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3365_));
NAND3X1 NAND3X1_178 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2867_), .B(AES_CORE_DATAPATH__abc_15863_new_n2869_), .C(AES_CORE_DATAPATH__abc_15863_new_n3371_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3372_));
NAND3X1 NAND3X1_179 ( .A(AES_CORE_DATAPATH_col_0__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3384_));
NAND3X1 NAND3X1_18 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2746_));
NAND3X1 NAND3X1_180 ( .A(AES_CORE_DATAPATH_col_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3385_));
NAND3X1 NAND3X1_181 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3386_));
NAND3X1 NAND3X1_182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3384_), .B(AES_CORE_DATAPATH__abc_15863_new_n3386_), .C(AES_CORE_DATAPATH__abc_15863_new_n3385_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3387_));
NAND3X1 NAND3X1_183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2875_), .B(AES_CORE_DATAPATH__abc_15863_new_n2879_), .C(AES_CORE_DATAPATH__abc_15863_new_n3391_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3392_));
NAND3X1 NAND3X1_184 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3392_), .C(AES_CORE_DATAPATH__abc_15863_new_n3394_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3395_));
NAND3X1 NAND3X1_185 ( .A(AES_CORE_DATAPATH_col_0__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3406_));
NAND3X1 NAND3X1_186 ( .A(AES_CORE_DATAPATH_col_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3407_));
NAND3X1 NAND3X1_187 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3408_));
NAND3X1 NAND3X1_188 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3406_), .B(AES_CORE_DATAPATH__abc_15863_new_n3408_), .C(AES_CORE_DATAPATH__abc_15863_new_n3407_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3409_));
NAND3X1 NAND3X1_189 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2887_), .B(AES_CORE_DATAPATH__abc_15863_new_n2889_), .C(AES_CORE_DATAPATH__abc_15863_new_n3415_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3416_));
NAND3X1 NAND3X1_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2745_), .B(AES_CORE_DATAPATH__abc_15863_new_n2746_), .C(AES_CORE_DATAPATH__abc_15863_new_n2747_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2748_));
NAND3X1 NAND3X1_190 ( .A(AES_CORE_DATAPATH_col_0__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3428_));
NAND3X1 NAND3X1_191 ( .A(AES_CORE_DATAPATH_col_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3429_));
NAND3X1 NAND3X1_192 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3430_));
NAND3X1 NAND3X1_193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3428_), .B(AES_CORE_DATAPATH__abc_15863_new_n3430_), .C(AES_CORE_DATAPATH__abc_15863_new_n3429_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3431_));
NAND3X1 NAND3X1_194 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2895_), .B(AES_CORE_DATAPATH__abc_15863_new_n2899_), .C(AES_CORE_DATAPATH__abc_15863_new_n3435_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3436_));
NAND3X1 NAND3X1_195 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3436_), .C(AES_CORE_DATAPATH__abc_15863_new_n3438_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3439_));
NAND3X1 NAND3X1_196 ( .A(AES_CORE_DATAPATH_col_0__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3450_));
NAND3X1 NAND3X1_197 ( .A(AES_CORE_DATAPATH_col_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3451_));
NAND3X1 NAND3X1_198 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3452_));
NAND3X1 NAND3X1_199 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3450_), .B(AES_CORE_DATAPATH__abc_15863_new_n3452_), .C(AES_CORE_DATAPATH__abc_15863_new_n3451_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3453_));
NAND3X1 NAND3X1_2 ( .A(AES_CORE_CONTROL_UNIT_state_0_), .B(start), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n97_));
NAND3X1 NAND3X1_20 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2758_));
NAND3X1 NAND3X1_200 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2906_), .B(AES_CORE_DATAPATH__abc_15863_new_n2910_), .C(AES_CORE_DATAPATH__abc_15863_new_n3459_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3460_));
NAND3X1 NAND3X1_201 ( .A(AES_CORE_DATAPATH_col_0__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3472_));
NAND3X1 NAND3X1_202 ( .A(AES_CORE_DATAPATH_col_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3473_));
NAND3X1 NAND3X1_203 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3474_));
NAND3X1 NAND3X1_204 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3472_), .B(AES_CORE_DATAPATH__abc_15863_new_n3474_), .C(AES_CORE_DATAPATH__abc_15863_new_n3473_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3475_));
NAND3X1 NAND3X1_205 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2915_), .B(AES_CORE_DATAPATH__abc_15863_new_n2919_), .C(AES_CORE_DATAPATH__abc_15863_new_n3479_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3480_));
NAND3X1 NAND3X1_206 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3480_), .C(AES_CORE_DATAPATH__abc_15863_new_n3482_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3483_));
NAND3X1 NAND3X1_207 ( .A(AES_CORE_DATAPATH_col_0__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3494_));
NAND3X1 NAND3X1_208 ( .A(AES_CORE_DATAPATH_col_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3495_));
NAND3X1 NAND3X1_209 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3496_));
NAND3X1 NAND3X1_21 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2759_));
NAND3X1 NAND3X1_210 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3494_), .B(AES_CORE_DATAPATH__abc_15863_new_n3496_), .C(AES_CORE_DATAPATH__abc_15863_new_n3495_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3497_));
NAND3X1 NAND3X1_211 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2925_), .B(AES_CORE_DATAPATH__abc_15863_new_n2929_), .C(AES_CORE_DATAPATH__abc_15863_new_n3503_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3504_));
NAND3X1 NAND3X1_212 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3504_), .C(AES_CORE_DATAPATH__abc_15863_new_n3502_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3505_));
NAND3X1 NAND3X1_213 ( .A(AES_CORE_DATAPATH_col_0__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3516_));
NAND3X1 NAND3X1_214 ( .A(AES_CORE_DATAPATH_col_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3517_));
NAND3X1 NAND3X1_215 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3518_));
NAND3X1 NAND3X1_216 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3516_), .B(AES_CORE_DATAPATH__abc_15863_new_n3518_), .C(AES_CORE_DATAPATH__abc_15863_new_n3517_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3519_));
NAND3X1 NAND3X1_217 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2935_), .B(AES_CORE_DATAPATH__abc_15863_new_n2939_), .C(AES_CORE_DATAPATH__abc_15863_new_n3523_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3524_));
NAND3X1 NAND3X1_218 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3524_), .C(AES_CORE_DATAPATH__abc_15863_new_n3526_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3527_));
NAND3X1 NAND3X1_219 ( .A(AES_CORE_DATAPATH_col_0__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3538_));
NAND3X1 NAND3X1_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2758_), .B(AES_CORE_DATAPATH__abc_15863_new_n2759_), .C(AES_CORE_DATAPATH__abc_15863_new_n2760_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2761_));
NAND3X1 NAND3X1_220 ( .A(AES_CORE_DATAPATH_col_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3539_));
NAND3X1 NAND3X1_221 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3540_));
NAND3X1 NAND3X1_222 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3538_), .B(AES_CORE_DATAPATH__abc_15863_new_n3540_), .C(AES_CORE_DATAPATH__abc_15863_new_n3539_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3541_));
NAND3X1 NAND3X1_223 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2946_), .B(AES_CORE_DATAPATH__abc_15863_new_n2950_), .C(AES_CORE_DATAPATH__abc_15863_new_n3547_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3548_));
NAND3X1 NAND3X1_224 ( .A(AES_CORE_DATAPATH_col_0__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3560_));
NAND3X1 NAND3X1_225 ( .A(AES_CORE_DATAPATH_col_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3561_));
NAND3X1 NAND3X1_226 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3562_));
NAND3X1 NAND3X1_227 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3560_), .B(AES_CORE_DATAPATH__abc_15863_new_n3562_), .C(AES_CORE_DATAPATH__abc_15863_new_n3561_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3563_));
NAND3X1 NAND3X1_228 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2958_), .B(AES_CORE_DATAPATH__abc_15863_new_n2962_), .C(AES_CORE_DATAPATH__abc_15863_new_n3567_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3568_));
NAND3X1 NAND3X1_229 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3568_), .C(AES_CORE_DATAPATH__abc_15863_new_n3570_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3571_));
NAND3X1 NAND3X1_23 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2770_));
NAND3X1 NAND3X1_230 ( .A(AES_CORE_DATAPATH_col_0__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3582_));
NAND3X1 NAND3X1_231 ( .A(AES_CORE_DATAPATH_col_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3583_));
NAND3X1 NAND3X1_232 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3584_));
NAND3X1 NAND3X1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3582_), .B(AES_CORE_DATAPATH__abc_15863_new_n3584_), .C(AES_CORE_DATAPATH__abc_15863_new_n3583_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3585_));
NAND3X1 NAND3X1_234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2968_), .B(AES_CORE_DATAPATH__abc_15863_new_n2972_), .C(AES_CORE_DATAPATH__abc_15863_new_n3591_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3592_));
NAND3X1 NAND3X1_235 ( .A(AES_CORE_DATAPATH_col_0__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3604_));
NAND3X1 NAND3X1_236 ( .A(AES_CORE_DATAPATH_col_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3605_));
NAND3X1 NAND3X1_237 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3606_));
NAND3X1 NAND3X1_238 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3604_), .B(AES_CORE_DATAPATH__abc_15863_new_n3606_), .C(AES_CORE_DATAPATH__abc_15863_new_n3605_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3607_));
NAND3X1 NAND3X1_239 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2979_), .B(AES_CORE_DATAPATH__abc_15863_new_n2983_), .C(AES_CORE_DATAPATH__abc_15863_new_n3613_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3614_));
NAND3X1 NAND3X1_24 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2771_));
NAND3X1 NAND3X1_240 ( .A(AES_CORE_DATAPATH_col_0__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3626_));
NAND3X1 NAND3X1_241 ( .A(AES_CORE_DATAPATH_col_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3627_));
NAND3X1 NAND3X1_242 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3628_));
NAND3X1 NAND3X1_243 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3626_), .B(AES_CORE_DATAPATH__abc_15863_new_n3628_), .C(AES_CORE_DATAPATH__abc_15863_new_n3627_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3629_));
NAND3X1 NAND3X1_244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2994_), .B(AES_CORE_DATAPATH__abc_15863_new_n2996_), .C(AES_CORE_DATAPATH__abc_15863_new_n3635_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3636_));
NAND3X1 NAND3X1_245 ( .A(AES_CORE_DATAPATH_col_0__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3648_));
NAND3X1 NAND3X1_246 ( .A(AES_CORE_DATAPATH_col_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3649_));
NAND3X1 NAND3X1_247 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3650_));
NAND3X1 NAND3X1_248 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3648_), .B(AES_CORE_DATAPATH__abc_15863_new_n3650_), .C(AES_CORE_DATAPATH__abc_15863_new_n3649_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3651_));
NAND3X1 NAND3X1_249 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3006_), .B(AES_CORE_DATAPATH__abc_15863_new_n3008_), .C(AES_CORE_DATAPATH__abc_15863_new_n3655_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3656_));
NAND3X1 NAND3X1_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2770_), .B(AES_CORE_DATAPATH__abc_15863_new_n2771_), .C(AES_CORE_DATAPATH__abc_15863_new_n2772_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2773_));
NAND3X1 NAND3X1_250 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3656_), .C(AES_CORE_DATAPATH__abc_15863_new_n3658_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3659_));
NAND3X1 NAND3X1_251 ( .A(AES_CORE_DATAPATH_col_0__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3670_));
NAND3X1 NAND3X1_252 ( .A(AES_CORE_DATAPATH_col_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3671_));
NAND3X1 NAND3X1_253 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3672_));
NAND3X1 NAND3X1_254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3670_), .B(AES_CORE_DATAPATH__abc_15863_new_n3672_), .C(AES_CORE_DATAPATH__abc_15863_new_n3671_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3673_));
NAND3X1 NAND3X1_255 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3016_), .B(AES_CORE_DATAPATH__abc_15863_new_n3018_), .C(AES_CORE_DATAPATH__abc_15863_new_n3679_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3680_));
NAND3X1 NAND3X1_256 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3680_), .C(AES_CORE_DATAPATH__abc_15863_new_n3678_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3681_));
NAND3X1 NAND3X1_257 ( .A(AES_CORE_DATAPATH_col_0__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3692_));
NAND3X1 NAND3X1_258 ( .A(AES_CORE_DATAPATH_col_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3693_));
NAND3X1 NAND3X1_259 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3694_));
NAND3X1 NAND3X1_26 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2780_));
NAND3X1 NAND3X1_260 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3692_), .B(AES_CORE_DATAPATH__abc_15863_new_n3694_), .C(AES_CORE_DATAPATH__abc_15863_new_n3693_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3695_));
NAND3X1 NAND3X1_261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3026_), .B(AES_CORE_DATAPATH__abc_15863_new_n3028_), .C(AES_CORE_DATAPATH__abc_15863_new_n3701_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3702_));
NAND3X1 NAND3X1_262 ( .A(AES_CORE_DATAPATH_col_0__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3714_));
NAND3X1 NAND3X1_263 ( .A(AES_CORE_DATAPATH_col_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3715_));
NAND3X1 NAND3X1_264 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3716_));
NAND3X1 NAND3X1_265 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3714_), .B(AES_CORE_DATAPATH__abc_15863_new_n3716_), .C(AES_CORE_DATAPATH__abc_15863_new_n3715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3717_));
NAND3X1 NAND3X1_266 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3037_), .B(AES_CORE_DATAPATH__abc_15863_new_n3039_), .C(AES_CORE_DATAPATH__abc_15863_new_n3721_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3722_));
NAND3X1 NAND3X1_267 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3722_), .C(AES_CORE_DATAPATH__abc_15863_new_n3724_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3725_));
NAND3X1 NAND3X1_268 ( .A(AES_CORE_DATAPATH_col_0__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3736_));
NAND3X1 NAND3X1_269 ( .A(AES_CORE_DATAPATH_col_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3737_));
NAND3X1 NAND3X1_27 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2781_));
NAND3X1 NAND3X1_270 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3738_));
NAND3X1 NAND3X1_271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3736_), .B(AES_CORE_DATAPATH__abc_15863_new_n3738_), .C(AES_CORE_DATAPATH__abc_15863_new_n3737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3739_));
NAND3X1 NAND3X1_272 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3047_), .B(AES_CORE_DATAPATH__abc_15863_new_n3049_), .C(AES_CORE_DATAPATH__abc_15863_new_n3745_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3746_));
NAND3X1 NAND3X1_273 ( .A(AES_CORE_DATAPATH_col_0__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3758_));
NAND3X1 NAND3X1_274 ( .A(AES_CORE_DATAPATH_col_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3759_));
NAND3X1 NAND3X1_275 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3760_));
NAND3X1 NAND3X1_276 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3758_), .B(AES_CORE_DATAPATH__abc_15863_new_n3760_), .C(AES_CORE_DATAPATH__abc_15863_new_n3759_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3761_));
NAND3X1 NAND3X1_277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3057_), .B(AES_CORE_DATAPATH__abc_15863_new_n3059_), .C(AES_CORE_DATAPATH__abc_15863_new_n3767_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3768_));
NAND3X1 NAND3X1_278 ( .A(AES_CORE_DATAPATH_col_0__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n3087_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3780_));
NAND3X1 NAND3X1_279 ( .A(AES_CORE_DATAPATH_col_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3094_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3781_));
NAND3X1 NAND3X1_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2780_), .B(AES_CORE_DATAPATH__abc_15863_new_n2781_), .C(AES_CORE_DATAPATH__abc_15863_new_n2782_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2783_));
NAND3X1 NAND3X1_280 ( .A(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .B(AES_CORE_DATAPATH__abc_15863_new_n3082_), .C(AES_CORE_DATAPATH__abc_15863_new_n3091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3782_));
NAND3X1 NAND3X1_281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3780_), .B(AES_CORE_DATAPATH__abc_15863_new_n3782_), .C(AES_CORE_DATAPATH__abc_15863_new_n3781_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3783_));
NAND3X1 NAND3X1_282 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3064_), .B(AES_CORE_DATAPATH__abc_15863_new_n3068_), .C(AES_CORE_DATAPATH__abc_15863_new_n3787_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3788_));
NAND3X1 NAND3X1_283 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n3788_), .C(AES_CORE_DATAPATH__abc_15863_new_n3790_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3791_));
NAND3X1 NAND3X1_284 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4591_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4590_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4594_));
NAND3X1 NAND3X1_285 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4595_), .B(AES_CORE_DATAPATH__abc_15863_new_n4609_), .C(AES_CORE_DATAPATH__abc_15863_new_n4594_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4610_));
NAND3X1 NAND3X1_286 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4613_), .B(AES_CORE_DATAPATH__abc_15863_new_n4615_), .C(AES_CORE_DATAPATH__abc_15863_new_n4611_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4616_));
NAND3X1 NAND3X1_287 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4583_), .B(AES_CORE_DATAPATH__abc_15863_new_n4586_), .C(AES_CORE_DATAPATH__abc_15863_new_n4629_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4630_));
NAND3X1 NAND3X1_288 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4639_), .B(AES_CORE_DATAPATH__abc_15863_new_n4650_), .C(AES_CORE_DATAPATH__abc_15863_new_n4637_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4651_));
NAND3X1 NAND3X1_289 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2748_), .B(AES_CORE_DATAPATH__abc_15863_new_n2750_), .C(AES_CORE_DATAPATH__abc_15863_new_n3126_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4652_));
NAND3X1 NAND3X1_29 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2788_));
NAND3X1 NAND3X1_290 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n4652_), .C(AES_CORE_DATAPATH__abc_15863_new_n4653_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4654_));
NAND3X1 NAND3X1_291 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4636_), .B(AES_CORE_DATAPATH__abc_15863_new_n4668_), .C(AES_CORE_DATAPATH__abc_15863_new_n4667_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4669_));
NAND3X1 NAND3X1_292 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4678_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4677_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4679_));
NAND3X1 NAND3X1_293 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4680_), .B(AES_CORE_DATAPATH__abc_15863_new_n4691_), .C(AES_CORE_DATAPATH__abc_15863_new_n4679_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4692_));
NAND3X1 NAND3X1_294 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4695_), .B(AES_CORE_DATAPATH__abc_15863_new_n4697_), .C(AES_CORE_DATAPATH__abc_15863_new_n4693_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4698_));
NAND3X1 NAND3X1_295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4675_), .B(AES_CORE_DATAPATH__abc_15863_new_n4707_), .C(AES_CORE_DATAPATH__abc_15863_new_n4706_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4708_));
NAND3X1 NAND3X1_296 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2769_), .B(AES_CORE_DATAPATH__abc_15863_new_n2773_), .C(AES_CORE_DATAPATH__abc_15863_new_n3173_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4716_));
NAND3X1 NAND3X1_297 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4720_), .B(AES_CORE_DATAPATH__abc_15863_new_n4731_), .C(AES_CORE_DATAPATH__abc_15863_new_n4718_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4732_));
NAND3X1 NAND3X1_298 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4714_), .B(AES_CORE_DATAPATH__abc_15863_new_n4747_), .C(AES_CORE_DATAPATH__abc_15863_new_n4744_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4748_));
NAND3X1 NAND3X1_299 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4757_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4756_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4758_));
NAND3X1 NAND3X1_3 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .B(AES_CORE_CONTROL_UNIT_state_12_), .C(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n100_));
NAND3X1 NAND3X1_30 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2789_));
NAND3X1 NAND3X1_300 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4759_), .B(AES_CORE_DATAPATH__abc_15863_new_n4767_), .C(AES_CORE_DATAPATH__abc_15863_new_n4758_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4768_));
NAND3X1 NAND3X1_301 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4771_), .B(AES_CORE_DATAPATH__abc_15863_new_n4773_), .C(AES_CORE_DATAPATH__abc_15863_new_n4769_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4774_));
NAND3X1 NAND3X1_302 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4754_), .B(AES_CORE_DATAPATH__abc_15863_new_n4783_), .C(AES_CORE_DATAPATH__abc_15863_new_n4782_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4784_));
NAND3X1 NAND3X1_303 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4793_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4792_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4794_));
NAND3X1 NAND3X1_304 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4795_), .B(AES_CORE_DATAPATH__abc_15863_new_n4806_), .C(AES_CORE_DATAPATH__abc_15863_new_n4794_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4807_));
NAND3X1 NAND3X1_305 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4810_), .B(AES_CORE_DATAPATH__abc_15863_new_n4812_), .C(AES_CORE_DATAPATH__abc_15863_new_n4808_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4813_));
NAND3X1 NAND3X1_306 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4790_), .B(AES_CORE_DATAPATH__abc_15863_new_n4822_), .C(AES_CORE_DATAPATH__abc_15863_new_n4821_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4823_));
NAND3X1 NAND3X1_307 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4832_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4831_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4833_));
NAND3X1 NAND3X1_308 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4834_), .B(AES_CORE_DATAPATH__abc_15863_new_n4842_), .C(AES_CORE_DATAPATH__abc_15863_new_n4833_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4843_));
NAND3X1 NAND3X1_309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4846_), .B(AES_CORE_DATAPATH__abc_15863_new_n4847_), .C(AES_CORE_DATAPATH__abc_15863_new_n4844_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4848_));
NAND3X1 NAND3X1_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2788_), .B(AES_CORE_DATAPATH__abc_15863_new_n2789_), .C(AES_CORE_DATAPATH__abc_15863_new_n2790_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2791_));
NAND3X1 NAND3X1_310 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4829_), .B(AES_CORE_DATAPATH__abc_15863_new_n4857_), .C(AES_CORE_DATAPATH__abc_15863_new_n4856_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4858_));
NAND3X1 NAND3X1_311 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4867_), .B(AES_CORE_DATAPATH__abc_15863_new_n4878_), .C(AES_CORE_DATAPATH__abc_15863_new_n4865_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4879_));
NAND3X1 NAND3X1_312 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2812_), .B(AES_CORE_DATAPATH__abc_15863_new_n2814_), .C(AES_CORE_DATAPATH__abc_15863_new_n3259_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4880_));
NAND3X1 NAND3X1_313 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n4880_), .C(AES_CORE_DATAPATH__abc_15863_new_n4881_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4882_));
NAND3X1 NAND3X1_314 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4864_), .B(AES_CORE_DATAPATH__abc_15863_new_n4896_), .C(AES_CORE_DATAPATH__abc_15863_new_n4895_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4897_));
NAND3X1 NAND3X1_315 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4906_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4905_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4907_));
NAND3X1 NAND3X1_316 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4908_), .B(AES_CORE_DATAPATH__abc_15863_new_n4916_), .C(AES_CORE_DATAPATH__abc_15863_new_n4907_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4917_));
NAND3X1 NAND3X1_317 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4920_), .B(AES_CORE_DATAPATH__abc_15863_new_n4921_), .C(AES_CORE_DATAPATH__abc_15863_new_n4918_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4922_));
NAND3X1 NAND3X1_318 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4903_), .B(AES_CORE_DATAPATH__abc_15863_new_n4931_), .C(AES_CORE_DATAPATH__abc_15863_new_n4930_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4932_));
NAND3X1 NAND3X1_319 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2837_), .B(AES_CORE_DATAPATH__abc_15863_new_n2839_), .C(AES_CORE_DATAPATH__abc_15863_new_n3305_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4940_));
NAND3X1 NAND3X1_32 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2800_));
NAND3X1 NAND3X1_320 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4944_), .B(AES_CORE_DATAPATH__abc_15863_new_n4955_), .C(AES_CORE_DATAPATH__abc_15863_new_n4942_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4956_));
NAND3X1 NAND3X1_321 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4938_), .B(AES_CORE_DATAPATH__abc_15863_new_n4970_), .C(AES_CORE_DATAPATH__abc_15863_new_n4968_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4971_));
NAND3X1 NAND3X1_322 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4980_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4979_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4981_));
NAND3X1 NAND3X1_323 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4982_), .B(AES_CORE_DATAPATH__abc_15863_new_n4993_), .C(AES_CORE_DATAPATH__abc_15863_new_n4981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4994_));
NAND3X1 NAND3X1_324 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4997_), .B(AES_CORE_DATAPATH__abc_15863_new_n4999_), .C(AES_CORE_DATAPATH__abc_15863_new_n4995_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5000_));
NAND3X1 NAND3X1_325 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4977_), .B(AES_CORE_DATAPATH__abc_15863_new_n5009_), .C(AES_CORE_DATAPATH__abc_15863_new_n5008_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5010_));
NAND3X1 NAND3X1_326 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2857_), .B(AES_CORE_DATAPATH__abc_15863_new_n2859_), .C(AES_CORE_DATAPATH__abc_15863_new_n3349_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5018_));
NAND3X1 NAND3X1_327 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5022_), .B(AES_CORE_DATAPATH__abc_15863_new_n5033_), .C(AES_CORE_DATAPATH__abc_15863_new_n5020_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5034_));
NAND3X1 NAND3X1_328 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5016_), .B(AES_CORE_DATAPATH__abc_15863_new_n5048_), .C(AES_CORE_DATAPATH__abc_15863_new_n5046_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5049_));
NAND3X1 NAND3X1_329 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5058_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5057_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5059_));
NAND3X1 NAND3X1_33 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2801_));
NAND3X1 NAND3X1_330 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5060_), .B(AES_CORE_DATAPATH__abc_15863_new_n5071_), .C(AES_CORE_DATAPATH__abc_15863_new_n5059_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5072_));
NAND3X1 NAND3X1_331 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5075_), .B(AES_CORE_DATAPATH__abc_15863_new_n5077_), .C(AES_CORE_DATAPATH__abc_15863_new_n5073_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5078_));
NAND3X1 NAND3X1_332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5055_), .B(AES_CORE_DATAPATH__abc_15863_new_n5087_), .C(AES_CORE_DATAPATH__abc_15863_new_n5086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5088_));
NAND3X1 NAND3X1_333 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2875_), .B(AES_CORE_DATAPATH__abc_15863_new_n2879_), .C(AES_CORE_DATAPATH__abc_15863_new_n3393_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5096_));
NAND3X1 NAND3X1_334 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5100_), .B(AES_CORE_DATAPATH__abc_15863_new_n5111_), .C(AES_CORE_DATAPATH__abc_15863_new_n5098_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5112_));
NAND3X1 NAND3X1_335 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5094_), .B(AES_CORE_DATAPATH__abc_15863_new_n5126_), .C(AES_CORE_DATAPATH__abc_15863_new_n5124_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5127_));
NAND3X1 NAND3X1_336 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5136_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5135_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5137_));
NAND3X1 NAND3X1_337 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5138_), .B(AES_CORE_DATAPATH__abc_15863_new_n5146_), .C(AES_CORE_DATAPATH__abc_15863_new_n5137_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5147_));
NAND3X1 NAND3X1_338 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5150_), .B(AES_CORE_DATAPATH__abc_15863_new_n5152_), .C(AES_CORE_DATAPATH__abc_15863_new_n5148_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5153_));
NAND3X1 NAND3X1_339 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5133_), .B(AES_CORE_DATAPATH__abc_15863_new_n5162_), .C(AES_CORE_DATAPATH__abc_15863_new_n5161_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5163_));
NAND3X1 NAND3X1_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2800_), .B(AES_CORE_DATAPATH__abc_15863_new_n2801_), .C(AES_CORE_DATAPATH__abc_15863_new_n2802_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2803_));
NAND3X1 NAND3X1_340 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2895_), .B(AES_CORE_DATAPATH__abc_15863_new_n2899_), .C(AES_CORE_DATAPATH__abc_15863_new_n3437_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5171_));
NAND3X1 NAND3X1_341 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5175_), .B(AES_CORE_DATAPATH__abc_15863_new_n5186_), .C(AES_CORE_DATAPATH__abc_15863_new_n5173_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5187_));
NAND3X1 NAND3X1_342 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5169_), .B(AES_CORE_DATAPATH__abc_15863_new_n5201_), .C(AES_CORE_DATAPATH__abc_15863_new_n5199_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5202_));
NAND3X1 NAND3X1_343 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5211_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5210_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5212_));
NAND3X1 NAND3X1_344 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5213_), .B(AES_CORE_DATAPATH__abc_15863_new_n5224_), .C(AES_CORE_DATAPATH__abc_15863_new_n5212_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5225_));
NAND3X1 NAND3X1_345 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5228_), .B(AES_CORE_DATAPATH__abc_15863_new_n5230_), .C(AES_CORE_DATAPATH__abc_15863_new_n5226_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5231_));
NAND3X1 NAND3X1_346 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5208_), .B(AES_CORE_DATAPATH__abc_15863_new_n5240_), .C(AES_CORE_DATAPATH__abc_15863_new_n5239_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5241_));
NAND3X1 NAND3X1_347 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2915_), .B(AES_CORE_DATAPATH__abc_15863_new_n2919_), .C(AES_CORE_DATAPATH__abc_15863_new_n3481_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5249_));
NAND3X1 NAND3X1_348 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5253_), .B(AES_CORE_DATAPATH__abc_15863_new_n5264_), .C(AES_CORE_DATAPATH__abc_15863_new_n5251_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5265_));
NAND3X1 NAND3X1_349 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5247_), .B(AES_CORE_DATAPATH__abc_15863_new_n5279_), .C(AES_CORE_DATAPATH__abc_15863_new_n5277_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5280_));
NAND3X1 NAND3X1_35 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2809_));
NAND3X1 NAND3X1_350 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2925_), .B(AES_CORE_DATAPATH__abc_15863_new_n2929_), .C(AES_CORE_DATAPATH__abc_15863_new_n3501_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5288_));
NAND3X1 NAND3X1_351 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5292_), .B(AES_CORE_DATAPATH__abc_15863_new_n5303_), .C(AES_CORE_DATAPATH__abc_15863_new_n5290_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5304_));
NAND3X1 NAND3X1_352 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5286_), .B(AES_CORE_DATAPATH__abc_15863_new_n5318_), .C(AES_CORE_DATAPATH__abc_15863_new_n5316_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5319_));
NAND3X1 NAND3X1_353 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2935_), .B(AES_CORE_DATAPATH__abc_15863_new_n2939_), .C(AES_CORE_DATAPATH__abc_15863_new_n3525_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5327_));
NAND3X1 NAND3X1_354 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5331_), .B(AES_CORE_DATAPATH__abc_15863_new_n5342_), .C(AES_CORE_DATAPATH__abc_15863_new_n5329_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5343_));
NAND3X1 NAND3X1_355 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5325_), .B(AES_CORE_DATAPATH__abc_15863_new_n5357_), .C(AES_CORE_DATAPATH__abc_15863_new_n5355_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5358_));
NAND3X1 NAND3X1_356 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5367_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5366_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5368_));
NAND3X1 NAND3X1_357 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5369_), .B(AES_CORE_DATAPATH__abc_15863_new_n5380_), .C(AES_CORE_DATAPATH__abc_15863_new_n5368_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5381_));
NAND3X1 NAND3X1_358 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5384_), .B(AES_CORE_DATAPATH__abc_15863_new_n5386_), .C(AES_CORE_DATAPATH__abc_15863_new_n5382_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5387_));
NAND3X1 NAND3X1_359 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5364_), .B(AES_CORE_DATAPATH__abc_15863_new_n5396_), .C(AES_CORE_DATAPATH__abc_15863_new_n5395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5397_));
NAND3X1 NAND3X1_36 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2810_));
NAND3X1 NAND3X1_360 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2958_), .B(AES_CORE_DATAPATH__abc_15863_new_n2962_), .C(AES_CORE_DATAPATH__abc_15863_new_n3569_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5405_));
NAND3X1 NAND3X1_361 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5409_), .B(AES_CORE_DATAPATH__abc_15863_new_n5420_), .C(AES_CORE_DATAPATH__abc_15863_new_n5407_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5421_));
NAND3X1 NAND3X1_362 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5403_), .B(AES_CORE_DATAPATH__abc_15863_new_n5435_), .C(AES_CORE_DATAPATH__abc_15863_new_n5433_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5436_));
NAND3X1 NAND3X1_363 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5445_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5444_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5446_));
NAND3X1 NAND3X1_364 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5447_), .B(AES_CORE_DATAPATH__abc_15863_new_n5455_), .C(AES_CORE_DATAPATH__abc_15863_new_n5446_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5456_));
NAND3X1 NAND3X1_365 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5459_), .B(AES_CORE_DATAPATH__abc_15863_new_n5461_), .C(AES_CORE_DATAPATH__abc_15863_new_n5457_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5462_));
NAND3X1 NAND3X1_366 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5442_), .B(AES_CORE_DATAPATH__abc_15863_new_n5471_), .C(AES_CORE_DATAPATH__abc_15863_new_n5470_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5472_));
NAND3X1 NAND3X1_367 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5481_), .B(AES_CORE_DATAPATH__abc_15863_new_n5492_), .C(AES_CORE_DATAPATH__abc_15863_new_n5479_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5493_));
NAND3X1 NAND3X1_368 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2979_), .B(AES_CORE_DATAPATH__abc_15863_new_n2983_), .C(AES_CORE_DATAPATH__abc_15863_new_n3611_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5494_));
NAND3X1 NAND3X1_369 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3168_), .B(AES_CORE_DATAPATH__abc_15863_new_n5494_), .C(AES_CORE_DATAPATH__abc_15863_new_n5495_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5496_));
NAND3X1 NAND3X1_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2809_), .B(AES_CORE_DATAPATH__abc_15863_new_n2810_), .C(AES_CORE_DATAPATH__abc_15863_new_n2811_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2812_));
NAND3X1 NAND3X1_370 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5478_), .B(AES_CORE_DATAPATH__abc_15863_new_n5510_), .C(AES_CORE_DATAPATH__abc_15863_new_n5509_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5511_));
NAND3X1 NAND3X1_371 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5520_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5519_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5521_));
NAND3X1 NAND3X1_372 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5522_), .B(AES_CORE_DATAPATH__abc_15863_new_n5533_), .C(AES_CORE_DATAPATH__abc_15863_new_n5521_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5534_));
NAND3X1 NAND3X1_373 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5537_), .B(AES_CORE_DATAPATH__abc_15863_new_n5539_), .C(AES_CORE_DATAPATH__abc_15863_new_n5535_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5540_));
NAND3X1 NAND3X1_374 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5517_), .B(AES_CORE_DATAPATH__abc_15863_new_n5549_), .C(AES_CORE_DATAPATH__abc_15863_new_n5548_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5550_));
NAND3X1 NAND3X1_375 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3006_), .B(AES_CORE_DATAPATH__abc_15863_new_n3008_), .C(AES_CORE_DATAPATH__abc_15863_new_n3657_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5558_));
NAND3X1 NAND3X1_376 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5562_), .B(AES_CORE_DATAPATH__abc_15863_new_n5573_), .C(AES_CORE_DATAPATH__abc_15863_new_n5560_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5574_));
NAND3X1 NAND3X1_377 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5556_), .B(AES_CORE_DATAPATH__abc_15863_new_n5588_), .C(AES_CORE_DATAPATH__abc_15863_new_n5586_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5589_));
NAND3X1 NAND3X1_378 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3016_), .B(AES_CORE_DATAPATH__abc_15863_new_n3018_), .C(AES_CORE_DATAPATH__abc_15863_new_n3677_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5597_));
NAND3X1 NAND3X1_379 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5601_), .B(AES_CORE_DATAPATH__abc_15863_new_n5612_), .C(AES_CORE_DATAPATH__abc_15863_new_n5599_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5613_));
NAND3X1 NAND3X1_38 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2822_));
NAND3X1 NAND3X1_380 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5595_), .B(AES_CORE_DATAPATH__abc_15863_new_n5627_), .C(AES_CORE_DATAPATH__abc_15863_new_n5625_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5628_));
NAND3X1 NAND3X1_381 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5637_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5636_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5638_));
NAND3X1 NAND3X1_382 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5639_), .B(AES_CORE_DATAPATH__abc_15863_new_n5650_), .C(AES_CORE_DATAPATH__abc_15863_new_n5638_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5651_));
NAND3X1 NAND3X1_383 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5654_), .B(AES_CORE_DATAPATH__abc_15863_new_n5656_), .C(AES_CORE_DATAPATH__abc_15863_new_n5652_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5657_));
NAND3X1 NAND3X1_384 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5634_), .B(AES_CORE_DATAPATH__abc_15863_new_n5666_), .C(AES_CORE_DATAPATH__abc_15863_new_n5665_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5667_));
NAND3X1 NAND3X1_385 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3037_), .B(AES_CORE_DATAPATH__abc_15863_new_n3039_), .C(AES_CORE_DATAPATH__abc_15863_new_n3723_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5675_));
NAND3X1 NAND3X1_386 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5679_), .B(AES_CORE_DATAPATH__abc_15863_new_n5690_), .C(AES_CORE_DATAPATH__abc_15863_new_n5677_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5691_));
NAND3X1 NAND3X1_387 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5673_), .B(AES_CORE_DATAPATH__abc_15863_new_n5705_), .C(AES_CORE_DATAPATH__abc_15863_new_n5703_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5706_));
NAND3X1 NAND3X1_388 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5715_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5714_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5716_));
NAND3X1 NAND3X1_389 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5717_), .B(AES_CORE_DATAPATH__abc_15863_new_n5725_), .C(AES_CORE_DATAPATH__abc_15863_new_n5716_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5726_));
NAND3X1 NAND3X1_39 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2823_));
NAND3X1 NAND3X1_390 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5729_), .B(AES_CORE_DATAPATH__abc_15863_new_n5731_), .C(AES_CORE_DATAPATH__abc_15863_new_n5727_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5732_));
NAND3X1 NAND3X1_391 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5712_), .B(AES_CORE_DATAPATH__abc_15863_new_n5741_), .C(AES_CORE_DATAPATH__abc_15863_new_n5740_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5742_));
NAND3X1 NAND3X1_392 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5751_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .C(AES_CORE_DATAPATH__abc_15863_new_n5750_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5752_));
NAND3X1 NAND3X1_393 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5753_), .B(AES_CORE_DATAPATH__abc_15863_new_n5764_), .C(AES_CORE_DATAPATH__abc_15863_new_n5752_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5765_));
NAND3X1 NAND3X1_394 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5768_), .B(AES_CORE_DATAPATH__abc_15863_new_n5770_), .C(AES_CORE_DATAPATH__abc_15863_new_n5766_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5771_));
NAND3X1 NAND3X1_395 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5748_), .B(AES_CORE_DATAPATH__abc_15863_new_n5780_), .C(AES_CORE_DATAPATH__abc_15863_new_n5779_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5781_));
NAND3X1 NAND3X1_396 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3064_), .B(AES_CORE_DATAPATH__abc_15863_new_n3068_), .C(AES_CORE_DATAPATH__abc_15863_new_n3789_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5789_));
NAND3X1 NAND3X1_397 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5793_), .B(AES_CORE_DATAPATH__abc_15863_new_n5804_), .C(AES_CORE_DATAPATH__abc_15863_new_n5791_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5805_));
NAND3X1 NAND3X1_398 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5787_), .B(AES_CORE_DATAPATH__abc_15863_new_n5819_), .C(AES_CORE_DATAPATH__abc_15863_new_n5817_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5820_));
NAND3X1 NAND3X1_399 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4586_), .B(AES_CORE_DATAPATH__abc_15863_new_n6054_), .C(AES_CORE_DATAPATH__abc_15863_new_n4629_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6055_));
NAND3X1 NAND3X1_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n99_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n100_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n96_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_2_));
NAND3X1 NAND3X1_40 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2822_), .B(AES_CORE_DATAPATH__abc_15863_new_n2823_), .C(AES_CORE_DATAPATH__abc_15863_new_n2824_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2825_));
NAND3X1 NAND3X1_400 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4668_), .B(AES_CORE_DATAPATH__abc_15863_new_n6061_), .C(AES_CORE_DATAPATH__abc_15863_new_n4667_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6062_));
NAND3X1 NAND3X1_401 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4707_), .B(AES_CORE_DATAPATH__abc_15863_new_n6068_), .C(AES_CORE_DATAPATH__abc_15863_new_n4706_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6069_));
NAND3X1 NAND3X1_402 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4747_), .B(AES_CORE_DATAPATH__abc_15863_new_n6075_), .C(AES_CORE_DATAPATH__abc_15863_new_n4744_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6076_));
NAND3X1 NAND3X1_403 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4783_), .B(AES_CORE_DATAPATH__abc_15863_new_n6082_), .C(AES_CORE_DATAPATH__abc_15863_new_n4782_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6083_));
NAND3X1 NAND3X1_404 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4822_), .B(AES_CORE_DATAPATH__abc_15863_new_n6089_), .C(AES_CORE_DATAPATH__abc_15863_new_n4821_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6090_));
NAND3X1 NAND3X1_405 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4857_), .B(AES_CORE_DATAPATH__abc_15863_new_n6096_), .C(AES_CORE_DATAPATH__abc_15863_new_n4856_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6097_));
NAND3X1 NAND3X1_406 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4896_), .B(AES_CORE_DATAPATH__abc_15863_new_n6103_), .C(AES_CORE_DATAPATH__abc_15863_new_n4895_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6104_));
NAND3X1 NAND3X1_407 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4931_), .B(AES_CORE_DATAPATH__abc_15863_new_n6110_), .C(AES_CORE_DATAPATH__abc_15863_new_n4930_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6111_));
NAND3X1 NAND3X1_408 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4970_), .B(AES_CORE_DATAPATH__abc_15863_new_n6117_), .C(AES_CORE_DATAPATH__abc_15863_new_n4968_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6118_));
NAND3X1 NAND3X1_409 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5009_), .B(AES_CORE_DATAPATH__abc_15863_new_n6124_), .C(AES_CORE_DATAPATH__abc_15863_new_n5008_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6125_));
NAND3X1 NAND3X1_41 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2834_));
NAND3X1 NAND3X1_410 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5048_), .B(AES_CORE_DATAPATH__abc_15863_new_n6131_), .C(AES_CORE_DATAPATH__abc_15863_new_n5046_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6132_));
NAND3X1 NAND3X1_411 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5087_), .B(AES_CORE_DATAPATH__abc_15863_new_n6138_), .C(AES_CORE_DATAPATH__abc_15863_new_n5086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6139_));
NAND3X1 NAND3X1_412 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5126_), .B(AES_CORE_DATAPATH__abc_15863_new_n6145_), .C(AES_CORE_DATAPATH__abc_15863_new_n5124_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6146_));
NAND3X1 NAND3X1_413 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5162_), .B(AES_CORE_DATAPATH__abc_15863_new_n6152_), .C(AES_CORE_DATAPATH__abc_15863_new_n5161_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6153_));
NAND3X1 NAND3X1_414 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5201_), .B(AES_CORE_DATAPATH__abc_15863_new_n6159_), .C(AES_CORE_DATAPATH__abc_15863_new_n5199_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6160_));
NAND3X1 NAND3X1_415 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5240_), .B(AES_CORE_DATAPATH__abc_15863_new_n6166_), .C(AES_CORE_DATAPATH__abc_15863_new_n5239_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6167_));
NAND3X1 NAND3X1_416 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5279_), .B(AES_CORE_DATAPATH__abc_15863_new_n6173_), .C(AES_CORE_DATAPATH__abc_15863_new_n5277_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6174_));
NAND3X1 NAND3X1_417 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5318_), .B(AES_CORE_DATAPATH__abc_15863_new_n6180_), .C(AES_CORE_DATAPATH__abc_15863_new_n5316_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6181_));
NAND3X1 NAND3X1_418 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5357_), .B(AES_CORE_DATAPATH__abc_15863_new_n6187_), .C(AES_CORE_DATAPATH__abc_15863_new_n5355_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6188_));
NAND3X1 NAND3X1_419 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5396_), .B(AES_CORE_DATAPATH__abc_15863_new_n6194_), .C(AES_CORE_DATAPATH__abc_15863_new_n5395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6195_));
NAND3X1 NAND3X1_42 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2835_));
NAND3X1 NAND3X1_420 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5435_), .B(AES_CORE_DATAPATH__abc_15863_new_n6201_), .C(AES_CORE_DATAPATH__abc_15863_new_n5433_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6202_));
NAND3X1 NAND3X1_421 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5471_), .B(AES_CORE_DATAPATH__abc_15863_new_n6208_), .C(AES_CORE_DATAPATH__abc_15863_new_n5470_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6209_));
NAND3X1 NAND3X1_422 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5510_), .B(AES_CORE_DATAPATH__abc_15863_new_n6215_), .C(AES_CORE_DATAPATH__abc_15863_new_n5509_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6216_));
NAND3X1 NAND3X1_423 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5549_), .B(AES_CORE_DATAPATH__abc_15863_new_n6222_), .C(AES_CORE_DATAPATH__abc_15863_new_n5548_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6223_));
NAND3X1 NAND3X1_424 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5588_), .B(AES_CORE_DATAPATH__abc_15863_new_n6229_), .C(AES_CORE_DATAPATH__abc_15863_new_n5586_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6230_));
NAND3X1 NAND3X1_425 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5627_), .B(AES_CORE_DATAPATH__abc_15863_new_n6236_), .C(AES_CORE_DATAPATH__abc_15863_new_n5625_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6237_));
NAND3X1 NAND3X1_426 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5666_), .B(AES_CORE_DATAPATH__abc_15863_new_n6243_), .C(AES_CORE_DATAPATH__abc_15863_new_n5665_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6244_));
NAND3X1 NAND3X1_427 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5705_), .B(AES_CORE_DATAPATH__abc_15863_new_n6250_), .C(AES_CORE_DATAPATH__abc_15863_new_n5703_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6251_));
NAND3X1 NAND3X1_428 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5741_), .B(AES_CORE_DATAPATH__abc_15863_new_n6257_), .C(AES_CORE_DATAPATH__abc_15863_new_n5740_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6258_));
NAND3X1 NAND3X1_429 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5780_), .B(AES_CORE_DATAPATH__abc_15863_new_n6264_), .C(AES_CORE_DATAPATH__abc_15863_new_n5779_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6265_));
NAND3X1 NAND3X1_43 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2834_), .B(AES_CORE_DATAPATH__abc_15863_new_n2835_), .C(AES_CORE_DATAPATH__abc_15863_new_n2836_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2837_));
NAND3X1 NAND3X1_430 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5819_), .B(AES_CORE_DATAPATH__abc_15863_new_n6271_), .C(AES_CORE_DATAPATH__abc_15863_new_n5817_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6272_));
NAND3X1 NAND3X1_431 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4586_), .B(AES_CORE_DATAPATH__abc_15863_new_n6278_), .C(AES_CORE_DATAPATH__abc_15863_new_n4629_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6279_));
NAND3X1 NAND3X1_432 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4668_), .B(AES_CORE_DATAPATH__abc_15863_new_n6285_), .C(AES_CORE_DATAPATH__abc_15863_new_n4667_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6286_));
NAND3X1 NAND3X1_433 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4707_), .B(AES_CORE_DATAPATH__abc_15863_new_n6292_), .C(AES_CORE_DATAPATH__abc_15863_new_n4706_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6293_));
NAND3X1 NAND3X1_434 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4747_), .B(AES_CORE_DATAPATH__abc_15863_new_n6299_), .C(AES_CORE_DATAPATH__abc_15863_new_n4744_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6300_));
NAND3X1 NAND3X1_435 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4783_), .B(AES_CORE_DATAPATH__abc_15863_new_n6306_), .C(AES_CORE_DATAPATH__abc_15863_new_n4782_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6307_));
NAND3X1 NAND3X1_436 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4822_), .B(AES_CORE_DATAPATH__abc_15863_new_n6313_), .C(AES_CORE_DATAPATH__abc_15863_new_n4821_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6314_));
NAND3X1 NAND3X1_437 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4857_), .B(AES_CORE_DATAPATH__abc_15863_new_n6320_), .C(AES_CORE_DATAPATH__abc_15863_new_n4856_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6321_));
NAND3X1 NAND3X1_438 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4896_), .B(AES_CORE_DATAPATH__abc_15863_new_n6327_), .C(AES_CORE_DATAPATH__abc_15863_new_n4895_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6328_));
NAND3X1 NAND3X1_439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4931_), .B(AES_CORE_DATAPATH__abc_15863_new_n6334_), .C(AES_CORE_DATAPATH__abc_15863_new_n4930_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6335_));
NAND3X1 NAND3X1_44 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2845_));
NAND3X1 NAND3X1_440 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4970_), .B(AES_CORE_DATAPATH__abc_15863_new_n6341_), .C(AES_CORE_DATAPATH__abc_15863_new_n4968_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6342_));
NAND3X1 NAND3X1_441 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5009_), .B(AES_CORE_DATAPATH__abc_15863_new_n6348_), .C(AES_CORE_DATAPATH__abc_15863_new_n5008_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6349_));
NAND3X1 NAND3X1_442 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5048_), .B(AES_CORE_DATAPATH__abc_15863_new_n6355_), .C(AES_CORE_DATAPATH__abc_15863_new_n5046_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6356_));
NAND3X1 NAND3X1_443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5087_), .B(AES_CORE_DATAPATH__abc_15863_new_n6362_), .C(AES_CORE_DATAPATH__abc_15863_new_n5086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6363_));
NAND3X1 NAND3X1_444 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5126_), .B(AES_CORE_DATAPATH__abc_15863_new_n6369_), .C(AES_CORE_DATAPATH__abc_15863_new_n5124_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6370_));
NAND3X1 NAND3X1_445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5162_), .B(AES_CORE_DATAPATH__abc_15863_new_n6376_), .C(AES_CORE_DATAPATH__abc_15863_new_n5161_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6377_));
NAND3X1 NAND3X1_446 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5201_), .B(AES_CORE_DATAPATH__abc_15863_new_n6383_), .C(AES_CORE_DATAPATH__abc_15863_new_n5199_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6384_));
NAND3X1 NAND3X1_447 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5240_), .B(AES_CORE_DATAPATH__abc_15863_new_n6390_), .C(AES_CORE_DATAPATH__abc_15863_new_n5239_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6391_));
NAND3X1 NAND3X1_448 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5279_), .B(AES_CORE_DATAPATH__abc_15863_new_n6397_), .C(AES_CORE_DATAPATH__abc_15863_new_n5277_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6398_));
NAND3X1 NAND3X1_449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5318_), .B(AES_CORE_DATAPATH__abc_15863_new_n6404_), .C(AES_CORE_DATAPATH__abc_15863_new_n5316_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6405_));
NAND3X1 NAND3X1_45 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2846_));
NAND3X1 NAND3X1_450 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5357_), .B(AES_CORE_DATAPATH__abc_15863_new_n6411_), .C(AES_CORE_DATAPATH__abc_15863_new_n5355_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6412_));
NAND3X1 NAND3X1_451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5396_), .B(AES_CORE_DATAPATH__abc_15863_new_n6418_), .C(AES_CORE_DATAPATH__abc_15863_new_n5395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6419_));
NAND3X1 NAND3X1_452 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5435_), .B(AES_CORE_DATAPATH__abc_15863_new_n6425_), .C(AES_CORE_DATAPATH__abc_15863_new_n5433_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6426_));
NAND3X1 NAND3X1_453 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5471_), .B(AES_CORE_DATAPATH__abc_15863_new_n6432_), .C(AES_CORE_DATAPATH__abc_15863_new_n5470_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6433_));
NAND3X1 NAND3X1_454 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5510_), .B(AES_CORE_DATAPATH__abc_15863_new_n6439_), .C(AES_CORE_DATAPATH__abc_15863_new_n5509_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6440_));
NAND3X1 NAND3X1_455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5549_), .B(AES_CORE_DATAPATH__abc_15863_new_n6446_), .C(AES_CORE_DATAPATH__abc_15863_new_n5548_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6447_));
NAND3X1 NAND3X1_456 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5588_), .B(AES_CORE_DATAPATH__abc_15863_new_n6453_), .C(AES_CORE_DATAPATH__abc_15863_new_n5586_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6454_));
NAND3X1 NAND3X1_457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5627_), .B(AES_CORE_DATAPATH__abc_15863_new_n6460_), .C(AES_CORE_DATAPATH__abc_15863_new_n5625_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6461_));
NAND3X1 NAND3X1_458 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5666_), .B(AES_CORE_DATAPATH__abc_15863_new_n6467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5665_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6468_));
NAND3X1 NAND3X1_459 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5705_), .B(AES_CORE_DATAPATH__abc_15863_new_n6474_), .C(AES_CORE_DATAPATH__abc_15863_new_n5703_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6475_));
NAND3X1 NAND3X1_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2845_), .B(AES_CORE_DATAPATH__abc_15863_new_n2846_), .C(AES_CORE_DATAPATH__abc_15863_new_n2847_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2848_));
NAND3X1 NAND3X1_460 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5741_), .B(AES_CORE_DATAPATH__abc_15863_new_n6481_), .C(AES_CORE_DATAPATH__abc_15863_new_n5740_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6482_));
NAND3X1 NAND3X1_461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5780_), .B(AES_CORE_DATAPATH__abc_15863_new_n6488_), .C(AES_CORE_DATAPATH__abc_15863_new_n5779_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6489_));
NAND3X1 NAND3X1_462 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5819_), .B(AES_CORE_DATAPATH__abc_15863_new_n6495_), .C(AES_CORE_DATAPATH__abc_15863_new_n5817_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6496_));
NAND3X1 NAND3X1_463 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4586_), .B(AES_CORE_DATAPATH__abc_15863_new_n6503_), .C(AES_CORE_DATAPATH__abc_15863_new_n4629_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6504_));
NAND3X1 NAND3X1_464 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4668_), .B(AES_CORE_DATAPATH__abc_15863_new_n6509_), .C(AES_CORE_DATAPATH__abc_15863_new_n4667_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6510_));
NAND3X1 NAND3X1_465 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4707_), .B(AES_CORE_DATAPATH__abc_15863_new_n6516_), .C(AES_CORE_DATAPATH__abc_15863_new_n4706_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6517_));
NAND3X1 NAND3X1_466 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4747_), .B(AES_CORE_DATAPATH__abc_15863_new_n6522_), .C(AES_CORE_DATAPATH__abc_15863_new_n4744_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6523_));
NAND3X1 NAND3X1_467 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4783_), .B(AES_CORE_DATAPATH__abc_15863_new_n6529_), .C(AES_CORE_DATAPATH__abc_15863_new_n4782_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6530_));
NAND3X1 NAND3X1_468 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4822_), .B(AES_CORE_DATAPATH__abc_15863_new_n6536_), .C(AES_CORE_DATAPATH__abc_15863_new_n4821_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6537_));
NAND3X1 NAND3X1_469 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4857_), .B(AES_CORE_DATAPATH__abc_15863_new_n6543_), .C(AES_CORE_DATAPATH__abc_15863_new_n4856_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6544_));
NAND3X1 NAND3X1_47 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2854_));
NAND3X1 NAND3X1_470 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4896_), .B(AES_CORE_DATAPATH__abc_15863_new_n6549_), .C(AES_CORE_DATAPATH__abc_15863_new_n4895_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6550_));
NAND3X1 NAND3X1_471 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4931_), .B(AES_CORE_DATAPATH__abc_15863_new_n6556_), .C(AES_CORE_DATAPATH__abc_15863_new_n4930_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6557_));
NAND3X1 NAND3X1_472 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4970_), .B(AES_CORE_DATAPATH__abc_15863_new_n6562_), .C(AES_CORE_DATAPATH__abc_15863_new_n4968_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6563_));
NAND3X1 NAND3X1_473 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5009_), .B(AES_CORE_DATAPATH__abc_15863_new_n6569_), .C(AES_CORE_DATAPATH__abc_15863_new_n5008_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6570_));
NAND3X1 NAND3X1_474 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5048_), .B(AES_CORE_DATAPATH__abc_15863_new_n6575_), .C(AES_CORE_DATAPATH__abc_15863_new_n5046_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6576_));
NAND3X1 NAND3X1_475 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5087_), .B(AES_CORE_DATAPATH__abc_15863_new_n6582_), .C(AES_CORE_DATAPATH__abc_15863_new_n5086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6583_));
NAND3X1 NAND3X1_476 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5126_), .B(AES_CORE_DATAPATH__abc_15863_new_n6588_), .C(AES_CORE_DATAPATH__abc_15863_new_n5124_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6589_));
NAND3X1 NAND3X1_477 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5162_), .B(AES_CORE_DATAPATH__abc_15863_new_n6595_), .C(AES_CORE_DATAPATH__abc_15863_new_n5161_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6596_));
NAND3X1 NAND3X1_478 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5201_), .B(AES_CORE_DATAPATH__abc_15863_new_n6601_), .C(AES_CORE_DATAPATH__abc_15863_new_n5199_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6602_));
NAND3X1 NAND3X1_479 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5240_), .B(AES_CORE_DATAPATH__abc_15863_new_n6608_), .C(AES_CORE_DATAPATH__abc_15863_new_n5239_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6609_));
NAND3X1 NAND3X1_48 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2855_));
NAND3X1 NAND3X1_480 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5279_), .B(AES_CORE_DATAPATH__abc_15863_new_n6614_), .C(AES_CORE_DATAPATH__abc_15863_new_n5277_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6615_));
NAND3X1 NAND3X1_481 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5318_), .B(AES_CORE_DATAPATH__abc_15863_new_n6620_), .C(AES_CORE_DATAPATH__abc_15863_new_n5316_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6621_));
NAND3X1 NAND3X1_482 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5357_), .B(AES_CORE_DATAPATH__abc_15863_new_n6626_), .C(AES_CORE_DATAPATH__abc_15863_new_n5355_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6627_));
NAND3X1 NAND3X1_483 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5396_), .B(AES_CORE_DATAPATH__abc_15863_new_n6633_), .C(AES_CORE_DATAPATH__abc_15863_new_n5395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6634_));
NAND3X1 NAND3X1_484 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5435_), .B(AES_CORE_DATAPATH__abc_15863_new_n6639_), .C(AES_CORE_DATAPATH__abc_15863_new_n5433_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6640_));
NAND3X1 NAND3X1_485 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5471_), .B(AES_CORE_DATAPATH__abc_15863_new_n6646_), .C(AES_CORE_DATAPATH__abc_15863_new_n5470_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6647_));
NAND3X1 NAND3X1_486 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5510_), .B(AES_CORE_DATAPATH__abc_15863_new_n6652_), .C(AES_CORE_DATAPATH__abc_15863_new_n5509_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6653_));
NAND3X1 NAND3X1_487 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5549_), .B(AES_CORE_DATAPATH__abc_15863_new_n6659_), .C(AES_CORE_DATAPATH__abc_15863_new_n5548_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6660_));
NAND3X1 NAND3X1_488 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5588_), .B(AES_CORE_DATAPATH__abc_15863_new_n6665_), .C(AES_CORE_DATAPATH__abc_15863_new_n5586_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6666_));
NAND3X1 NAND3X1_489 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5627_), .B(AES_CORE_DATAPATH__abc_15863_new_n6671_), .C(AES_CORE_DATAPATH__abc_15863_new_n5625_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6672_));
NAND3X1 NAND3X1_49 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2854_), .B(AES_CORE_DATAPATH__abc_15863_new_n2855_), .C(AES_CORE_DATAPATH__abc_15863_new_n2856_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2857_));
NAND3X1 NAND3X1_490 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5666_), .B(AES_CORE_DATAPATH__abc_15863_new_n6678_), .C(AES_CORE_DATAPATH__abc_15863_new_n5665_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6679_));
NAND3X1 NAND3X1_491 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5705_), .B(AES_CORE_DATAPATH__abc_15863_new_n6684_), .C(AES_CORE_DATAPATH__abc_15863_new_n5703_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6685_));
NAND3X1 NAND3X1_492 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5741_), .B(AES_CORE_DATAPATH__abc_15863_new_n6691_), .C(AES_CORE_DATAPATH__abc_15863_new_n5740_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6692_));
NAND3X1 NAND3X1_493 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5780_), .B(AES_CORE_DATAPATH__abc_15863_new_n6698_), .C(AES_CORE_DATAPATH__abc_15863_new_n5779_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6699_));
NAND3X1 NAND3X1_494 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5819_), .B(AES_CORE_DATAPATH__abc_15863_new_n6704_), .C(AES_CORE_DATAPATH__abc_15863_new_n5817_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6705_));
NAND3X1 NAND3X1_495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6981_), .B(AES_CORE_DATAPATH__abc_15863_new_n7061_), .C(AES_CORE_DATAPATH__abc_15863_new_n7060_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7062_));
NAND3X1 NAND3X1_496 ( .A(AES_CORE_DATAPATH_iv_3__17_), .B(AES_CORE_DATAPATH_iv_3__18_), .C(AES_CORE_DATAPATH__abc_15863_new_n7085_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7097_));
NAND3X1 NAND3X1_497 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6981_), .B(AES_CORE_DATAPATH__abc_15863_new_n7096_), .C(AES_CORE_DATAPATH__abc_15863_new_n7097_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7098_));
NAND3X1 NAND3X1_498 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7109_), .B(AES_CORE_DATAPATH__abc_15863_new_n7110_), .C(AES_CORE_DATAPATH__abc_15863_new_n7108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7111_));
NAND3X1 NAND3X1_499 ( .A(AES_CORE_DATAPATH_iv_3__26_), .B(AES_CORE_DATAPATH_iv_3__27_), .C(AES_CORE_DATAPATH__abc_15863_new_n7163_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7179_));
NAND3X1 NAND3X1_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n126_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n169_), .Y(AES_CORE_CONTROL_UNIT_col_en_0_));
NAND3X1 NAND3X1_50 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2864_));
NAND3X1 NAND3X1_500 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n419_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n417_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n420_));
NAND3X1 NAND3X1_501 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n420_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n428_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n429_));
NAND3X1 NAND3X1_502 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n434_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n435_));
NAND3X1 NAND3X1_503 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n437_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n435_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n438_));
NAND3X1 NAND3X1_504 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n433_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n438_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n442_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n443_));
NAND3X1 NAND3X1_505 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n400_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n401_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n445_));
NAND3X1 NAND3X1_506 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n432_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n449_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n450_));
NAND3X1 NAND3X1_507 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n438_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n442_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n451_));
NAND3X1 NAND3X1_508 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n451_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n452_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n453_));
NAND3X1 NAND3X1_509 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n461_));
NAND3X1 NAND3X1_51 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2865_));
NAND3X1 NAND3X1_510 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n462_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n461_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n463_));
NAND3X1 NAND3X1_511 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n458_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n463_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n460_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n464_));
NAND3X1 NAND3X1_512 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n457_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n468_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n469_));
NAND3X1 NAND3X1_513 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n463_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n460_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n470_));
NAND3X1 NAND3X1_514 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n470_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n471_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n472_));
NAND3X1 NAND3X1_515 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n476_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n477_));
NAND3X1 NAND3X1_516 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n424_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n436_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n478_));
NAND3X1 NAND3X1_517 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n480_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n486_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n487_));
NAND3X1 NAND3X1_518 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n489_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n490_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n491_));
NAND3X1 NAND3X1_519 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n437_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n478_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n496_));
NAND3X1 NAND3X1_52 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2864_), .B(AES_CORE_DATAPATH__abc_15863_new_n2865_), .C(AES_CORE_DATAPATH__abc_15863_new_n2866_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2867_));
NAND3X1 NAND3X1_520 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n495_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n496_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n497_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n498_));
NAND3X1 NAND3X1_521 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n494_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n501_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n502_));
NAND3X1 NAND3X1_522 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n496_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n497_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n503_));
NAND3X1 NAND3X1_523 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n503_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n504_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n505_));
NAND3X1 NAND3X1_524 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n510_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n511_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n512_));
NAND3X1 NAND3X1_525 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n512_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n515_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n516_));
NAND3X1 NAND3X1_526 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n520_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n519_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n521_));
NAND3X1 NAND3X1_527 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n521_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n524_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n525_));
NAND3X1 NAND3X1_528 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n443_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n448_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n682_));
NAND3X1 NAND3X1_529 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n498_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n500_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n688_));
NAND3X1 NAND3X1_53 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2876_));
NAND3X1 NAND3X1_530 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n138_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n143_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n146_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n147_));
NAND3X1 NAND3X1_531 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n127_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n147_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n153_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n154_));
NAND3X1 NAND3X1_532 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n150_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n143_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n146_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n156_));
NAND3X1 NAND3X1_533 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n156_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n155_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n157_));
NAND3X1 NAND3X1_534 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n169_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n183_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n186_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n187_));
NAND3X1 NAND3X1_535 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n190_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n192_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n191_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n193_));
NAND3X1 NAND3X1_536 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n205_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n208_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n209_));
NAND3X1 NAND3X1_537 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n210_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n211_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n212_));
NAND3X1 NAND3X1_538 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n223_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n209_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n212_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n224_));
NAND3X1 NAND3X1_539 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n210_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n211_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n225_));
NAND3X1 NAND3X1_54 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2877_));
NAND3X1 NAND3X1_540 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n205_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n208_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n226_));
NAND3X1 NAND3X1_541 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n222_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n225_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n226_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n227_));
NAND3X1 NAND3X1_542 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n201_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n224_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n227_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n228_));
NAND3X1 NAND3X1_543 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n222_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n209_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n212_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n229_));
NAND3X1 NAND3X1_544 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n223_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n225_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n226_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n230_));
NAND3X1 NAND3X1_545 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n229_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n230_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n231_));
NAND3X1 NAND3X1_546 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n266_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n275_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n276_));
NAND3X1 NAND3X1_547 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n244_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n276_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n261_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n277_));
NAND3X1 NAND3X1_548 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n266_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n275_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n281_));
NAND3X1 NAND3X1_549 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n280_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n281_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n282_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n283_));
NAND3X1 NAND3X1_55 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2876_), .B(AES_CORE_DATAPATH__abc_15863_new_n2877_), .C(AES_CORE_DATAPATH__abc_15863_new_n2878_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2879_));
NAND3X1 NAND3X1_550 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n277_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n283_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n284_));
NAND3X1 NAND3X1_551 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n244_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n281_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n282_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n286_));
NAND3X1 NAND3X1_552 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n280_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n276_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n261_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n287_));
NAND3X1 NAND3X1_553 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n285_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n286_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n287_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n288_));
NAND3X1 NAND3X1_554 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n300_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n301_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n280_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n302_));
NAND3X1 NAND3X1_555 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n298_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n309_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n310_));
NAND3X1 NAND3X1_556 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n300_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n301_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n244_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n315_));
NAND3X1 NAND3X1_557 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n313_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n314_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n315_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n316_));
NAND3X1 NAND3X1_558 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n292_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n310_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n316_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n317_));
NAND3X1 NAND3X1_559 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n331_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n329_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n332_));
NAND3X1 NAND3X1_56 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2884_));
NAND3X1 NAND3X1_560 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n333_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n335_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n334_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n336_));
NAND3X1 NAND3X1_561 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n332_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n336_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n326_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n337_));
NAND3X1 NAND3X1_562 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n333_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n331_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n329_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n338_));
NAND3X1 NAND3X1_563 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n335_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n334_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n339_));
NAND3X1 NAND3X1_564 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n338_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n339_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n340_));
NAND3X1 NAND3X1_565 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n119_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n113_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n364_));
NAND3X1 NAND3X1_566 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n364_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n368_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n369_));
NAND3X1 NAND3X1_567 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n374_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n192_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n191_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n375_));
NAND3X1 NAND3X1_568 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n376_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n183_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n186_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n377_));
NAND3X1 NAND3X1_569 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n259_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n209_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n212_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n389_));
NAND3X1 NAND3X1_57 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2885_));
NAND3X1 NAND3X1_570 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n274_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n225_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n226_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n390_));
NAND3X1 NAND3X1_571 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n384_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n389_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n390_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n391_));
NAND3X1 NAND3X1_572 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n276_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n398_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n261_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n399_));
NAND3X1 NAND3X1_573 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n281_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n400_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n282_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n401_));
NAND3X1 NAND3X1_574 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n397_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n399_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n401_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n402_));
NAND3X1 NAND3X1_575 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n276_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n400_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n261_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n403_));
NAND3X1 NAND3X1_576 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n281_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n398_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n282_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n404_));
NAND3X1 NAND3X1_577 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n403_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n404_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n405_));
NAND3X1 NAND3X1_578 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n328_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n314_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n315_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n412_));
NAND3X1 NAND3X1_579 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n330_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n309_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n413_));
NAND3X1 NAND3X1_58 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2884_), .B(AES_CORE_DATAPATH__abc_15863_new_n2885_), .C(AES_CORE_DATAPATH__abc_15863_new_n2886_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2887_));
NAND3X1 NAND3X1_580 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n411_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n412_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n413_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n414_));
NAND3X1 NAND3X1_581 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n328_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n309_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n415_));
NAND3X1 NAND3X1_582 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n330_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n314_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n315_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n416_));
NAND3X1 NAND3X1_583 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n415_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n416_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n417_));
NAND3X1 NAND3X1_584 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n423_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n331_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n329_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n424_));
NAND3X1 NAND3X1_585 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n349_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n335_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n334_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n425_));
NAND3X1 NAND3X1_586 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n423_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n335_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n334_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n427_));
NAND3X1 NAND3X1_587 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n349_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n331_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n329_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n428_));
NAND3X1 NAND3X1_588 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n147_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n445_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n153_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n446_));
NAND3X1 NAND3X1_589 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n156_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n155_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n447_));
NAND3X1 NAND3X1_59 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2896_));
NAND3X1 NAND3X1_590 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n456_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n224_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n227_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n457_));
NAND3X1 NAND3X1_591 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n229_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n230_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n458_));
NAND3X1 NAND3X1_592 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n277_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n283_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n464_));
NAND3X1 NAND3X1_593 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n465_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n286_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n287_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n466_));
NAND3X1 NAND3X1_594 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n469_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n310_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n316_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n471_));
NAND3X1 NAND3X1_595 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n476_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n332_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n336_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n478_));
NAND3X1 NAND3X1_596 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n338_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n339_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n479_));
NAND3X1 NAND3X1_597 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n364_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n368_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n494_));
NAND3X1 NAND3X1_598 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n502_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n389_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n390_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n504_));
NAND3X1 NAND3X1_599 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n510_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n399_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n401_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n511_));
NAND3X1 NAND3X1_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n169_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_), .Y(AES_CORE_CONTROL_UNIT_col_en_1_));
NAND3X1 NAND3X1_60 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2897_));
NAND3X1 NAND3X1_600 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n403_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n404_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n512_));
NAND3X1 NAND3X1_601 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n516_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n412_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n413_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n518_));
NAND3X1 NAND3X1_602 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n415_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n416_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n519_));
NAND3X1 NAND3X1_603 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n61_));
NAND3X1 NAND3X1_604 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n65_));
NAND3X1 NAND3X1_605 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n77_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n109_));
NAND3X1 NAND3X1_606 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n111_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n112_));
NAND3X1 NAND3X1_607 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n112_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n109_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n113_));
NAND3X1 NAND3X1_608 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n114_));
NAND3X1 NAND3X1_609 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n115_));
NAND3X1 NAND3X1_61 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2896_), .B(AES_CORE_DATAPATH__abc_15863_new_n2897_), .C(AES_CORE_DATAPATH__abc_15863_new_n2898_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2899_));
NAND3X1 NAND3X1_610 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n114_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n116_));
NAND3X1 NAND3X1_611 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n116_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n118_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n119_));
NAND3X1 NAND3X1_612 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n130_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n133_));
NAND3X1 NAND3X1_613 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n144_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n148_));
NAND3X1 NAND3X1_614 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n148_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n143_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n149_));
NAND3X1 NAND3X1_615 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n164_));
NAND3X1 NAND3X1_616 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n169_));
NAND3X1 NAND3X1_617 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_));
NAND3X1 NAND3X1_618 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n178_));
NAND3X1 NAND3X1_619 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n142_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n181_));
NAND3X1 NAND3X1_62 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2907_));
NAND3X1 NAND3X1_620 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n182_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n183_));
NAND3X1 NAND3X1_621 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_));
NAND3X1 NAND3X1_622 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n156_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n198_));
NAND3X1 NAND3X1_623 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n198_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n183_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n178_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n199_));
NAND3X1 NAND3X1_624 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n207_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n211_));
NAND3X1 NAND3X1_625 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n219_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n222_));
NAND3X1 NAND3X1_626 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n235_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n236_));
NAND3X1 NAND3X1_627 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n238_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n239_));
NAND3X1 NAND3X1_628 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n255_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n256_));
NAND3X1 NAND3X1_629 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n257_));
NAND3X1 NAND3X1_63 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2908_));
NAND3X1 NAND3X1_630 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n194_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n259_));
NAND3X1 NAND3X1_631 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n263_));
NAND3X1 NAND3X1_632 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n267_));
NAND3X1 NAND3X1_633 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n269_));
NAND3X1 NAND3X1_634 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n272_));
NAND3X1 NAND3X1_635 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n273_));
NAND3X1 NAND3X1_636 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n238_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n296_));
NAND3X1 NAND3X1_637 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n297_));
NAND3X1 NAND3X1_638 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n230_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n298_));
NAND3X1 NAND3X1_639 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n298_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n296_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n299_));
NAND3X1 NAND3X1_64 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2907_), .B(AES_CORE_DATAPATH__abc_15863_new_n2908_), .C(AES_CORE_DATAPATH__abc_15863_new_n2909_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2910_));
NAND3X1 NAND3X1_640 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n315_));
NAND3X1 NAND3X1_641 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n318_));
NAND3X1 NAND3X1_642 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n318_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n320_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n321_));
NAND3X1 NAND3X1_643 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n322_));
NAND3X1 NAND3X1_644 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n323_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n324_));
NAND3X1 NAND3X1_645 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n308_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n340_));
NAND3X1 NAND3X1_646 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n341_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n342_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n344_));
NAND3X1 NAND3X1_647 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n320_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n348_));
NAND3X1 NAND3X1_648 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n323_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n349_));
NAND3X1 NAND3X1_649 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n334_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n352_));
NAND3X1 NAND3X1_65 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2916_));
NAND3X1 NAND3X1_650 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n354_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n356_));
NAND3X1 NAND3X1_651 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n357_));
NAND3X1 NAND3X1_652 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n358_));
NAND3X1 NAND3X1_653 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n359_));
NAND3X1 NAND3X1_654 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n360_));
NAND3X1 NAND3X1_655 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n361_));
NAND3X1 NAND3X1_656 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n319_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n362_));
NAND3X1 NAND3X1_657 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n365_));
NAND3X1 NAND3X1_658 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n366_));
NAND3X1 NAND3X1_659 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n377_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n378_));
NAND3X1 NAND3X1_66 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2917_));
NAND3X1 NAND3X1_660 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n381_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n383_));
NAND3X1 NAND3X1_661 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n386_));
NAND3X1 NAND3X1_662 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n91_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n389_));
NAND3X1 NAND3X1_663 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n390_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n391_));
NAND3X1 NAND3X1_664 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n392_));
NAND3X1 NAND3X1_665 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n408_));
NAND3X1 NAND3X1_666 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n409_));
NAND3X1 NAND3X1_667 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n423_));
NAND3X1 NAND3X1_668 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n424_));
NAND3X1 NAND3X1_669 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n424_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n426_));
NAND3X1 NAND3X1_67 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2916_), .B(AES_CORE_DATAPATH__abc_15863_new_n2917_), .C(AES_CORE_DATAPATH__abc_15863_new_n2918_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2919_));
NAND3X1 NAND3X1_670 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n427_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n431_));
NAND3X1 NAND3X1_671 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n434_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n435_));
NAND3X1 NAND3X1_672 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n392_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n437_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n438_));
NAND3X1 NAND3X1_673 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n438_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n439_));
NAND3X1 NAND3X1_674 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n440_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n441_));
NAND3X1 NAND3X1_675 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n423_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n443_));
NAND3X1 NAND3X1_676 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n442_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n447_));
NAND3X1 NAND3X1_677 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n446_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n452_));
NAND3X1 NAND3X1_678 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n444_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n453_));
NAND3X1 NAND3X1_679 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n453_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n452_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n454_));
NAND3X1 NAND3X1_68 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2926_));
NAND3X1 NAND3X1_680 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n459_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n458_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n413_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n460_));
NAND3X1 NAND3X1_681 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n463_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n464_));
NAND3X1 NAND3X1_682 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n457_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n465_));
NAND3X1 NAND3X1_683 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n462_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n468_));
NAND3X1 NAND3X1_684 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n468_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n470_));
NAND3X1 NAND3X1_685 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n470_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n465_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n471_));
NAND3X1 NAND3X1_686 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n472_));
NAND3X1 NAND3X1_687 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n457_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n473_));
NAND3X1 NAND3X1_688 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n473_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n474_));
NAND3X1 NAND3X1_689 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n477_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n480_));
NAND3X1 NAND3X1_69 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2927_));
NAND3X1 NAND3X1_690 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n479_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n481_));
NAND3X1 NAND3X1_691 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n478_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n483_));
NAND3X1 NAND3X1_692 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n483_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n484_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n485_));
NAND3X1 NAND3X1_693 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n451_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n481_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n486_));
NAND3X1 NAND3X1_694 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n483_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n484_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n487_));
NAND3X1 NAND3X1_695 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n480_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n488_));
NAND3X1 NAND3X1_696 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n488_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n489_));
NAND3X1 NAND3X1_697 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n383_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n498_));
NAND3X1 NAND3X1_698 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n61_));
NAND3X1 NAND3X1_699 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n65_));
NAND3X1 NAND3X1_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n169_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n176_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_), .Y(AES_CORE_CONTROL_UNIT_col_en_2_));
NAND3X1 NAND3X1_70 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2926_), .B(AES_CORE_DATAPATH__abc_15863_new_n2927_), .C(AES_CORE_DATAPATH__abc_15863_new_n2928_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2929_));
NAND3X1 NAND3X1_700 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n77_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n109_));
NAND3X1 NAND3X1_701 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n111_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n112_));
NAND3X1 NAND3X1_702 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n112_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n109_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n113_));
NAND3X1 NAND3X1_703 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n114_));
NAND3X1 NAND3X1_704 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n115_));
NAND3X1 NAND3X1_705 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n114_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n116_));
NAND3X1 NAND3X1_706 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n116_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n118_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n119_));
NAND3X1 NAND3X1_707 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n130_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n133_));
NAND3X1 NAND3X1_708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n144_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n148_));
NAND3X1 NAND3X1_709 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n148_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n143_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n149_));
NAND3X1 NAND3X1_71 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2936_));
NAND3X1 NAND3X1_710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n164_));
NAND3X1 NAND3X1_711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n169_));
NAND3X1 NAND3X1_712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_));
NAND3X1 NAND3X1_713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n178_));
NAND3X1 NAND3X1_714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n142_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n181_));
NAND3X1 NAND3X1_715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n182_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n183_));
NAND3X1 NAND3X1_716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_));
NAND3X1 NAND3X1_717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n156_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n198_));
NAND3X1 NAND3X1_718 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n198_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n183_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n178_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n199_));
NAND3X1 NAND3X1_719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n207_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n211_));
NAND3X1 NAND3X1_72 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2937_));
NAND3X1 NAND3X1_720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n219_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n222_));
NAND3X1 NAND3X1_721 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n235_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n236_));
NAND3X1 NAND3X1_722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n238_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n239_));
NAND3X1 NAND3X1_723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n255_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n256_));
NAND3X1 NAND3X1_724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n257_));
NAND3X1 NAND3X1_725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n194_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n259_));
NAND3X1 NAND3X1_726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n263_));
NAND3X1 NAND3X1_727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n267_));
NAND3X1 NAND3X1_728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n269_));
NAND3X1 NAND3X1_729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n272_));
NAND3X1 NAND3X1_73 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2936_), .B(AES_CORE_DATAPATH__abc_15863_new_n2937_), .C(AES_CORE_DATAPATH__abc_15863_new_n2938_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2939_));
NAND3X1 NAND3X1_730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n273_));
NAND3X1 NAND3X1_731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n238_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n296_));
NAND3X1 NAND3X1_732 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n297_));
NAND3X1 NAND3X1_733 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n230_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n298_));
NAND3X1 NAND3X1_734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n298_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n296_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n299_));
NAND3X1 NAND3X1_735 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n315_));
NAND3X1 NAND3X1_736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n318_));
NAND3X1 NAND3X1_737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n318_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n320_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n321_));
NAND3X1 NAND3X1_738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n322_));
NAND3X1 NAND3X1_739 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n323_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n324_));
NAND3X1 NAND3X1_74 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2947_));
NAND3X1 NAND3X1_740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n308_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n340_));
NAND3X1 NAND3X1_741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n341_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n342_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n344_));
NAND3X1 NAND3X1_742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n320_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n348_));
NAND3X1 NAND3X1_743 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n323_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n349_));
NAND3X1 NAND3X1_744 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n334_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n352_));
NAND3X1 NAND3X1_745 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n354_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n356_));
NAND3X1 NAND3X1_746 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n357_));
NAND3X1 NAND3X1_747 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n358_));
NAND3X1 NAND3X1_748 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n359_));
NAND3X1 NAND3X1_749 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n360_));
NAND3X1 NAND3X1_75 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2948_));
NAND3X1 NAND3X1_750 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n361_));
NAND3X1 NAND3X1_751 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n319_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n362_));
NAND3X1 NAND3X1_752 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n365_));
NAND3X1 NAND3X1_753 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n366_));
NAND3X1 NAND3X1_754 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n377_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n378_));
NAND3X1 NAND3X1_755 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n381_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n383_));
NAND3X1 NAND3X1_756 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n386_));
NAND3X1 NAND3X1_757 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n91_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n389_));
NAND3X1 NAND3X1_758 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n390_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n391_));
NAND3X1 NAND3X1_759 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n392_));
NAND3X1 NAND3X1_76 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2947_), .B(AES_CORE_DATAPATH__abc_15863_new_n2948_), .C(AES_CORE_DATAPATH__abc_15863_new_n2949_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2950_));
NAND3X1 NAND3X1_760 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n408_));
NAND3X1 NAND3X1_761 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n409_));
NAND3X1 NAND3X1_762 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n423_));
NAND3X1 NAND3X1_763 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n424_));
NAND3X1 NAND3X1_764 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n424_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n426_));
NAND3X1 NAND3X1_765 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n427_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n431_));
NAND3X1 NAND3X1_766 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n434_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n435_));
NAND3X1 NAND3X1_767 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n392_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n437_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n438_));
NAND3X1 NAND3X1_768 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n438_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n439_));
NAND3X1 NAND3X1_769 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n440_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n441_));
NAND3X1 NAND3X1_77 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2959_));
NAND3X1 NAND3X1_770 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n423_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n443_));
NAND3X1 NAND3X1_771 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n442_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n447_));
NAND3X1 NAND3X1_772 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n446_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n452_));
NAND3X1 NAND3X1_773 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n444_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n453_));
NAND3X1 NAND3X1_774 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n453_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n452_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n454_));
NAND3X1 NAND3X1_775 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n459_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n458_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n413_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n460_));
NAND3X1 NAND3X1_776 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n463_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n464_));
NAND3X1 NAND3X1_777 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n457_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n465_));
NAND3X1 NAND3X1_778 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n462_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n468_));
NAND3X1 NAND3X1_779 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n468_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n470_));
NAND3X1 NAND3X1_78 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2960_));
NAND3X1 NAND3X1_780 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n470_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n465_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n471_));
NAND3X1 NAND3X1_781 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n472_));
NAND3X1 NAND3X1_782 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n457_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n473_));
NAND3X1 NAND3X1_783 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n473_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n474_));
NAND3X1 NAND3X1_784 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n477_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n480_));
NAND3X1 NAND3X1_785 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n479_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n481_));
NAND3X1 NAND3X1_786 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n478_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n483_));
NAND3X1 NAND3X1_787 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n483_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n484_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n485_));
NAND3X1 NAND3X1_788 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n451_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n481_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n486_));
NAND3X1 NAND3X1_789 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n483_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n484_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n487_));
NAND3X1 NAND3X1_79 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2959_), .B(AES_CORE_DATAPATH__abc_15863_new_n2960_), .C(AES_CORE_DATAPATH__abc_15863_new_n2961_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2962_));
NAND3X1 NAND3X1_790 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n480_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n488_));
NAND3X1 NAND3X1_791 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n488_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n489_));
NAND3X1 NAND3X1_792 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n383_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n498_));
NAND3X1 NAND3X1_793 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n61_));
NAND3X1 NAND3X1_794 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n65_));
NAND3X1 NAND3X1_795 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n77_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n109_));
NAND3X1 NAND3X1_796 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n111_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n112_));
NAND3X1 NAND3X1_797 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n112_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n109_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n113_));
NAND3X1 NAND3X1_798 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n114_));
NAND3X1 NAND3X1_799 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n115_));
NAND3X1 NAND3X1_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n123_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n190_));
NAND3X1 NAND3X1_80 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2969_));
NAND3X1 NAND3X1_800 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n114_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n116_));
NAND3X1 NAND3X1_801 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n116_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n118_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n119_));
NAND3X1 NAND3X1_802 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n130_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n133_));
NAND3X1 NAND3X1_803 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n144_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n148_));
NAND3X1 NAND3X1_804 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n148_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n143_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n149_));
NAND3X1 NAND3X1_805 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n164_));
NAND3X1 NAND3X1_806 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n169_));
NAND3X1 NAND3X1_807 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_));
NAND3X1 NAND3X1_808 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n178_));
NAND3X1 NAND3X1_809 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n142_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n181_));
NAND3X1 NAND3X1_81 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2970_));
NAND3X1 NAND3X1_810 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n182_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n183_));
NAND3X1 NAND3X1_811 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_));
NAND3X1 NAND3X1_812 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n156_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n198_));
NAND3X1 NAND3X1_813 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n198_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n183_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n178_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n199_));
NAND3X1 NAND3X1_814 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n207_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n211_));
NAND3X1 NAND3X1_815 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n219_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n222_));
NAND3X1 NAND3X1_816 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n235_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n236_));
NAND3X1 NAND3X1_817 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n238_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n239_));
NAND3X1 NAND3X1_818 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n255_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n256_));
NAND3X1 NAND3X1_819 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n257_));
NAND3X1 NAND3X1_82 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2969_), .B(AES_CORE_DATAPATH__abc_15863_new_n2970_), .C(AES_CORE_DATAPATH__abc_15863_new_n2971_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2972_));
NAND3X1 NAND3X1_820 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n194_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n259_));
NAND3X1 NAND3X1_821 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n263_));
NAND3X1 NAND3X1_822 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n267_));
NAND3X1 NAND3X1_823 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n269_));
NAND3X1 NAND3X1_824 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n272_));
NAND3X1 NAND3X1_825 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n273_));
NAND3X1 NAND3X1_826 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n238_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n296_));
NAND3X1 NAND3X1_827 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n297_));
NAND3X1 NAND3X1_828 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n230_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n298_));
NAND3X1 NAND3X1_829 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n298_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n296_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n299_));
NAND3X1 NAND3X1_83 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2980_));
NAND3X1 NAND3X1_830 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n315_));
NAND3X1 NAND3X1_831 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n318_));
NAND3X1 NAND3X1_832 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n318_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n320_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n321_));
NAND3X1 NAND3X1_833 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n322_));
NAND3X1 NAND3X1_834 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n323_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n324_));
NAND3X1 NAND3X1_835 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n308_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n340_));
NAND3X1 NAND3X1_836 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n341_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n342_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n344_));
NAND3X1 NAND3X1_837 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n320_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n348_));
NAND3X1 NAND3X1_838 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n323_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n349_));
NAND3X1 NAND3X1_839 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n334_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n352_));
NAND3X1 NAND3X1_84 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2981_));
NAND3X1 NAND3X1_840 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n354_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n356_));
NAND3X1 NAND3X1_841 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n357_));
NAND3X1 NAND3X1_842 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n358_));
NAND3X1 NAND3X1_843 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n359_));
NAND3X1 NAND3X1_844 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n360_));
NAND3X1 NAND3X1_845 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n361_));
NAND3X1 NAND3X1_846 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n319_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n362_));
NAND3X1 NAND3X1_847 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n365_));
NAND3X1 NAND3X1_848 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n366_));
NAND3X1 NAND3X1_849 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n377_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n378_));
NAND3X1 NAND3X1_85 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2980_), .B(AES_CORE_DATAPATH__abc_15863_new_n2981_), .C(AES_CORE_DATAPATH__abc_15863_new_n2982_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2983_));
NAND3X1 NAND3X1_850 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n381_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n383_));
NAND3X1 NAND3X1_851 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n386_));
NAND3X1 NAND3X1_852 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n91_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n389_));
NAND3X1 NAND3X1_853 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n390_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n391_));
NAND3X1 NAND3X1_854 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n392_));
NAND3X1 NAND3X1_855 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n408_));
NAND3X1 NAND3X1_856 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n409_));
NAND3X1 NAND3X1_857 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n423_));
NAND3X1 NAND3X1_858 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n424_));
NAND3X1 NAND3X1_859 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n424_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n426_));
NAND3X1 NAND3X1_86 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2991_));
NAND3X1 NAND3X1_860 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n427_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n431_));
NAND3X1 NAND3X1_861 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n434_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n435_));
NAND3X1 NAND3X1_862 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n392_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n437_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n438_));
NAND3X1 NAND3X1_863 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n438_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n439_));
NAND3X1 NAND3X1_864 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n440_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n441_));
NAND3X1 NAND3X1_865 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n423_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n443_));
NAND3X1 NAND3X1_866 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n442_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n447_));
NAND3X1 NAND3X1_867 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n446_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n452_));
NAND3X1 NAND3X1_868 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n444_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n453_));
NAND3X1 NAND3X1_869 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n453_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n452_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n454_));
NAND3X1 NAND3X1_87 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2992_));
NAND3X1 NAND3X1_870 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n459_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n458_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n413_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n460_));
NAND3X1 NAND3X1_871 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n463_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n464_));
NAND3X1 NAND3X1_872 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n457_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n465_));
NAND3X1 NAND3X1_873 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n462_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n468_));
NAND3X1 NAND3X1_874 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n468_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n470_));
NAND3X1 NAND3X1_875 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n470_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n465_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n471_));
NAND3X1 NAND3X1_876 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n472_));
NAND3X1 NAND3X1_877 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n457_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n473_));
NAND3X1 NAND3X1_878 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n473_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n474_));
NAND3X1 NAND3X1_879 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n477_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n480_));
NAND3X1 NAND3X1_88 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2991_), .B(AES_CORE_DATAPATH__abc_15863_new_n2992_), .C(AES_CORE_DATAPATH__abc_15863_new_n2993_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2994_));
NAND3X1 NAND3X1_880 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n479_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n481_));
NAND3X1 NAND3X1_881 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n478_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n483_));
NAND3X1 NAND3X1_882 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n483_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n484_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n485_));
NAND3X1 NAND3X1_883 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n451_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n481_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n486_));
NAND3X1 NAND3X1_884 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n483_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n484_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n487_));
NAND3X1 NAND3X1_885 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n480_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n488_));
NAND3X1 NAND3X1_886 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n488_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n489_));
NAND3X1 NAND3X1_887 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n383_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n498_));
NAND3X1 NAND3X1_888 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n61_));
NAND3X1 NAND3X1_889 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n65_));
NAND3X1 NAND3X1_89 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3003_));
NAND3X1 NAND3X1_890 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n73_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n77_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n109_));
NAND3X1 NAND3X1_891 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n110_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n111_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n112_));
NAND3X1 NAND3X1_892 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n112_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n109_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n113_));
NAND3X1 NAND3X1_893 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n64_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n114_));
NAND3X1 NAND3X1_894 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n60_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n115_));
NAND3X1 NAND3X1_895 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n114_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n116_));
NAND3X1 NAND3X1_896 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n116_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n118_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n119_));
NAND3X1 NAND3X1_897 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n130_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n133_));
NAND3X1 NAND3X1_898 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n144_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n148_));
NAND3X1 NAND3X1_899 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n148_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n143_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n149_));
NAND3X1 NAND3X1_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n136_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_), .Y(AES_CORE_CONTROL_UNIT_key_en_2_));
NAND3X1 NAND3X1_90 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3004_));
NAND3X1 NAND3X1_900 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n146_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n164_));
NAND3X1 NAND3X1_901 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n169_));
NAND3X1 NAND3X1_902 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n176_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_));
NAND3X1 NAND3X1_903 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n178_));
NAND3X1 NAND3X1_904 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n142_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n181_));
NAND3X1 NAND3X1_905 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n182_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n183_));
NAND3X1 NAND3X1_906 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n163_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n164_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_));
NAND3X1 NAND3X1_907 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n156_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n198_));
NAND3X1 NAND3X1_908 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n198_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n183_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n178_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n199_));
NAND3X1 NAND3X1_909 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n207_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n211_));
NAND3X1 NAND3X1_91 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3003_), .B(AES_CORE_DATAPATH__abc_15863_new_n3004_), .C(AES_CORE_DATAPATH__abc_15863_new_n3005_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3006_));
NAND3X1 NAND3X1_910 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n219_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n222_));
NAND3X1 NAND3X1_911 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n235_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n236_));
NAND3X1 NAND3X1_912 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n238_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n239_));
NAND3X1 NAND3X1_913 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n149_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n255_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n256_));
NAND3X1 NAND3X1_914 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n257_));
NAND3X1 NAND3X1_915 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n194_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n150_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n259_));
NAND3X1 NAND3X1_916 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n263_));
NAND3X1 NAND3X1_917 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n267_));
NAND3X1 NAND3X1_918 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n269_));
NAND3X1 NAND3X1_919 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n258_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n272_));
NAND3X1 NAND3X1_92 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3013_));
NAND3X1 NAND3X1_920 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n262_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n264_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n273_));
NAND3X1 NAND3X1_921 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n238_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n180_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n296_));
NAND3X1 NAND3X1_922 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n173_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n297_));
NAND3X1 NAND3X1_923 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n230_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n185_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n298_));
NAND3X1 NAND3X1_924 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n298_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n296_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n299_));
NAND3X1 NAND3X1_925 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n247_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n315_));
NAND3X1 NAND3X1_926 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n318_));
NAND3X1 NAND3X1_927 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n318_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n320_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n321_));
NAND3X1 NAND3X1_928 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n313_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n322_));
NAND3X1 NAND3X1_929 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n323_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n324_));
NAND3X1 NAND3X1_93 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3014_));
NAND3X1 NAND3X1_930 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n308_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n340_));
NAND3X1 NAND3X1_931 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n341_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n342_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n344_));
NAND3X1 NAND3X1_932 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n320_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n348_));
NAND3X1 NAND3X1_933 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n323_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n322_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n349_));
NAND3X1 NAND3X1_934 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n334_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n352_));
NAND3X1 NAND3X1_935 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n354_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n356_));
NAND3X1 NAND3X1_936 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n357_));
NAND3X1 NAND3X1_937 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n358_));
NAND3X1 NAND3X1_938 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n359_));
NAND3X1 NAND3X1_939 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n317_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n352_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n356_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n360_));
NAND3X1 NAND3X1_94 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3013_), .B(AES_CORE_DATAPATH__abc_15863_new_n3014_), .C(AES_CORE_DATAPATH__abc_15863_new_n3015_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3016_));
NAND3X1 NAND3X1_940 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n340_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n361_));
NAND3X1 NAND3X1_941 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n319_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n362_));
NAND3X1 NAND3X1_942 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n357_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n365_));
NAND3X1 NAND3X1_943 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n360_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n361_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n366_));
NAND3X1 NAND3X1_944 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n377_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n370_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n378_));
NAND3X1 NAND3X1_945 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n381_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n382_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n383_));
NAND3X1 NAND3X1_946 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n386_));
NAND3X1 NAND3X1_947 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n91_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n389_));
NAND3X1 NAND3X1_948 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n390_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n391_));
NAND3X1 NAND3X1_949 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n392_));
NAND3X1 NAND3X1_95 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3023_));
NAND3X1 NAND3X1_950 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n408_));
NAND3X1 NAND3X1_951 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n409_));
NAND3X1 NAND3X1_952 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n388_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n391_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n423_));
NAND3X1 NAND3X1_953 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n113_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n424_));
NAND3X1 NAND3X1_954 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n424_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n426_));
NAND3X1 NAND3X1_955 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n430_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n427_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n429_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n431_));
NAND3X1 NAND3X1_956 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n434_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n435_));
NAND3X1 NAND3X1_957 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n392_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n437_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n438_));
NAND3X1 NAND3X1_958 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n438_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n439_));
NAND3X1 NAND3X1_959 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n440_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n441_));
NAND3X1 NAND3X1_96 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3024_));
NAND3X1 NAND3X1_960 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n423_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n443_));
NAND3X1 NAND3X1_961 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n427_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n442_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n447_));
NAND3X1 NAND3X1_962 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n446_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n452_));
NAND3X1 NAND3X1_963 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n441_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n444_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n453_));
NAND3X1 NAND3X1_964 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n453_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n452_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n454_));
NAND3X1 NAND3X1_965 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n459_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n458_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n413_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n460_));
NAND3X1 NAND3X1_966 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n463_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n464_));
NAND3X1 NAND3X1_967 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n457_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n465_));
NAND3X1 NAND3X1_968 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n462_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n468_));
NAND3X1 NAND3X1_969 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n468_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n470_));
NAND3X1 NAND3X1_97 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3023_), .B(AES_CORE_DATAPATH__abc_15863_new_n3024_), .C(AES_CORE_DATAPATH__abc_15863_new_n3025_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3026_));
NAND3X1 NAND3X1_970 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n470_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n465_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n471_));
NAND3X1 NAND3X1_971 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n464_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n472_));
NAND3X1 NAND3X1_972 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n457_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n469_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n473_));
NAND3X1 NAND3X1_973 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n473_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n474_));
NAND3X1 NAND3X1_974 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n477_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n480_));
NAND3X1 NAND3X1_975 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n479_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n481_));
NAND3X1 NAND3X1_976 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n437_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n478_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n466_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n483_));
NAND3X1 NAND3X1_977 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n483_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n484_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n485_));
NAND3X1 NAND3X1_978 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n451_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n481_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n486_));
NAND3X1 NAND3X1_979 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n483_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n484_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n487_));
NAND3X1 NAND3X1_98 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .C(AES_CORE_DATAPATH__abc_15863_new_n2735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3034_));
NAND3X1 NAND3X1_980 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n480_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n488_));
NAND3X1 NAND3X1_981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n488_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n489_));
NAND3X1 NAND3X1_982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n343_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n383_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n498_));
NAND3X1 NAND3X1_983 ( .A(\data_type[0] ), .B(\bus_in[16] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n68_));
NAND3X1 NAND3X1_984 ( .A(\data_type[1] ), .B(\bus_in[24] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n70_));
NAND3X1 NAND3X1_985 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n68_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n70_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n73_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_));
NAND3X1 NAND3X1_986 ( .A(\data_type[0] ), .B(\bus_in[17] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n75_));
NAND3X1 NAND3X1_987 ( .A(\data_type[1] ), .B(\bus_in[25] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n76_));
NAND3X1 NAND3X1_988 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n75_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n76_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n77_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_));
NAND3X1 NAND3X1_989 ( .A(\data_type[0] ), .B(\bus_in[18] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n79_));
NAND3X1 NAND3X1_99 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n2721_), .C(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3035_));
NAND3X1 NAND3X1_990 ( .A(\data_type[1] ), .B(\bus_in[26] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n80_));
NAND3X1 NAND3X1_991 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n79_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n80_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n81_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_));
NAND3X1 NAND3X1_992 ( .A(\data_type[0] ), .B(\bus_in[19] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n83_));
NAND3X1 NAND3X1_993 ( .A(\data_type[1] ), .B(\bus_in[27] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n84_));
NAND3X1 NAND3X1_994 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n83_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n84_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n85_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_));
NAND3X1 NAND3X1_995 ( .A(\data_type[0] ), .B(\bus_in[20] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n87_));
NAND3X1 NAND3X1_996 ( .A(\data_type[1] ), .B(\bus_in[28] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n88_));
NAND3X1 NAND3X1_997 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n87_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n88_), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n89_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_));
NAND3X1 NAND3X1_998 ( .A(\data_type[0] ), .B(\bus_in[21] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n67_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n91_));
NAND3X1 NAND3X1_999 ( .A(\data_type[1] ), .B(\bus_in[29] ), .C(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n69_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n92_));
NOR2X1 NOR2X1_1 ( .A(\addr[1] ), .B(_abc_15574_new_n13_), .Y(AES_CORE_DATAPATH_col_en_host_1_));
NOR2X1 NOR2X1_10 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_));
NOR2X1 NOR2X1_100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4363_));
NOR2X1 NOR2X1_101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4368_));
NOR2X1 NOR2X1_102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4374_));
NOR2X1 NOR2X1_103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4378_));
NOR2X1 NOR2X1_104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4380_));
NOR2X1 NOR2X1_105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4382_));
NOR2X1 NOR2X1_106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4384_));
NOR2X1 NOR2X1_107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4386_));
NOR2X1 NOR2X1_108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4388_));
NOR2X1 NOR2X1_109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4390_));
NOR2X1 NOR2X1_11 ( .A(disable_core), .B(end_aes), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n112_));
NOR2X1 NOR2X1_110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4392_));
NOR2X1 NOR2X1_111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4394_));
NOR2X1 NOR2X1_112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4396_));
NOR2X1 NOR2X1_113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4398_));
NOR2X1 NOR2X1_114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4400_));
NOR2X1 NOR2X1_115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4402_));
NOR2X1 NOR2X1_116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4404_));
NOR2X1 NOR2X1_117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4406_));
NOR2X1 NOR2X1_118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4408_));
NOR2X1 NOR2X1_119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4410_));
NOR2X1 NOR2X1_12 ( .A(AES_CORE_CONTROL_UNIT_rd_count_1_), .B(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n114_));
NOR2X1 NOR2X1_120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4412_));
NOR2X1 NOR2X1_121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4414_));
NOR2X1 NOR2X1_122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4416_));
NOR2X1 NOR2X1_123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4418_));
NOR2X1 NOR2X1_124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4420_));
NOR2X1 NOR2X1_125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4422_));
NOR2X1 NOR2X1_126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4424_));
NOR2X1 NOR2X1_127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4426_));
NOR2X1 NOR2X1_128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4428_));
NOR2X1 NOR2X1_129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4430_));
NOR2X1 NOR2X1_13 ( .A(AES_CORE_CONTROL_UNIT_rd_count_3_), .B(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n115_));
NOR2X1 NOR2X1_130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4432_));
NOR2X1 NOR2X1_131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4434_));
NOR2X1 NOR2X1_132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4436_));
NOR2X1 NOR2X1_133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4438_));
NOR2X1 NOR2X1_134 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4575_), .B(AES_CORE_DATAPATH__abc_15863_new_n4578_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4579_));
NOR2X1 NOR2X1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4581_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4582_));
NOR2X1 NOR2X1_136 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4575_), .B(AES_CORE_DATAPATH__abc_15863_new_n4584_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4585_));
NOR2X1 NOR2X1_137 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n2715_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4592_));
NOR2X1 NOR2X1_138 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4597_));
NOR2X1 NOR2X1_139 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4618_));
NOR2X1 NOR2X1_14 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n123_));
NOR2X1 NOR2X1_140 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_15863_new_n4623_));
NOR2X1 NOR2X1_141 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4626_));
NOR2X1 NOR2X1_142 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4634_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4635_));
NOR2X1 NOR2X1_143 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4638_));
NOR2X1 NOR2X1_144 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4673_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4674_));
NOR2X1 NOR2X1_145 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4712_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4713_));
NOR2X1 NOR2X1_146 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4719_));
NOR2X1 NOR2X1_147 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3180_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4746_));
NOR2X1 NOR2X1_148 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4752_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4753_));
NOR2X1 NOR2X1_149 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4788_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4789_));
NOR2X1 NOR2X1_15 ( .A(AES_CORE_CONTROL_UNIT_state_8_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_));
NOR2X1 NOR2X1_150 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4827_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4828_));
NOR2X1 NOR2X1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4862_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4863_));
NOR2X1 NOR2X1_152 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4866_));
NOR2X1 NOR2X1_153 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4901_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4902_));
NOR2X1 NOR2X1_154 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4936_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4937_));
NOR2X1 NOR2X1_155 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4943_));
NOR2X1 NOR2X1_156 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3312_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4969_));
NOR2X1 NOR2X1_157 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4975_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4976_));
NOR2X1 NOR2X1_158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5014_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5015_));
NOR2X1 NOR2X1_159 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5021_));
NOR2X1 NOR2X1_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n129_));
NOR2X1 NOR2X1_160 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3356_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5047_));
NOR2X1 NOR2X1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5053_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5054_));
NOR2X1 NOR2X1_162 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5092_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5093_));
NOR2X1 NOR2X1_163 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5099_));
NOR2X1 NOR2X1_164 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3400_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5125_));
NOR2X1 NOR2X1_165 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5131_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5132_));
NOR2X1 NOR2X1_166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5167_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5168_));
NOR2X1 NOR2X1_167 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5174_));
NOR2X1 NOR2X1_168 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3444_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5200_));
NOR2X1 NOR2X1_169 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5206_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5207_));
NOR2X1 NOR2X1_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n129_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n127_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n130_));
NOR2X1 NOR2X1_170 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5245_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5246_));
NOR2X1 NOR2X1_171 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5252_));
NOR2X1 NOR2X1_172 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3488_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5278_));
NOR2X1 NOR2X1_173 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5284_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5285_));
NOR2X1 NOR2X1_174 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5291_));
NOR2X1 NOR2X1_175 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3510_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5317_));
NOR2X1 NOR2X1_176 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5323_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5324_));
NOR2X1 NOR2X1_177 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5330_));
NOR2X1 NOR2X1_178 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3532_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5356_));
NOR2X1 NOR2X1_179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5362_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5363_));
NOR2X1 NOR2X1_18 ( .A(disable_core), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n130_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_10_));
NOR2X1 NOR2X1_180 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5401_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5402_));
NOR2X1 NOR2X1_181 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5408_));
NOR2X1 NOR2X1_182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3576_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5434_));
NOR2X1 NOR2X1_183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5440_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5441_));
NOR2X1 NOR2X1_184 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5476_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5477_));
NOR2X1 NOR2X1_185 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5480_));
NOR2X1 NOR2X1_186 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5515_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5516_));
NOR2X1 NOR2X1_187 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5554_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5555_));
NOR2X1 NOR2X1_188 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5561_));
NOR2X1 NOR2X1_189 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3664_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5587_));
NOR2X1 NOR2X1_19 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n146_));
NOR2X1 NOR2X1_190 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5593_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5594_));
NOR2X1 NOR2X1_191 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5600_));
NOR2X1 NOR2X1_192 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3686_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5626_));
NOR2X1 NOR2X1_193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5632_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5633_));
NOR2X1 NOR2X1_194 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5671_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5672_));
NOR2X1 NOR2X1_195 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5678_));
NOR2X1 NOR2X1_196 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3730_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5704_));
NOR2X1 NOR2X1_197 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5710_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5711_));
NOR2X1 NOR2X1_198 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5746_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5747_));
NOR2X1 NOR2X1_199 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5785_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5786_));
NOR2X1 NOR2X1_2 ( .A(\aes_mode[0] ), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_), .Y(AES_CORE_CONTROL_UNIT_mode_ctr));
NOR2X1 NOR2X1_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n151_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n154_));
NOR2X1 NOR2X1_200 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5792_));
NOR2X1 NOR2X1_201 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4745_), .B(AES_CORE_DATAPATH__abc_15863_new_n3796_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5818_));
NOR2X1 NOR2X1_202 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5989_));
NOR2X1 NOR2X1_203 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5991_));
NOR2X1 NOR2X1_204 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5993_));
NOR2X1 NOR2X1_205 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5995_));
NOR2X1 NOR2X1_206 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5997_));
NOR2X1 NOR2X1_207 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5999_));
NOR2X1 NOR2X1_208 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6001_));
NOR2X1 NOR2X1_209 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6003_));
NOR2X1 NOR2X1_21 ( .A(AES_CORE_CONTROL_UNIT_state_14_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n161_));
NOR2X1 NOR2X1_210 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6005_));
NOR2X1 NOR2X1_211 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6007_));
NOR2X1 NOR2X1_212 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6009_));
NOR2X1 NOR2X1_213 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6011_));
NOR2X1 NOR2X1_214 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6013_));
NOR2X1 NOR2X1_215 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6015_));
NOR2X1 NOR2X1_216 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6017_));
NOR2X1 NOR2X1_217 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6019_));
NOR2X1 NOR2X1_218 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6021_));
NOR2X1 NOR2X1_219 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6023_));
NOR2X1 NOR2X1_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n163_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n162_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_));
NOR2X1 NOR2X1_220 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6025_));
NOR2X1 NOR2X1_221 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6027_));
NOR2X1 NOR2X1_222 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6029_));
NOR2X1 NOR2X1_223 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6031_));
NOR2X1 NOR2X1_224 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6033_));
NOR2X1 NOR2X1_225 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6035_));
NOR2X1 NOR2X1_226 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6037_));
NOR2X1 NOR2X1_227 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6039_));
NOR2X1 NOR2X1_228 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6041_));
NOR2X1 NOR2X1_229 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6043_));
NOR2X1 NOR2X1_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_), .Y(AES_CORE_CONTROL_UNIT_rk_sel_0_));
NOR2X1 NOR2X1_230 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6045_));
NOR2X1 NOR2X1_231 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6047_));
NOR2X1 NOR2X1_232 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6049_));
NOR2X1 NOR2X1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6052_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6053_));
NOR2X1 NOR2X1_234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6059_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6060_));
NOR2X1 NOR2X1_235 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6066_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6067_));
NOR2X1 NOR2X1_236 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6073_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6074_));
NOR2X1 NOR2X1_237 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6080_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6081_));
NOR2X1 NOR2X1_238 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6087_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6088_));
NOR2X1 NOR2X1_239 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6094_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6095_));
NOR2X1 NOR2X1_24 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_), .Y(AES_CORE_CONTROL_UNIT_rk_sel_1_));
NOR2X1 NOR2X1_240 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6101_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6102_));
NOR2X1 NOR2X1_241 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6108_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6109_));
NOR2X1 NOR2X1_242 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6115_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6116_));
NOR2X1 NOR2X1_243 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6122_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6123_));
NOR2X1 NOR2X1_244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6129_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6130_));
NOR2X1 NOR2X1_245 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6136_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6137_));
NOR2X1 NOR2X1_246 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6143_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6144_));
NOR2X1 NOR2X1_247 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6150_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6151_));
NOR2X1 NOR2X1_248 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6157_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6158_));
NOR2X1 NOR2X1_249 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6164_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6165_));
NOR2X1 NOR2X1_25 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n167_));
NOR2X1 NOR2X1_250 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6171_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6172_));
NOR2X1 NOR2X1_251 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6178_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6179_));
NOR2X1 NOR2X1_252 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6185_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6186_));
NOR2X1 NOR2X1_253 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6192_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6193_));
NOR2X1 NOR2X1_254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6199_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6200_));
NOR2X1 NOR2X1_255 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6206_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6207_));
NOR2X1 NOR2X1_256 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6213_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6214_));
NOR2X1 NOR2X1_257 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6220_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6221_));
NOR2X1 NOR2X1_258 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6227_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6228_));
NOR2X1 NOR2X1_259 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6234_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6235_));
NOR2X1 NOR2X1_26 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n172_));
NOR2X1 NOR2X1_260 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6241_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6242_));
NOR2X1 NOR2X1_261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6248_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6249_));
NOR2X1 NOR2X1_262 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6255_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6256_));
NOR2X1 NOR2X1_263 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6262_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6263_));
NOR2X1 NOR2X1_264 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6269_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6270_));
NOR2X1 NOR2X1_265 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6276_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6277_));
NOR2X1 NOR2X1_266 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6283_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6284_));
NOR2X1 NOR2X1_267 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6290_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6291_));
NOR2X1 NOR2X1_268 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6297_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6298_));
NOR2X1 NOR2X1_269 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6304_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6305_));
NOR2X1 NOR2X1_27 ( .A(AES_CORE_CONTROL_UNIT_state_4_), .B(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_));
NOR2X1 NOR2X1_270 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6311_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6312_));
NOR2X1 NOR2X1_271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6318_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6319_));
NOR2X1 NOR2X1_272 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6325_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6326_));
NOR2X1 NOR2X1_273 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6332_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6333_));
NOR2X1 NOR2X1_274 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6339_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6340_));
NOR2X1 NOR2X1_275 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6346_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6347_));
NOR2X1 NOR2X1_276 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6353_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6354_));
NOR2X1 NOR2X1_277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6360_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6361_));
NOR2X1 NOR2X1_278 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6367_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6368_));
NOR2X1 NOR2X1_279 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6374_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6375_));
NOR2X1 NOR2X1_28 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n176_));
NOR2X1 NOR2X1_280 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6381_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6382_));
NOR2X1 NOR2X1_281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6388_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6389_));
NOR2X1 NOR2X1_282 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6395_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6396_));
NOR2X1 NOR2X1_283 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6402_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6403_));
NOR2X1 NOR2X1_284 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6409_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6410_));
NOR2X1 NOR2X1_285 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6416_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6417_));
NOR2X1 NOR2X1_286 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6423_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6424_));
NOR2X1 NOR2X1_287 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6430_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6431_));
NOR2X1 NOR2X1_288 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6437_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6438_));
NOR2X1 NOR2X1_289 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6444_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6445_));
NOR2X1 NOR2X1_29 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_));
NOR2X1 NOR2X1_290 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6451_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6452_));
NOR2X1 NOR2X1_291 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6458_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6459_));
NOR2X1 NOR2X1_292 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6465_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6466_));
NOR2X1 NOR2X1_293 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6472_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6473_));
NOR2X1 NOR2X1_294 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6479_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6480_));
NOR2X1 NOR2X1_295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6486_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6487_));
NOR2X1 NOR2X1_296 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6493_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6494_));
NOR2X1 NOR2X1_297 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6501_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6502_));
NOR2X1 NOR2X1_298 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6507_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6508_));
NOR2X1 NOR2X1_299 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6514_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6515_));
NOR2X1 NOR2X1_3 ( .A(AES_CORE_CONTROL_UNIT_state_7_), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n78_));
NOR2X1 NOR2X1_30 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n182_));
NOR2X1 NOR2X1_300 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6520_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6521_));
NOR2X1 NOR2X1_301 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6527_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6528_));
NOR2X1 NOR2X1_302 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6534_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6535_));
NOR2X1 NOR2X1_303 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6541_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6542_));
NOR2X1 NOR2X1_304 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6547_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6548_));
NOR2X1 NOR2X1_305 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6554_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6555_));
NOR2X1 NOR2X1_306 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6560_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6561_));
NOR2X1 NOR2X1_307 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6567_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6568_));
NOR2X1 NOR2X1_308 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6573_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6574_));
NOR2X1 NOR2X1_309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6580_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6581_));
NOR2X1 NOR2X1_31 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n133_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n195_));
NOR2X1 NOR2X1_310 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6586_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6587_));
NOR2X1 NOR2X1_311 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6593_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6594_));
NOR2X1 NOR2X1_312 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6599_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6600_));
NOR2X1 NOR2X1_313 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6606_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6607_));
NOR2X1 NOR2X1_314 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6612_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6613_));
NOR2X1 NOR2X1_315 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6618_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6619_));
NOR2X1 NOR2X1_316 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6624_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6625_));
NOR2X1 NOR2X1_317 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6631_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6632_));
NOR2X1 NOR2X1_318 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6637_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6638_));
NOR2X1 NOR2X1_319 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6644_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6645_));
NOR2X1 NOR2X1_32 ( .A(disable_core), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1856));
NOR2X1 NOR2X1_320 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6650_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6651_));
NOR2X1 NOR2X1_321 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6657_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6658_));
NOR2X1 NOR2X1_322 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6663_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6664_));
NOR2X1 NOR2X1_323 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6669_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6670_));
NOR2X1 NOR2X1_324 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6676_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6677_));
NOR2X1 NOR2X1_325 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6682_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6683_));
NOR2X1 NOR2X1_326 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6689_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6690_));
NOR2X1 NOR2X1_327 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6696_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6697_));
NOR2X1 NOR2X1_328 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6702_), .B(AES_CORE_DATAPATH__abc_15863_new_n4580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6703_));
NOR2X1 NOR2X1_329 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n6708_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6710_));
NOR2X1 NOR2X1_33 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n139_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n116_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_));
NOR2X1 NOR2X1_330 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4612_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6782_));
NOR2X1 NOR2X1_331 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6782_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6783_));
NOR2X1 NOR2X1_332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6788_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6789_));
NOR2X1 NOR2X1_333 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4694_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6794_));
NOR2X1 NOR2X1_334 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6794_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6795_));
NOR2X1 NOR2X1_335 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6800_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6801_));
NOR2X1 NOR2X1_336 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4770_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6807_));
NOR2X1 NOR2X1_337 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6807_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6808_));
NOR2X1 NOR2X1_338 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4809_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6813_));
NOR2X1 NOR2X1_339 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6813_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6814_));
NOR2X1 NOR2X1_34 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n210_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n91_), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en));
NOR2X1 NOR2X1_340 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4845_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6820_));
NOR2X1 NOR2X1_341 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6820_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6821_));
NOR2X1 NOR2X1_342 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6826_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6827_));
NOR2X1 NOR2X1_343 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4919_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6833_));
NOR2X1 NOR2X1_344 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6833_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6834_));
NOR2X1 NOR2X1_345 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6839_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6840_));
NOR2X1 NOR2X1_346 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n4996_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6845_));
NOR2X1 NOR2X1_347 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6845_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6846_));
NOR2X1 NOR2X1_348 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6851_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6852_));
NOR2X1 NOR2X1_349 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5074_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6857_));
NOR2X1 NOR2X1_35 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n212_), .Y(AES_CORE_CONTROL_UNIT_iv_cnt_en));
NOR2X1 NOR2X1_350 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6857_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6858_));
NOR2X1 NOR2X1_351 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6863_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6864_));
NOR2X1 NOR2X1_352 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5149_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6870_));
NOR2X1 NOR2X1_353 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6870_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6871_));
NOR2X1 NOR2X1_354 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6876_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6877_));
NOR2X1 NOR2X1_355 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5227_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6882_));
NOR2X1 NOR2X1_356 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6882_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6883_));
NOR2X1 NOR2X1_357 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6888_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6889_));
NOR2X1 NOR2X1_358 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6894_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6895_));
NOR2X1 NOR2X1_359 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6900_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6901_));
NOR2X1 NOR2X1_36 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2463_));
NOR2X1 NOR2X1_360 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5383_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6906_));
NOR2X1 NOR2X1_361 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6906_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6907_));
NOR2X1 NOR2X1_362 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6912_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6913_));
NOR2X1 NOR2X1_363 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5458_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6919_));
NOR2X1 NOR2X1_364 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6919_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6920_));
NOR2X1 NOR2X1_365 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6925_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6926_));
NOR2X1 NOR2X1_366 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5536_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6931_));
NOR2X1 NOR2X1_367 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6931_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6932_));
NOR2X1 NOR2X1_368 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6937_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6938_));
NOR2X1 NOR2X1_369 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6943_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6944_));
NOR2X1 NOR2X1_37 ( .A(\iv_sel_rd[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2467_));
NOR2X1 NOR2X1_370 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5653_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6949_));
NOR2X1 NOR2X1_371 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6949_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6950_));
NOR2X1 NOR2X1_372 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6955_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6956_));
NOR2X1 NOR2X1_373 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6962_));
NOR2X1 NOR2X1_374 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6962_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6963_));
NOR2X1 NOR2X1_375 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n5767_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6968_));
NOR2X1 NOR2X1_376 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6968_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6969_));
NOR2X1 NOR2X1_377 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6974_), .B(AES_CORE_DATAPATH__abc_15863_new_n6713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6975_));
NOR2X1 NOR2X1_378 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(\iv_en[3] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n6977_));
NOR2X1 NOR2X1_379 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6981_));
NOR2X1 NOR2X1_38 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2721_), .B(AES_CORE_DATAPATH__abc_15863_new_n2728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2729_));
NOR2X1 NOR2X1_380 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2494_), .B(AES_CORE_DATAPATH__abc_15863_new_n6988_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6995_));
NOR2X1 NOR2X1_381 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6986_), .B(AES_CORE_DATAPATH__abc_15863_new_n7000_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7001_));
NOR2X1 NOR2X1_382 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2716_), .B(AES_CORE_DATAPATH__abc_15863_new_n7002_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7003_));
NOR2X1 NOR2X1_383 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2508_), .B(AES_CORE_DATAPATH__abc_15863_new_n7008_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7009_));
NOR2X1 NOR2X1_384 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2508_), .B(AES_CORE_DATAPATH__abc_15863_new_n2514_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7014_));
NOR2X1 NOR2X1_385 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2520_), .B(AES_CORE_DATAPATH__abc_15863_new_n7026_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7027_));
NOR2X1 NOR2X1_386 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6982_), .B(AES_CORE_DATAPATH__abc_15863_new_n7029_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7030_));
NOR2X1 NOR2X1_387 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2536_), .B(AES_CORE_DATAPATH__abc_15863_new_n7028_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7034_));
NOR2X1 NOR2X1_388 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6982_), .B(AES_CORE_DATAPATH__abc_15863_new_n7034_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7035_));
NOR2X1 NOR2X1_389 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7039_));
NOR2X1 NOR2X1_39 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .B(\key_out[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2753_));
NOR2X1 NOR2X1_390 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7041_), .B(AES_CORE_DATAPATH__abc_15863_new_n7028_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7042_));
NOR2X1 NOR2X1_391 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2560_), .B(AES_CORE_DATAPATH__abc_15863_new_n7048_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7055_));
NOR2X1 NOR2X1_392 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2574_), .B(AES_CORE_DATAPATH__abc_15863_new_n7060_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7071_));
NOR2X1 NOR2X1_393 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7041_), .B(AES_CORE_DATAPATH__abc_15863_new_n7107_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7108_));
NOR2X1 NOR2X1_394 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2568_), .B(AES_CORE_DATAPATH__abc_15863_new_n2574_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7109_));
NOR2X1 NOR2X1_395 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2582_), .B(AES_CORE_DATAPATH__abc_15863_new_n2588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7110_));
NOR2X1 NOR2X1_396 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7111_), .B(AES_CORE_DATAPATH__abc_15863_new_n7028_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7112_));
NOR2X1 NOR2X1_397 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2596_), .B(AES_CORE_DATAPATH__abc_15863_new_n2602_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7113_));
NOR2X1 NOR2X1_398 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2610_), .B(AES_CORE_DATAPATH__abc_15863_new_n2618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7114_));
NOR2X1 NOR2X1_399 ( .A(AES_CORE_DATAPATH_iv_3__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n7117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7118_));
NOR2X1 NOR2X1_4 ( .A(AES_CORE_CONTROL_UNIT_state_13_), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n79_));
NOR2X1 NOR2X1_40 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .B(\key_out[7] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2817_));
NOR2X1 NOR2X1_400 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2626_), .B(AES_CORE_DATAPATH__abc_15863_new_n7117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7123_));
NOR2X1 NOR2X1_401 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2632_), .B(AES_CORE_DATAPATH__abc_15863_new_n7123_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7124_));
NOR2X1 NOR2X1_402 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7130_), .B(AES_CORE_DATAPATH__abc_15863_new_n7117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7131_));
NOR2X1 NOR2X1_403 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2640_), .B(AES_CORE_DATAPATH__abc_15863_new_n7131_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7132_));
NOR2X1 NOR2X1_404 ( .A(AES_CORE_DATAPATH_iv_3__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n7139_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7140_));
NOR2X1 NOR2X1_405 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7130_), .B(AES_CORE_DATAPATH__abc_15863_new_n7145_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7146_));
NOR2X1 NOR2X1_406 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2654_), .B(AES_CORE_DATAPATH__abc_15863_new_n7149_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7150_));
NOR2X1 NOR2X1_407 ( .A(AES_CORE_DATAPATH_iv_3__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n7148_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7151_));
NOR2X1 NOR2X1_408 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2654_), .B(AES_CORE_DATAPATH__abc_15863_new_n7148_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7156_));
NOR2X1 NOR2X1_409 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2660_), .B(AES_CORE_DATAPATH__abc_15863_new_n7156_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7157_));
NOR2X1 NOR2X1_41 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .B(\key_out[8] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2830_));
NOR2X1 NOR2X1_410 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2654_), .B(AES_CORE_DATAPATH__abc_15863_new_n2660_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7163_));
NOR2X1 NOR2X1_411 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2668_), .B(AES_CORE_DATAPATH__abc_15863_new_n7165_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7166_));
NOR2X1 NOR2X1_412 ( .A(AES_CORE_DATAPATH_iv_3__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n7164_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7167_));
NOR2X1 NOR2X1_413 ( .A(AES_CORE_DATAPATH_iv_3__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n7173_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7174_));
NOR2X1 NOR2X1_414 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7179_), .B(AES_CORE_DATAPATH__abc_15863_new_n7148_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7180_));
NOR2X1 NOR2X1_415 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2682_), .B(AES_CORE_DATAPATH__abc_15863_new_n7180_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7181_));
NOR2X1 NOR2X1_416 ( .A(AES_CORE_DATAPATH_iv_3__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n7182_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7183_));
NOR2X1 NOR2X1_417 ( .A(AES_CORE_DATAPATH_iv_3__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n7189_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7190_));
NOR2X1 NOR2X1_418 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7195_), .B(AES_CORE_DATAPATH__abc_15863_new_n7182_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7196_));
NOR2X1 NOR2X1_419 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2696_), .B(AES_CORE_DATAPATH__abc_15863_new_n7196_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7197_));
NOR2X1 NOR2X1_42 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_), .B(\key_out[20] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2953_));
NOR2X1 NOR2X1_420 ( .A(AES_CORE_DATAPATH_iv_3__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n7204_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7205_));
NOR2X1 NOR2X1_421 ( .A(AES_CORE_DATAPATH_iv_2__2_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7214_));
NOR2X1 NOR2X1_422 ( .A(AES_CORE_DATAPATH_iv_2__4_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7218_));
NOR2X1 NOR2X1_423 ( .A(AES_CORE_DATAPATH_iv_2__5_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7220_));
NOR2X1 NOR2X1_424 ( .A(AES_CORE_DATAPATH_iv_2__12_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7234_));
NOR2X1 NOR2X1_425 ( .A(AES_CORE_DATAPATH_iv_2__14_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7238_));
NOR2X1 NOR2X1_426 ( .A(AES_CORE_DATAPATH_iv_2__16_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7242_));
NOR2X1 NOR2X1_427 ( .A(AES_CORE_DATAPATH_iv_2__20_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7250_));
NOR2X1 NOR2X1_428 ( .A(AES_CORE_DATAPATH_iv_2__22_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7254_));
NOR2X1 NOR2X1_429 ( .A(AES_CORE_DATAPATH_iv_2__24_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7258_));
NOR2X1 NOR2X1_43 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .B(\key_out[23] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2986_));
NOR2X1 NOR2X1_430 ( .A(AES_CORE_DATAPATH_iv_2__27_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7264_));
NOR2X1 NOR2X1_431 ( .A(AES_CORE_DATAPATH_iv_2__29_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7268_));
NOR2X1 NOR2X1_432 ( .A(AES_CORE_DATAPATH_iv_2__30_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7270_));
NOR2X1 NOR2X1_433 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6782_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7342_));
NOR2X1 NOR2X1_434 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6788_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7347_));
NOR2X1 NOR2X1_435 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6794_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7352_));
NOR2X1 NOR2X1_436 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6800_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7357_));
NOR2X1 NOR2X1_437 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6807_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7362_));
NOR2X1 NOR2X1_438 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6813_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7367_));
NOR2X1 NOR2X1_439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6820_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7372_));
NOR2X1 NOR2X1_44 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .B(\key_out[24] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n2999_));
NOR2X1 NOR2X1_440 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6826_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7377_));
NOR2X1 NOR2X1_441 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6833_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7382_));
NOR2X1 NOR2X1_442 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6839_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7387_));
NOR2X1 NOR2X1_443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6845_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7392_));
NOR2X1 NOR2X1_444 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6851_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7397_));
NOR2X1 NOR2X1_445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6857_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7402_));
NOR2X1 NOR2X1_446 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6863_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7407_));
NOR2X1 NOR2X1_447 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6870_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7412_));
NOR2X1 NOR2X1_448 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6876_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7417_));
NOR2X1 NOR2X1_449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6882_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7422_));
NOR2X1 NOR2X1_45 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3076_), .B(AES_CORE_DATAPATH__abc_15863_new_n3079_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3080_));
NOR2X1 NOR2X1_450 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6888_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7427_));
NOR2X1 NOR2X1_451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6894_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7432_));
NOR2X1 NOR2X1_452 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6900_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7437_));
NOR2X1 NOR2X1_453 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6906_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7442_));
NOR2X1 NOR2X1_454 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6912_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7447_));
NOR2X1 NOR2X1_455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6919_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7452_));
NOR2X1 NOR2X1_456 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6925_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7457_));
NOR2X1 NOR2X1_457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6931_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7462_));
NOR2X1 NOR2X1_458 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6937_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7467_));
NOR2X1 NOR2X1_459 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6943_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7472_));
NOR2X1 NOR2X1_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3082_), .B(AES_CORE_DATAPATH__abc_15863_new_n3084_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3085_));
NOR2X1 NOR2X1_460 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6949_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7477_));
NOR2X1 NOR2X1_461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6955_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7482_));
NOR2X1 NOR2X1_462 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6962_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7487_));
NOR2X1 NOR2X1_463 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6968_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7492_));
NOR2X1 NOR2X1_464 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6974_), .B(AES_CORE_DATAPATH__abc_15863_new_n7274_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7497_));
NOR2X1 NOR2X1_465 ( .A(AES_CORE_DATAPATH_iv_1__1_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7501_));
NOR2X1 NOR2X1_466 ( .A(AES_CORE_DATAPATH_iv_1__2_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7503_));
NOR2X1 NOR2X1_467 ( .A(AES_CORE_DATAPATH_iv_1__3_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7505_));
NOR2X1 NOR2X1_468 ( .A(AES_CORE_DATAPATH_iv_1__4_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7507_));
NOR2X1 NOR2X1_469 ( .A(AES_CORE_DATAPATH_iv_1__5_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7509_));
NOR2X1 NOR2X1_47 ( .A(AES_CORE_DATAPATH_col_sel_host_0_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3087_));
NOR2X1 NOR2X1_470 ( .A(AES_CORE_DATAPATH_iv_1__12_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7523_));
NOR2X1 NOR2X1_471 ( .A(AES_CORE_DATAPATH_iv_1__13_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7525_));
NOR2X1 NOR2X1_472 ( .A(AES_CORE_DATAPATH_iv_1__14_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7527_));
NOR2X1 NOR2X1_473 ( .A(AES_CORE_DATAPATH_iv_1__15_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7529_));
NOR2X1 NOR2X1_474 ( .A(AES_CORE_DATAPATH_iv_1__16_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7531_));
NOR2X1 NOR2X1_475 ( .A(AES_CORE_DATAPATH_iv_1__17_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7533_));
NOR2X1 NOR2X1_476 ( .A(AES_CORE_DATAPATH_iv_1__18_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7535_));
NOR2X1 NOR2X1_477 ( .A(AES_CORE_DATAPATH_iv_1__19_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7537_));
NOR2X1 NOR2X1_478 ( .A(AES_CORE_DATAPATH_iv_1__20_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7539_));
NOR2X1 NOR2X1_479 ( .A(AES_CORE_DATAPATH_iv_1__21_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7541_));
NOR2X1 NOR2X1_48 ( .A(AES_CORE_DATAPATH_col_sel_host_1_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3088_));
NOR2X1 NOR2X1_480 ( .A(AES_CORE_DATAPATH_iv_1__22_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7543_));
NOR2X1 NOR2X1_481 ( .A(AES_CORE_DATAPATH_iv_1__23_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7545_));
NOR2X1 NOR2X1_482 ( .A(AES_CORE_DATAPATH_iv_1__24_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7547_));
NOR2X1 NOR2X1_483 ( .A(AES_CORE_DATAPATH_iv_1__25_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7549_));
NOR2X1 NOR2X1_484 ( .A(AES_CORE_DATAPATH_iv_1__26_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7551_));
NOR2X1 NOR2X1_485 ( .A(AES_CORE_DATAPATH_iv_1__27_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7553_));
NOR2X1 NOR2X1_486 ( .A(AES_CORE_DATAPATH_iv_1__28_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7555_));
NOR2X1 NOR2X1_487 ( .A(AES_CORE_DATAPATH_iv_1__29_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7557_));
NOR2X1 NOR2X1_488 ( .A(AES_CORE_DATAPATH_iv_1__30_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7559_));
NOR2X1 NOR2X1_489 ( .A(AES_CORE_DATAPATH_iv_1__31_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7561_));
NOR2X1 NOR2X1_49 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n3088_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3094_));
NOR2X1 NOR2X1_490 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6510_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7567_));
NOR2X1 NOR2X1_491 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6523_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7572_));
NOR2X1 NOR2X1_492 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6550_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7581_));
NOR2X1 NOR2X1_493 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7586_));
NOR2X1 NOR2X1_494 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6576_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7591_));
NOR2X1 NOR2X1_495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6589_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7596_));
NOR2X1 NOR2X1_496 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6602_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7601_));
NOR2X1 NOR2X1_497 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6615_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7606_));
NOR2X1 NOR2X1_498 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6621_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7609_));
NOR2X1 NOR2X1_499 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6627_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7612_));
NOR2X1 NOR2X1_5 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n83_), .Y(AES_CORE_CONTROL_UNIT_last_round));
NOR2X1 NOR2X1_50 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3076_), .B(AES_CORE_DATAPATH__abc_15863_new_n3098_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3100_));
NOR2X1 NOR2X1_500 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6640_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7617_));
NOR2X1 NOR2X1_501 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6653_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7622_));
NOR2X1 NOR2X1_502 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6666_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7627_));
NOR2X1 NOR2X1_503 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6672_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7630_));
NOR2X1 NOR2X1_504 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6685_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7635_));
NOR2X1 NOR2X1_505 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6705_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7642_));
NOR2X1 NOR2X1_506 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6782_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7648_));
NOR2X1 NOR2X1_507 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6788_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7653_));
NOR2X1 NOR2X1_508 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6794_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7659_));
NOR2X1 NOR2X1_509 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6800_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7664_));
NOR2X1 NOR2X1_51 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_rk_out_sel_pp2), .Y(AES_CORE_DATAPATH__abc_15863_new_n3108_));
NOR2X1 NOR2X1_510 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6807_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7670_));
NOR2X1 NOR2X1_511 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6813_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7676_));
NOR2X1 NOR2X1_512 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6820_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7682_));
NOR2X1 NOR2X1_513 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6826_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7687_));
NOR2X1 NOR2X1_514 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6833_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7693_));
NOR2X1 NOR2X1_515 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6839_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7698_));
NOR2X1 NOR2X1_516 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6845_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7704_));
NOR2X1 NOR2X1_517 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6851_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7709_));
NOR2X1 NOR2X1_518 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6857_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7715_));
NOR2X1 NOR2X1_519 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6863_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7720_));
NOR2X1 NOR2X1_52 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3110_), .B(AES_CORE_DATAPATH__abc_15863_new_n3106_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3111_));
NOR2X1 NOR2X1_520 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6870_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7726_));
NOR2X1 NOR2X1_521 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6876_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7731_));
NOR2X1 NOR2X1_522 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6882_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7737_));
NOR2X1 NOR2X1_523 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6888_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7742_));
NOR2X1 NOR2X1_524 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6894_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7747_));
NOR2X1 NOR2X1_525 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6900_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7752_));
NOR2X1 NOR2X1_526 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6906_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7758_));
NOR2X1 NOR2X1_527 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6912_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7763_));
NOR2X1 NOR2X1_528 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6919_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7769_));
NOR2X1 NOR2X1_529 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6925_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7774_));
NOR2X1 NOR2X1_53 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3133_), .B(AES_CORE_DATAPATH__abc_15863_new_n3130_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3134_));
NOR2X1 NOR2X1_530 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6931_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7780_));
NOR2X1 NOR2X1_531 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6937_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7785_));
NOR2X1 NOR2X1_532 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6943_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7790_));
NOR2X1 NOR2X1_533 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6949_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7796_));
NOR2X1 NOR2X1_534 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6955_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7801_));
NOR2X1 NOR2X1_535 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6962_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7807_));
NOR2X1 NOR2X1_536 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6968_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7813_));
NOR2X1 NOR2X1_537 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6974_), .B(AES_CORE_DATAPATH__abc_15863_new_n7563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7818_));
NOR2X1 NOR2X1_538 ( .A(AES_CORE_DATAPATH_iv_0__0_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7820_));
NOR2X1 NOR2X1_539 ( .A(AES_CORE_DATAPATH_iv_0__1_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7822_));
NOR2X1 NOR2X1_54 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3155_), .B(AES_CORE_DATAPATH__abc_15863_new_n3152_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3156_));
NOR2X1 NOR2X1_540 ( .A(AES_CORE_DATAPATH_iv_0__2_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7824_));
NOR2X1 NOR2X1_541 ( .A(AES_CORE_DATAPATH_iv_0__3_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7826_));
NOR2X1 NOR2X1_542 ( .A(AES_CORE_DATAPATH_iv_0__4_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7828_));
NOR2X1 NOR2X1_543 ( .A(AES_CORE_DATAPATH_iv_0__5_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7830_));
NOR2X1 NOR2X1_544 ( .A(AES_CORE_DATAPATH_iv_0__12_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7850_));
NOR2X1 NOR2X1_545 ( .A(AES_CORE_DATAPATH_iv_0__13_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7852_));
NOR2X1 NOR2X1_546 ( .A(AES_CORE_DATAPATH_iv_0__14_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7854_));
NOR2X1 NOR2X1_547 ( .A(AES_CORE_DATAPATH_iv_0__15_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7856_));
NOR2X1 NOR2X1_548 ( .A(AES_CORE_DATAPATH_iv_0__16_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7858_));
NOR2X1 NOR2X1_549 ( .A(AES_CORE_DATAPATH_iv_0__17_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7860_));
NOR2X1 NOR2X1_55 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3200_), .B(AES_CORE_DATAPATH__abc_15863_new_n3197_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3201_));
NOR2X1 NOR2X1_550 ( .A(AES_CORE_DATAPATH_iv_0__18_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7862_));
NOR2X1 NOR2X1_551 ( .A(AES_CORE_DATAPATH_iv_0__19_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7864_));
NOR2X1 NOR2X1_552 ( .A(AES_CORE_DATAPATH_iv_0__20_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7866_));
NOR2X1 NOR2X1_553 ( .A(AES_CORE_DATAPATH_iv_0__21_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7868_));
NOR2X1 NOR2X1_554 ( .A(AES_CORE_DATAPATH_iv_0__22_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7870_));
NOR2X1 NOR2X1_555 ( .A(AES_CORE_DATAPATH_iv_0__23_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7872_));
NOR2X1 NOR2X1_556 ( .A(AES_CORE_DATAPATH_iv_0__24_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7874_));
NOR2X1 NOR2X1_557 ( .A(AES_CORE_DATAPATH_iv_0__25_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7876_));
NOR2X1 NOR2X1_558 ( .A(AES_CORE_DATAPATH_iv_0__26_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7878_));
NOR2X1 NOR2X1_559 ( .A(AES_CORE_DATAPATH_iv_0__27_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7880_));
NOR2X1 NOR2X1_56 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3222_), .B(AES_CORE_DATAPATH__abc_15863_new_n3219_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3223_));
NOR2X1 NOR2X1_560 ( .A(AES_CORE_DATAPATH_iv_0__28_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7882_));
NOR2X1 NOR2X1_561 ( .A(AES_CORE_DATAPATH_iv_0__29_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7884_));
NOR2X1 NOR2X1_562 ( .A(AES_CORE_DATAPATH_iv_0__30_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7886_));
NOR2X1 NOR2X1_563 ( .A(AES_CORE_DATAPATH_iv_0__31_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_15863_new_n7888_));
NOR2X1 NOR2X1_564 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6782_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7959_));
NOR2X1 NOR2X1_565 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6788_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7965_));
NOR2X1 NOR2X1_566 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6794_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7971_));
NOR2X1 NOR2X1_567 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6800_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7977_));
NOR2X1 NOR2X1_568 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6807_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7983_));
NOR2X1 NOR2X1_569 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6813_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7989_));
NOR2X1 NOR2X1_57 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3244_), .B(AES_CORE_DATAPATH__abc_15863_new_n3241_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3245_));
NOR2X1 NOR2X1_570 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6820_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7995_));
NOR2X1 NOR2X1_571 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6826_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8001_));
NOR2X1 NOR2X1_572 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6833_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8007_));
NOR2X1 NOR2X1_573 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6839_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8013_));
NOR2X1 NOR2X1_574 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6845_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8019_));
NOR2X1 NOR2X1_575 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6851_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8025_));
NOR2X1 NOR2X1_576 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6857_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8031_));
NOR2X1 NOR2X1_577 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6863_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8037_));
NOR2X1 NOR2X1_578 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6870_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8043_));
NOR2X1 NOR2X1_579 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6876_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8049_));
NOR2X1 NOR2X1_58 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3266_), .B(AES_CORE_DATAPATH__abc_15863_new_n3263_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3267_));
NOR2X1 NOR2X1_580 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6882_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8055_));
NOR2X1 NOR2X1_581 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6888_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8061_));
NOR2X1 NOR2X1_582 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6894_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8067_));
NOR2X1 NOR2X1_583 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6900_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8073_));
NOR2X1 NOR2X1_584 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6906_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8079_));
NOR2X1 NOR2X1_585 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6912_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8085_));
NOR2X1 NOR2X1_586 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6919_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8091_));
NOR2X1 NOR2X1_587 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6925_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8097_));
NOR2X1 NOR2X1_588 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6931_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8103_));
NOR2X1 NOR2X1_589 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6937_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8109_));
NOR2X1 NOR2X1_59 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3288_), .B(AES_CORE_DATAPATH__abc_15863_new_n3285_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3289_));
NOR2X1 NOR2X1_590 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6943_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8115_));
NOR2X1 NOR2X1_591 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6949_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8121_));
NOR2X1 NOR2X1_592 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6955_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8127_));
NOR2X1 NOR2X1_593 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6962_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8133_));
NOR2X1 NOR2X1_594 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6968_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8139_));
NOR2X1 NOR2X1_595 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6974_), .B(AES_CORE_DATAPATH__abc_15863_new_n7890_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8145_));
NOR2X1 NOR2X1_596 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n2712_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out));
NOR2X1 NOR2X1_597 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n412_));
NOR2X1 NOR2X1_598 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n414_));
NOR2X1 NOR2X1_599 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n416_));
NOR2X1 NOR2X1_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n89_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n91_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n92_));
NOR2X1 NOR2X1_60 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3332_), .B(AES_CORE_DATAPATH__abc_15863_new_n3329_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3333_));
NOR2X1 NOR2X1_600 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n436_));
NOR2X1 NOR2X1_601 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n444_));
NOR2X1 NOR2X1_602 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n465_));
NOR2X1 NOR2X1_603 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n476_));
NOR2X1 NOR2X1_604 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n423_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n483_));
NOR2X1 NOR2X1_605 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n107_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n109_));
NOR2X1 NOR2X1_606 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n114_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n115_));
NOR2X1 NOR2X1_607 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n116_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n117_));
NOR2X1 NOR2X1_608 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n132_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n137_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n138_));
NOR2X1 NOR2X1_609 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n139_));
NOR2X1 NOR2X1_61 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3376_), .B(AES_CORE_DATAPATH__abc_15863_new_n3373_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3377_));
NOR2X1 NOR2X1_610 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n139_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n140_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n141_));
NOR2X1 NOR2X1_611 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n149_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n148_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n150_));
NOR2X1 NOR2X1_612 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n145_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n151_));
NOR2X1 NOR2X1_613 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n142_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n152_));
NOR2X1 NOR2X1_614 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n163_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n164_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n165_));
NOR2X1 NOR2X1_615 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n167_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n166_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n168_));
NOR2X1 NOR2X1_616 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n165_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n168_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n169_));
NOR2X1 NOR2X1_617 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n174_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n176_));
NOR2X1 NOR2X1_618 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n141_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n182_));
NOR2X1 NOR2X1_619 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n141_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n184_));
NOR2X1 NOR2X1_62 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3420_), .B(AES_CORE_DATAPATH__abc_15863_new_n3417_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3421_));
NOR2X1 NOR2X1_620 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n174_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n185_));
NOR2X1 NOR2X1_621 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n163_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n167_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n188_));
NOR2X1 NOR2X1_622 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n164_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n166_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n189_));
NOR2X1 NOR2X1_623 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n188_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n189_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n190_));
NOR2X1 NOR2X1_624 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n97_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n202_));
NOR2X1 NOR2X1_625 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n203_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n204_));
NOR2X1 NOR2X1_626 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n97_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n206_));
NOR2X1 NOR2X1_627 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n203_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n207_));
NOR2X1 NOR2X1_628 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n213_));
NOR2X1 NOR2X1_629 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n217_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n218_));
NOR2X1 NOR2X1_63 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3464_), .B(AES_CORE_DATAPATH__abc_15863_new_n3461_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3465_));
NOR2X1 NOR2X1_630 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n219_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n220_));
NOR2X1 NOR2X1_631 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n247_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n248_));
NOR2X1 NOR2X1_632 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n249_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n250_));
NOR2X1 NOR2X1_633 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n251_));
NOR2X1 NOR2X1_634 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n171_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n252_));
NOR2X1 NOR2X1_635 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n254_));
NOR2X1 NOR2X1_636 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n264_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n265_));
NOR2X1 NOR2X1_637 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n271_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n273_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n274_));
NOR2X1 NOR2X1_638 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n207_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n206_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n374_));
NOR2X1 NOR2X1_639 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n202_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n204_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n376_));
NOR2X1 NOR2X1_64 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3552_), .B(AES_CORE_DATAPATH__abc_15863_new_n3549_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3553_));
NOR2X1 NOR2X1_640 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n305_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n308_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n400_));
NOR2X1 NOR2X1_641 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n426_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n429_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_));
NOR2X1 NOR2X1_642 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n525_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n524_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_));
NOR2X1 NOR2X1_643 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n56_));
NOR2X1 NOR2X1_644 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n67_));
NOR2X1 NOR2X1_645 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n81_));
NOR2X1 NOR2X1_646 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n82_));
NOR2X1 NOR2X1_647 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_));
NOR2X1 NOR2X1_648 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n106_));
NOR2X1 NOR2X1_649 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n137_));
NOR2X1 NOR2X1_65 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3596_), .B(AES_CORE_DATAPATH__abc_15863_new_n3593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3597_));
NOR2X1 NOR2X1_650 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n140_));
NOR2X1 NOR2X1_651 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n286_));
NOR2X1 NOR2X1_652 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n287_));
NOR2X1 NOR2X1_653 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n327_));
NOR2X1 NOR2X1_654 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n328_));
NOR2X1 NOR2X1_655 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n339_));
NOR2X1 NOR2X1_656 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n336_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n343_));
NOR2X1 NOR2X1_657 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n351_));
NOR2X1 NOR2X1_658 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n312_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n353_));
NOR2X1 NOR2X1_659 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n371_));
NOR2X1 NOR2X1_66 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3618_), .B(AES_CORE_DATAPATH__abc_15863_new_n3615_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3619_));
NOR2X1 NOR2X1_660 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n200_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n372_));
NOR2X1 NOR2X1_661 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n379_));
NOR2X1 NOR2X1_662 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n380_));
NOR2X1 NOR2X1_663 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n394_));
NOR2X1 NOR2X1_664 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n400_));
NOR2X1 NOR2X1_665 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n414_));
NOR2X1 NOR2X1_666 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n416_));
NOR2X1 NOR2X1_667 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n420_));
NOR2X1 NOR2X1_668 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n432_));
NOR2X1 NOR2X1_669 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n457_));
NOR2X1 NOR2X1_67 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3640_), .B(AES_CORE_DATAPATH__abc_15863_new_n3637_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3641_));
NOR2X1 NOR2X1_670 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n482_));
NOR2X1 NOR2X1_671 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n500_));
NOR2X1 NOR2X1_672 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n56_));
NOR2X1 NOR2X1_673 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n67_));
NOR2X1 NOR2X1_674 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n81_));
NOR2X1 NOR2X1_675 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n82_));
NOR2X1 NOR2X1_676 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_));
NOR2X1 NOR2X1_677 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n106_));
NOR2X1 NOR2X1_678 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n137_));
NOR2X1 NOR2X1_679 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n140_));
NOR2X1 NOR2X1_68 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3706_), .B(AES_CORE_DATAPATH__abc_15863_new_n3703_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3707_));
NOR2X1 NOR2X1_680 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n286_));
NOR2X1 NOR2X1_681 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n287_));
NOR2X1 NOR2X1_682 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n327_));
NOR2X1 NOR2X1_683 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n328_));
NOR2X1 NOR2X1_684 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n339_));
NOR2X1 NOR2X1_685 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n336_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n343_));
NOR2X1 NOR2X1_686 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n351_));
NOR2X1 NOR2X1_687 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n312_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n353_));
NOR2X1 NOR2X1_688 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n371_));
NOR2X1 NOR2X1_689 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n200_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n372_));
NOR2X1 NOR2X1_69 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3750_), .B(AES_CORE_DATAPATH__abc_15863_new_n3747_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3751_));
NOR2X1 NOR2X1_690 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n379_));
NOR2X1 NOR2X1_691 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n380_));
NOR2X1 NOR2X1_692 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n394_));
NOR2X1 NOR2X1_693 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n400_));
NOR2X1 NOR2X1_694 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n414_));
NOR2X1 NOR2X1_695 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n416_));
NOR2X1 NOR2X1_696 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n420_));
NOR2X1 NOR2X1_697 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n432_));
NOR2X1 NOR2X1_698 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n457_));
NOR2X1 NOR2X1_699 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n482_));
NOR2X1 NOR2X1_7 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n92_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n93_));
NOR2X1 NOR2X1_70 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3772_), .B(AES_CORE_DATAPATH__abc_15863_new_n3769_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3773_));
NOR2X1 NOR2X1_700 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n500_));
NOR2X1 NOR2X1_701 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n56_));
NOR2X1 NOR2X1_702 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n67_));
NOR2X1 NOR2X1_703 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n81_));
NOR2X1 NOR2X1_704 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n82_));
NOR2X1 NOR2X1_705 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_));
NOR2X1 NOR2X1_706 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n106_));
NOR2X1 NOR2X1_707 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n137_));
NOR2X1 NOR2X1_708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n140_));
NOR2X1 NOR2X1_709 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n286_));
NOR2X1 NOR2X1_71 ( .A(\key_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4033_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4034_));
NOR2X1 NOR2X1_710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n287_));
NOR2X1 NOR2X1_711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n327_));
NOR2X1 NOR2X1_712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n328_));
NOR2X1 NOR2X1_713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n339_));
NOR2X1 NOR2X1_714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n336_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n343_));
NOR2X1 NOR2X1_715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n351_));
NOR2X1 NOR2X1_716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n312_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n353_));
NOR2X1 NOR2X1_717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n371_));
NOR2X1 NOR2X1_718 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n200_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n372_));
NOR2X1 NOR2X1_719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n379_));
NOR2X1 NOR2X1_72 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4235_));
NOR2X1 NOR2X1_720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n380_));
NOR2X1 NOR2X1_721 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n394_));
NOR2X1 NOR2X1_722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n400_));
NOR2X1 NOR2X1_723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n414_));
NOR2X1 NOR2X1_724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n416_));
NOR2X1 NOR2X1_725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n420_));
NOR2X1 NOR2X1_726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n432_));
NOR2X1 NOR2X1_727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n457_));
NOR2X1 NOR2X1_728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n482_));
NOR2X1 NOR2X1_729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n500_));
NOR2X1 NOR2X1_73 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4240_));
NOR2X1 NOR2X1_730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n56_));
NOR2X1 NOR2X1_731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n67_));
NOR2X1 NOR2X1_732 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n81_));
NOR2X1 NOR2X1_733 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n82_));
NOR2X1 NOR2X1_734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_));
NOR2X1 NOR2X1_735 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n106_));
NOR2X1 NOR2X1_736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n137_));
NOR2X1 NOR2X1_737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n140_));
NOR2X1 NOR2X1_738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n286_));
NOR2X1 NOR2X1_739 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n287_));
NOR2X1 NOR2X1_74 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4245_));
NOR2X1 NOR2X1_740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n327_));
NOR2X1 NOR2X1_741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n328_));
NOR2X1 NOR2X1_742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n339_));
NOR2X1 NOR2X1_743 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n336_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n343_));
NOR2X1 NOR2X1_744 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n351_));
NOR2X1 NOR2X1_745 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n312_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n353_));
NOR2X1 NOR2X1_746 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n371_));
NOR2X1 NOR2X1_747 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n196_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n200_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n372_));
NOR2X1 NOR2X1_748 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n242_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n379_));
NOR2X1 NOR2X1_749 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n373_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n246_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n380_));
NOR2X1 NOR2X1_75 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4250_));
NOR2X1 NOR2X1_750 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n394_));
NOR2X1 NOR2X1_751 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n400_));
NOR2X1 NOR2X1_752 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n413_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n412_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n414_));
NOR2X1 NOR2X1_753 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n414_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n411_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n416_));
NOR2X1 NOR2X1_754 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n418_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n414_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n420_));
NOR2X1 NOR2X1_755 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n432_));
NOR2X1 NOR2X1_756 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n457_));
NOR2X1 NOR2X1_757 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n410_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n406_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n482_));
NOR2X1 NOR2X1_758 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n500_));
NOR2X1 NOR2X1_759 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15730_new_n71_));
NOR2X1 NOR2X1_76 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4255_));
NOR2X1 NOR2X1_760 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15730_new_n71_));
NOR2X1 NOR2X1_77 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4260_));
NOR2X1 NOR2X1_78 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4263_));
NOR2X1 NOR2X1_79 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4266_));
NOR2X1 NOR2X1_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n89_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n85_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n95_));
NOR2X1 NOR2X1_80 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4269_));
NOR2X1 NOR2X1_81 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4272_));
NOR2X1 NOR2X1_82 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4275_));
NOR2X1 NOR2X1_83 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4278_));
NOR2X1 NOR2X1_84 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4283_));
NOR2X1 NOR2X1_85 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4288_));
NOR2X1 NOR2X1_86 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4293_));
NOR2X1 NOR2X1_87 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4298_));
NOR2X1 NOR2X1_88 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4303_));
NOR2X1 NOR2X1_89 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4308_));
NOR2X1 NOR2X1_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n97_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n98_));
NOR2X1 NOR2X1_90 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4313_));
NOR2X1 NOR2X1_91 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4318_));
NOR2X1 NOR2X1_92 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4323_));
NOR2X1 NOR2X1_93 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4328_));
NOR2X1 NOR2X1_94 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4333_));
NOR2X1 NOR2X1_95 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4338_));
NOR2X1 NOR2X1_96 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4343_));
NOR2X1 NOR2X1_97 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4348_));
NOR2X1 NOR2X1_98 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4353_));
NOR2X1 NOR2X1_99 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4198_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4358_));
NOR3X1 NOR3X1_1 ( .A(\addr[1] ), .B(\addr[0] ), .C(_abc_15574_new_n11_), .Y(AES_CORE_DATAPATH_col_en_host_0_));
NOR3X1 NOR3X1_2 ( .A(\addr[0] ), .B(_abc_15574_new_n15_), .C(_abc_15574_new_n11_), .Y(AES_CORE_DATAPATH_col_en_host_2_));
NOR3X1 NOR3X1_3 ( .A(AES_CORE_DATAPATH_col_sel_host_1_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_1_), .C(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3091_));
OAI21X1 OAI21X1_1 ( .A(\aes_mode[0] ), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_), .C(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_));
OAI21X1 OAI21X1_10 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .C(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n135_));
OAI21X1 OAI21X1_100 ( .A(AES_CORE_DATAPATH_iv_2__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2657_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2658_));
OAI21X1 OAI21X1_1000 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5610_), .C(AES_CORE_DATAPATH__abc_15863_new_n5611_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5612_));
OAI21X1 OAI21X1_1001 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5610_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5615_));
OAI21X1 OAI21X1_1002 ( .A(\iv_out[26] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5615_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5616_));
OAI21X1 OAI21X1_1003 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5600_), .B(AES_CORE_DATAPATH__abc_15863_new_n5614_), .C(AES_CORE_DATAPATH__abc_15863_new_n5616_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5617_));
OAI21X1 OAI21X1_1004 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[26] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5619_));
OAI21X1 OAI21X1_1005 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5622_));
OAI21X1 OAI21X1_1006 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5622_), .B(AES_CORE_DATAPATH__abc_15863_new_n5621_), .C(AES_CORE_DATAPATH__abc_15863_new_n5623_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5624_));
OAI21X1 OAI21X1_1007 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5620_), .B(AES_CORE_DATAPATH__abc_15863_new_n5624_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5625_));
OAI21X1 OAI21X1_1008 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5629_), .C(AES_CORE_DATAPATH__abc_15863_new_n5592_), .Y(AES_CORE_DATAPATH__0col_0__31_0__26_));
OAI21X1 OAI21X1_1009 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3029_), .B(AES_CORE_DATAPATH__abc_15863_new_n3701_), .C(AES_CORE_DATAPATH__abc_15863_new_n5635_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5636_));
OAI21X1 OAI21X1_101 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2661_));
OAI21X1 OAI21X1_1010 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5641_));
OAI21X1 OAI21X1_1011 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5642_));
OAI21X1 OAI21X1_1012 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5642_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5641_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5643_));
OAI21X1 OAI21X1_1013 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5640_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5644_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5645_));
OAI21X1 OAI21X1_1014 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5646_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5647_));
OAI21X1 OAI21X1_1015 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5645_), .C(AES_CORE_DATAPATH__abc_15863_new_n5647_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5648_));
OAI21X1 OAI21X1_1016 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5648_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5649_));
OAI21X1 OAI21X1_1017 ( .A(\iv_out[27] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5649_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5650_));
OAI21X1 OAI21X1_1018 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3706_), .B(AES_CORE_DATAPATH__abc_15863_new_n3703_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5652_));
OAI21X1 OAI21X1_1019 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5648_), .C(AES_CORE_DATAPATH__abc_15863_new_n5655_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5656_));
OAI21X1 OAI21X1_102 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2661_), .C(AES_CORE_DATAPATH__abc_15863_new_n2662_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2663_));
OAI21X1 OAI21X1_1020 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[27] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5659_));
OAI21X1 OAI21X1_1021 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5662_));
OAI21X1 OAI21X1_1022 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5662_), .B(AES_CORE_DATAPATH__abc_15863_new_n5661_), .C(AES_CORE_DATAPATH__abc_15863_new_n5663_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5664_));
OAI21X1 OAI21X1_1023 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5660_), .B(AES_CORE_DATAPATH__abc_15863_new_n5664_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5665_));
OAI21X1 OAI21X1_1024 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5668_), .C(AES_CORE_DATAPATH__abc_15863_new_n5631_), .Y(AES_CORE_DATAPATH__0col_0__31_0__27_));
OAI21X1 OAI21X1_1025 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3728_), .B(AES_CORE_DATAPATH__abc_15863_new_n5676_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5677_));
OAI21X1 OAI21X1_1026 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5681_));
OAI21X1 OAI21X1_1027 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5682_));
OAI21X1 OAI21X1_1028 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5682_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5681_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5683_));
OAI21X1 OAI21X1_1029 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5680_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5684_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5685_));
OAI21X1 OAI21X1_103 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2660_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2666_), .Y(\iv_out[25] ));
OAI21X1 OAI21X1_1030 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5686_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5687_));
OAI21X1 OAI21X1_1031 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5685_), .C(AES_CORE_DATAPATH__abc_15863_new_n5687_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5688_));
OAI21X1 OAI21X1_1032 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5688_), .C(AES_CORE_DATAPATH__abc_15863_new_n5689_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5690_));
OAI21X1 OAI21X1_1033 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5688_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5693_));
OAI21X1 OAI21X1_1034 ( .A(\iv_out[28] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5693_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5694_));
OAI21X1 OAI21X1_1035 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5678_), .B(AES_CORE_DATAPATH__abc_15863_new_n5692_), .C(AES_CORE_DATAPATH__abc_15863_new_n5694_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5695_));
OAI21X1 OAI21X1_1036 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[28] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5697_));
OAI21X1 OAI21X1_1037 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5700_));
OAI21X1 OAI21X1_1038 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5700_), .B(AES_CORE_DATAPATH__abc_15863_new_n5699_), .C(AES_CORE_DATAPATH__abc_15863_new_n5701_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5702_));
OAI21X1 OAI21X1_1039 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5698_), .B(AES_CORE_DATAPATH__abc_15863_new_n5702_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5703_));
OAI21X1 OAI21X1_104 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2669_));
OAI21X1 OAI21X1_1040 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5707_), .C(AES_CORE_DATAPATH__abc_15863_new_n5670_), .Y(AES_CORE_DATAPATH__0col_0__31_0__28_));
OAI21X1 OAI21X1_1041 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3050_), .B(AES_CORE_DATAPATH__abc_15863_new_n3745_), .C(AES_CORE_DATAPATH__abc_15863_new_n5713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5714_));
OAI21X1 OAI21X1_1042 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5718_));
OAI21X1 OAI21X1_1043 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n5718_), .C(AES_CORE_DATAPATH__abc_15863_new_n5719_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5720_));
OAI21X1 OAI21X1_1044 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5723_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5724_));
OAI21X1 OAI21X1_1045 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4598_), .B(\iv_out[29] ), .C(AES_CORE_DATAPATH__abc_15863_new_n5724_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5725_));
OAI21X1 OAI21X1_1046 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3750_), .B(AES_CORE_DATAPATH__abc_15863_new_n3747_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5727_));
OAI21X1 OAI21X1_1047 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5723_), .C(AES_CORE_DATAPATH__abc_15863_new_n5730_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5731_));
OAI21X1 OAI21X1_1048 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[29] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5734_));
OAI21X1 OAI21X1_1049 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5737_));
OAI21X1 OAI21X1_105 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2669_), .C(AES_CORE_DATAPATH__abc_15863_new_n2670_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2671_));
OAI21X1 OAI21X1_1050 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5737_), .B(AES_CORE_DATAPATH__abc_15863_new_n5736_), .C(AES_CORE_DATAPATH__abc_15863_new_n5738_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5739_));
OAI21X1 OAI21X1_1051 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5735_), .B(AES_CORE_DATAPATH__abc_15863_new_n5739_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5740_));
OAI21X1 OAI21X1_1052 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5743_), .C(AES_CORE_DATAPATH__abc_15863_new_n5709_), .Y(AES_CORE_DATAPATH__0col_0__31_0__29_));
OAI21X1 OAI21X1_1053 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3060_), .B(AES_CORE_DATAPATH__abc_15863_new_n3767_), .C(AES_CORE_DATAPATH__abc_15863_new_n5749_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5750_));
OAI21X1 OAI21X1_1054 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5755_));
OAI21X1 OAI21X1_1055 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5756_));
OAI21X1 OAI21X1_1056 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5756_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5757_));
OAI21X1 OAI21X1_1057 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5754_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5758_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5759_));
OAI21X1 OAI21X1_1058 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5760_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5761_));
OAI21X1 OAI21X1_1059 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5759_), .C(AES_CORE_DATAPATH__abc_15863_new_n5761_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5762_));
OAI21X1 OAI21X1_106 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2668_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2674_), .Y(\iv_out[26] ));
OAI21X1 OAI21X1_1060 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5762_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5763_));
OAI21X1 OAI21X1_1061 ( .A(\iv_out[30] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5763_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5764_));
OAI21X1 OAI21X1_1062 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3772_), .B(AES_CORE_DATAPATH__abc_15863_new_n3769_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5766_));
OAI21X1 OAI21X1_1063 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5762_), .C(AES_CORE_DATAPATH__abc_15863_new_n5769_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5770_));
OAI21X1 OAI21X1_1064 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[30] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5773_));
OAI21X1 OAI21X1_1065 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5776_));
OAI21X1 OAI21X1_1066 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5776_), .B(AES_CORE_DATAPATH__abc_15863_new_n5775_), .C(AES_CORE_DATAPATH__abc_15863_new_n5777_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5778_));
OAI21X1 OAI21X1_1067 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5774_), .B(AES_CORE_DATAPATH__abc_15863_new_n5778_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5779_));
OAI21X1 OAI21X1_1068 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5782_), .C(AES_CORE_DATAPATH__abc_15863_new_n5745_), .Y(AES_CORE_DATAPATH__0col_0__31_0__30_));
OAI21X1 OAI21X1_1069 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3794_), .B(AES_CORE_DATAPATH__abc_15863_new_n5790_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5791_));
OAI21X1 OAI21X1_107 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2677_));
OAI21X1 OAI21X1_1070 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5795_));
OAI21X1 OAI21X1_1071 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5796_));
OAI21X1 OAI21X1_1072 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5796_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5795_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5797_));
OAI21X1 OAI21X1_1073 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5794_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5798_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5799_));
OAI21X1 OAI21X1_1074 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5800_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5801_));
OAI21X1 OAI21X1_1075 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5799_), .C(AES_CORE_DATAPATH__abc_15863_new_n5801_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5802_));
OAI21X1 OAI21X1_1076 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5802_), .C(AES_CORE_DATAPATH__abc_15863_new_n5803_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5804_));
OAI21X1 OAI21X1_1077 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5802_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5807_));
OAI21X1 OAI21X1_1078 ( .A(\iv_out[31] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5807_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5808_));
OAI21X1 OAI21X1_1079 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5792_), .B(AES_CORE_DATAPATH__abc_15863_new_n5806_), .C(AES_CORE_DATAPATH__abc_15863_new_n5808_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5809_));
OAI21X1 OAI21X1_108 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2677_), .C(AES_CORE_DATAPATH__abc_15863_new_n2678_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2679_));
OAI21X1 OAI21X1_1080 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[31] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5811_));
OAI21X1 OAI21X1_1081 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5814_));
OAI21X1 OAI21X1_1082 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5814_), .B(AES_CORE_DATAPATH__abc_15863_new_n5813_), .C(AES_CORE_DATAPATH__abc_15863_new_n5815_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5816_));
OAI21X1 OAI21X1_1083 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5812_), .B(AES_CORE_DATAPATH__abc_15863_new_n5816_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5817_));
OAI21X1 OAI21X1_1084 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5821_), .C(AES_CORE_DATAPATH__abc_15863_new_n5784_), .Y(AES_CORE_DATAPATH__0col_0__31_0__31_));
OAI21X1 OAI21X1_1085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5827_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5828_));
OAI21X1 OAI21X1_1086 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5828_), .C(AES_CORE_DATAPATH__abc_15863_new_n5829_), .Y(AES_CORE_DATAPATH__0key_3__31_0__0_));
OAI21X1 OAI21X1_1087 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5832_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5833_));
OAI21X1 OAI21X1_1088 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5833_), .C(AES_CORE_DATAPATH__abc_15863_new_n5834_), .Y(AES_CORE_DATAPATH__0key_3__31_0__1_));
OAI21X1 OAI21X1_1089 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5837_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5838_));
OAI21X1 OAI21X1_109 ( .A(AES_CORE_DATAPATH_iv_2__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2679_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2680_));
OAI21X1 OAI21X1_1090 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5838_), .C(AES_CORE_DATAPATH__abc_15863_new_n5839_), .Y(AES_CORE_DATAPATH__0key_3__31_0__2_));
OAI21X1 OAI21X1_1091 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5842_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5843_));
OAI21X1 OAI21X1_1092 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5843_), .C(AES_CORE_DATAPATH__abc_15863_new_n5844_), .Y(AES_CORE_DATAPATH__0key_3__31_0__3_));
OAI21X1 OAI21X1_1093 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5847_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5848_));
OAI21X1 OAI21X1_1094 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5848_), .C(AES_CORE_DATAPATH__abc_15863_new_n5849_), .Y(AES_CORE_DATAPATH__0key_3__31_0__4_));
OAI21X1 OAI21X1_1095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5852_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5853_));
OAI21X1 OAI21X1_1096 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5853_), .C(AES_CORE_DATAPATH__abc_15863_new_n5854_), .Y(AES_CORE_DATAPATH__0key_3__31_0__5_));
OAI21X1 OAI21X1_1097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5857_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5858_));
OAI21X1 OAI21X1_1098 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5858_), .C(AES_CORE_DATAPATH__abc_15863_new_n5859_), .Y(AES_CORE_DATAPATH__0key_3__31_0__6_));
OAI21X1 OAI21X1_1099 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5862_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5863_));
OAI21X1 OAI21X1_11 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n83_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n139_));
OAI21X1 OAI21X1_110 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2683_));
OAI21X1 OAI21X1_1100 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5863_), .C(AES_CORE_DATAPATH__abc_15863_new_n5864_), .Y(AES_CORE_DATAPATH__0key_3__31_0__7_));
OAI21X1 OAI21X1_1101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5867_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5868_));
OAI21X1 OAI21X1_1102 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5868_), .C(AES_CORE_DATAPATH__abc_15863_new_n5869_), .Y(AES_CORE_DATAPATH__0key_3__31_0__8_));
OAI21X1 OAI21X1_1103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5872_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5873_));
OAI21X1 OAI21X1_1104 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5873_), .C(AES_CORE_DATAPATH__abc_15863_new_n5874_), .Y(AES_CORE_DATAPATH__0key_3__31_0__9_));
OAI21X1 OAI21X1_1105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5877_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5878_));
OAI21X1 OAI21X1_1106 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5878_), .C(AES_CORE_DATAPATH__abc_15863_new_n5879_), .Y(AES_CORE_DATAPATH__0key_3__31_0__10_));
OAI21X1 OAI21X1_1107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5882_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5883_));
OAI21X1 OAI21X1_1108 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5883_), .C(AES_CORE_DATAPATH__abc_15863_new_n5884_), .Y(AES_CORE_DATAPATH__0key_3__31_0__11_));
OAI21X1 OAI21X1_1109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5887_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5888_));
OAI21X1 OAI21X1_111 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2683_), .C(AES_CORE_DATAPATH__abc_15863_new_n2684_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2685_));
OAI21X1 OAI21X1_1110 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5888_), .C(AES_CORE_DATAPATH__abc_15863_new_n5889_), .Y(AES_CORE_DATAPATH__0key_3__31_0__12_));
OAI21X1 OAI21X1_1111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5892_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5893_));
OAI21X1 OAI21X1_1112 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5893_), .C(AES_CORE_DATAPATH__abc_15863_new_n5894_), .Y(AES_CORE_DATAPATH__0key_3__31_0__13_));
OAI21X1 OAI21X1_1113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5897_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5898_));
OAI21X1 OAI21X1_1114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5898_), .C(AES_CORE_DATAPATH__abc_15863_new_n5899_), .Y(AES_CORE_DATAPATH__0key_3__31_0__14_));
OAI21X1 OAI21X1_1115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5902_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5903_));
OAI21X1 OAI21X1_1116 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5903_), .C(AES_CORE_DATAPATH__abc_15863_new_n5904_), .Y(AES_CORE_DATAPATH__0key_3__31_0__15_));
OAI21X1 OAI21X1_1117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5907_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5908_));
OAI21X1 OAI21X1_1118 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5908_), .C(AES_CORE_DATAPATH__abc_15863_new_n5909_), .Y(AES_CORE_DATAPATH__0key_3__31_0__16_));
OAI21X1 OAI21X1_1119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5912_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5913_));
OAI21X1 OAI21X1_112 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2682_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2688_), .Y(\iv_out[28] ));
OAI21X1 OAI21X1_1120 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5913_), .C(AES_CORE_DATAPATH__abc_15863_new_n5914_), .Y(AES_CORE_DATAPATH__0key_3__31_0__17_));
OAI21X1 OAI21X1_1121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5917_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5918_));
OAI21X1 OAI21X1_1122 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5918_), .C(AES_CORE_DATAPATH__abc_15863_new_n5919_), .Y(AES_CORE_DATAPATH__0key_3__31_0__18_));
OAI21X1 OAI21X1_1123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5922_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5923_));
OAI21X1 OAI21X1_1124 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5923_), .C(AES_CORE_DATAPATH__abc_15863_new_n5924_), .Y(AES_CORE_DATAPATH__0key_3__31_0__19_));
OAI21X1 OAI21X1_1125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5927_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5928_));
OAI21X1 OAI21X1_1126 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5928_), .C(AES_CORE_DATAPATH__abc_15863_new_n5929_), .Y(AES_CORE_DATAPATH__0key_3__31_0__20_));
OAI21X1 OAI21X1_1127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5932_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5933_));
OAI21X1 OAI21X1_1128 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5933_), .C(AES_CORE_DATAPATH__abc_15863_new_n5934_), .Y(AES_CORE_DATAPATH__0key_3__31_0__21_));
OAI21X1 OAI21X1_1129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5937_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5938_));
OAI21X1 OAI21X1_113 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2691_));
OAI21X1 OAI21X1_1130 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5938_), .C(AES_CORE_DATAPATH__abc_15863_new_n5939_), .Y(AES_CORE_DATAPATH__0key_3__31_0__22_));
OAI21X1 OAI21X1_1131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5942_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5943_));
OAI21X1 OAI21X1_1132 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5943_), .C(AES_CORE_DATAPATH__abc_15863_new_n5944_), .Y(AES_CORE_DATAPATH__0key_3__31_0__23_));
OAI21X1 OAI21X1_1133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5947_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5948_));
OAI21X1 OAI21X1_1134 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5948_), .C(AES_CORE_DATAPATH__abc_15863_new_n5949_), .Y(AES_CORE_DATAPATH__0key_3__31_0__24_));
OAI21X1 OAI21X1_1135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5952_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5953_));
OAI21X1 OAI21X1_1136 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5953_), .C(AES_CORE_DATAPATH__abc_15863_new_n5954_), .Y(AES_CORE_DATAPATH__0key_3__31_0__25_));
OAI21X1 OAI21X1_1137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5957_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5958_));
OAI21X1 OAI21X1_1138 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5958_), .C(AES_CORE_DATAPATH__abc_15863_new_n5959_), .Y(AES_CORE_DATAPATH__0key_3__31_0__26_));
OAI21X1 OAI21X1_1139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5962_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5963_));
OAI21X1 OAI21X1_114 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2691_), .C(AES_CORE_DATAPATH__abc_15863_new_n2692_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2693_));
OAI21X1 OAI21X1_1140 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5963_), .C(AES_CORE_DATAPATH__abc_15863_new_n5964_), .Y(AES_CORE_DATAPATH__0key_3__31_0__27_));
OAI21X1 OAI21X1_1141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5967_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5968_));
OAI21X1 OAI21X1_1142 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5968_), .C(AES_CORE_DATAPATH__abc_15863_new_n5969_), .Y(AES_CORE_DATAPATH__0key_3__31_0__28_));
OAI21X1 OAI21X1_1143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5972_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5973_));
OAI21X1 OAI21X1_1144 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5973_), .C(AES_CORE_DATAPATH__abc_15863_new_n5974_), .Y(AES_CORE_DATAPATH__0key_3__31_0__29_));
OAI21X1 OAI21X1_1145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5977_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5978_));
OAI21X1 OAI21X1_1146 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5978_), .C(AES_CORE_DATAPATH__abc_15863_new_n5979_), .Y(AES_CORE_DATAPATH__0key_3__31_0__30_));
OAI21X1 OAI21X1_1147 ( .A(\key_en[3] ), .B(AES_CORE_DATAPATH_key_host_3__31_), .C(AES_CORE_DATAPATH__abc_15863_new_n5981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5982_));
OAI21X1 OAI21X1_1148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n5983_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5984_));
OAI21X1 OAI21X1_1149 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5825_), .B(AES_CORE_DATAPATH__abc_15863_new_n5984_), .C(AES_CORE_DATAPATH__abc_15863_new_n5985_), .Y(AES_CORE_DATAPATH__0key_3__31_0__31_));
OAI21X1 OAI21X1_115 ( .A(AES_CORE_DATAPATH_iv_2__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2693_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2694_));
OAI21X1 OAI21X1_1150 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .B(AES_CORE_DATAPATH__abc_15863_new_n5826_), .C(AES_CORE_DATAPATH__abc_15863_new_n5987_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__0_));
OAI21X1 OAI21X1_1151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6056_), .C(AES_CORE_DATAPATH__abc_15863_new_n6051_), .Y(AES_CORE_DATAPATH__0col_3__31_0__0_));
OAI21X1 OAI21X1_1152 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6063_), .C(AES_CORE_DATAPATH__abc_15863_new_n6058_), .Y(AES_CORE_DATAPATH__0col_3__31_0__1_));
OAI21X1 OAI21X1_1153 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6070_), .C(AES_CORE_DATAPATH__abc_15863_new_n6065_), .Y(AES_CORE_DATAPATH__0col_3__31_0__2_));
OAI21X1 OAI21X1_1154 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6077_), .C(AES_CORE_DATAPATH__abc_15863_new_n6072_), .Y(AES_CORE_DATAPATH__0col_3__31_0__3_));
OAI21X1 OAI21X1_1155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6084_), .C(AES_CORE_DATAPATH__abc_15863_new_n6079_), .Y(AES_CORE_DATAPATH__0col_3__31_0__4_));
OAI21X1 OAI21X1_1156 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6091_), .C(AES_CORE_DATAPATH__abc_15863_new_n6086_), .Y(AES_CORE_DATAPATH__0col_3__31_0__5_));
OAI21X1 OAI21X1_1157 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6098_), .C(AES_CORE_DATAPATH__abc_15863_new_n6093_), .Y(AES_CORE_DATAPATH__0col_3__31_0__6_));
OAI21X1 OAI21X1_1158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6105_), .C(AES_CORE_DATAPATH__abc_15863_new_n6100_), .Y(AES_CORE_DATAPATH__0col_3__31_0__7_));
OAI21X1 OAI21X1_1159 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6112_), .C(AES_CORE_DATAPATH__abc_15863_new_n6107_), .Y(AES_CORE_DATAPATH__0col_3__31_0__8_));
OAI21X1 OAI21X1_116 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2697_));
OAI21X1 OAI21X1_1160 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6119_), .C(AES_CORE_DATAPATH__abc_15863_new_n6114_), .Y(AES_CORE_DATAPATH__0col_3__31_0__9_));
OAI21X1 OAI21X1_1161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6126_), .C(AES_CORE_DATAPATH__abc_15863_new_n6121_), .Y(AES_CORE_DATAPATH__0col_3__31_0__10_));
OAI21X1 OAI21X1_1162 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6133_), .C(AES_CORE_DATAPATH__abc_15863_new_n6128_), .Y(AES_CORE_DATAPATH__0col_3__31_0__11_));
OAI21X1 OAI21X1_1163 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6140_), .C(AES_CORE_DATAPATH__abc_15863_new_n6135_), .Y(AES_CORE_DATAPATH__0col_3__31_0__12_));
OAI21X1 OAI21X1_1164 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6147_), .C(AES_CORE_DATAPATH__abc_15863_new_n6142_), .Y(AES_CORE_DATAPATH__0col_3__31_0__13_));
OAI21X1 OAI21X1_1165 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6154_), .C(AES_CORE_DATAPATH__abc_15863_new_n6149_), .Y(AES_CORE_DATAPATH__0col_3__31_0__14_));
OAI21X1 OAI21X1_1166 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6161_), .C(AES_CORE_DATAPATH__abc_15863_new_n6156_), .Y(AES_CORE_DATAPATH__0col_3__31_0__15_));
OAI21X1 OAI21X1_1167 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6168_), .C(AES_CORE_DATAPATH__abc_15863_new_n6163_), .Y(AES_CORE_DATAPATH__0col_3__31_0__16_));
OAI21X1 OAI21X1_1168 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6175_), .C(AES_CORE_DATAPATH__abc_15863_new_n6170_), .Y(AES_CORE_DATAPATH__0col_3__31_0__17_));
OAI21X1 OAI21X1_1169 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6182_), .C(AES_CORE_DATAPATH__abc_15863_new_n6177_), .Y(AES_CORE_DATAPATH__0col_3__31_0__18_));
OAI21X1 OAI21X1_117 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2697_), .C(AES_CORE_DATAPATH__abc_15863_new_n2698_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2699_));
OAI21X1 OAI21X1_1170 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6189_), .C(AES_CORE_DATAPATH__abc_15863_new_n6184_), .Y(AES_CORE_DATAPATH__0col_3__31_0__19_));
OAI21X1 OAI21X1_1171 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6196_), .C(AES_CORE_DATAPATH__abc_15863_new_n6191_), .Y(AES_CORE_DATAPATH__0col_3__31_0__20_));
OAI21X1 OAI21X1_1172 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6203_), .C(AES_CORE_DATAPATH__abc_15863_new_n6198_), .Y(AES_CORE_DATAPATH__0col_3__31_0__21_));
OAI21X1 OAI21X1_1173 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6210_), .C(AES_CORE_DATAPATH__abc_15863_new_n6205_), .Y(AES_CORE_DATAPATH__0col_3__31_0__22_));
OAI21X1 OAI21X1_1174 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6217_), .C(AES_CORE_DATAPATH__abc_15863_new_n6212_), .Y(AES_CORE_DATAPATH__0col_3__31_0__23_));
OAI21X1 OAI21X1_1175 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6224_), .C(AES_CORE_DATAPATH__abc_15863_new_n6219_), .Y(AES_CORE_DATAPATH__0col_3__31_0__24_));
OAI21X1 OAI21X1_1176 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6231_), .C(AES_CORE_DATAPATH__abc_15863_new_n6226_), .Y(AES_CORE_DATAPATH__0col_3__31_0__25_));
OAI21X1 OAI21X1_1177 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6238_), .C(AES_CORE_DATAPATH__abc_15863_new_n6233_), .Y(AES_CORE_DATAPATH__0col_3__31_0__26_));
OAI21X1 OAI21X1_1178 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6245_), .C(AES_CORE_DATAPATH__abc_15863_new_n6240_), .Y(AES_CORE_DATAPATH__0col_3__31_0__27_));
OAI21X1 OAI21X1_1179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6252_), .C(AES_CORE_DATAPATH__abc_15863_new_n6247_), .Y(AES_CORE_DATAPATH__0col_3__31_0__28_));
OAI21X1 OAI21X1_118 ( .A(AES_CORE_DATAPATH_iv_2__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2699_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2700_));
OAI21X1 OAI21X1_1180 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6259_), .C(AES_CORE_DATAPATH__abc_15863_new_n6254_), .Y(AES_CORE_DATAPATH__0col_3__31_0__29_));
OAI21X1 OAI21X1_1181 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6266_), .C(AES_CORE_DATAPATH__abc_15863_new_n6261_), .Y(AES_CORE_DATAPATH__0col_3__31_0__30_));
OAI21X1 OAI21X1_1182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2461_), .B(AES_CORE_DATAPATH__abc_15863_new_n6273_), .C(AES_CORE_DATAPATH__abc_15863_new_n6268_), .Y(AES_CORE_DATAPATH__0col_3__31_0__31_));
OAI21X1 OAI21X1_1183 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6280_), .C(AES_CORE_DATAPATH__abc_15863_new_n6275_), .Y(AES_CORE_DATAPATH__0col_1__31_0__0_));
OAI21X1 OAI21X1_1184 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6287_), .C(AES_CORE_DATAPATH__abc_15863_new_n6282_), .Y(AES_CORE_DATAPATH__0col_1__31_0__1_));
OAI21X1 OAI21X1_1185 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6294_), .C(AES_CORE_DATAPATH__abc_15863_new_n6289_), .Y(AES_CORE_DATAPATH__0col_1__31_0__2_));
OAI21X1 OAI21X1_1186 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6301_), .C(AES_CORE_DATAPATH__abc_15863_new_n6296_), .Y(AES_CORE_DATAPATH__0col_1__31_0__3_));
OAI21X1 OAI21X1_1187 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6308_), .C(AES_CORE_DATAPATH__abc_15863_new_n6303_), .Y(AES_CORE_DATAPATH__0col_1__31_0__4_));
OAI21X1 OAI21X1_1188 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6315_), .C(AES_CORE_DATAPATH__abc_15863_new_n6310_), .Y(AES_CORE_DATAPATH__0col_1__31_0__5_));
OAI21X1 OAI21X1_1189 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6322_), .C(AES_CORE_DATAPATH__abc_15863_new_n6317_), .Y(AES_CORE_DATAPATH__0col_1__31_0__6_));
OAI21X1 OAI21X1_119 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2703_));
OAI21X1 OAI21X1_1190 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6329_), .C(AES_CORE_DATAPATH__abc_15863_new_n6324_), .Y(AES_CORE_DATAPATH__0col_1__31_0__7_));
OAI21X1 OAI21X1_1191 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6336_), .C(AES_CORE_DATAPATH__abc_15863_new_n6331_), .Y(AES_CORE_DATAPATH__0col_1__31_0__8_));
OAI21X1 OAI21X1_1192 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6343_), .C(AES_CORE_DATAPATH__abc_15863_new_n6338_), .Y(AES_CORE_DATAPATH__0col_1__31_0__9_));
OAI21X1 OAI21X1_1193 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6350_), .C(AES_CORE_DATAPATH__abc_15863_new_n6345_), .Y(AES_CORE_DATAPATH__0col_1__31_0__10_));
OAI21X1 OAI21X1_1194 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6357_), .C(AES_CORE_DATAPATH__abc_15863_new_n6352_), .Y(AES_CORE_DATAPATH__0col_1__31_0__11_));
OAI21X1 OAI21X1_1195 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6364_), .C(AES_CORE_DATAPATH__abc_15863_new_n6359_), .Y(AES_CORE_DATAPATH__0col_1__31_0__12_));
OAI21X1 OAI21X1_1196 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6371_), .C(AES_CORE_DATAPATH__abc_15863_new_n6366_), .Y(AES_CORE_DATAPATH__0col_1__31_0__13_));
OAI21X1 OAI21X1_1197 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6378_), .C(AES_CORE_DATAPATH__abc_15863_new_n6373_), .Y(AES_CORE_DATAPATH__0col_1__31_0__14_));
OAI21X1 OAI21X1_1198 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6385_), .C(AES_CORE_DATAPATH__abc_15863_new_n6380_), .Y(AES_CORE_DATAPATH__0col_1__31_0__15_));
OAI21X1 OAI21X1_1199 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6392_), .C(AES_CORE_DATAPATH__abc_15863_new_n6387_), .Y(AES_CORE_DATAPATH__0col_1__31_0__16_));
OAI21X1 OAI21X1_12 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n146_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n148_));
OAI21X1 OAI21X1_120 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2703_), .C(AES_CORE_DATAPATH__abc_15863_new_n2704_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2705_));
OAI21X1 OAI21X1_1200 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6399_), .C(AES_CORE_DATAPATH__abc_15863_new_n6394_), .Y(AES_CORE_DATAPATH__0col_1__31_0__17_));
OAI21X1 OAI21X1_1201 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6406_), .C(AES_CORE_DATAPATH__abc_15863_new_n6401_), .Y(AES_CORE_DATAPATH__0col_1__31_0__18_));
OAI21X1 OAI21X1_1202 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6413_), .C(AES_CORE_DATAPATH__abc_15863_new_n6408_), .Y(AES_CORE_DATAPATH__0col_1__31_0__19_));
OAI21X1 OAI21X1_1203 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6420_), .C(AES_CORE_DATAPATH__abc_15863_new_n6415_), .Y(AES_CORE_DATAPATH__0col_1__31_0__20_));
OAI21X1 OAI21X1_1204 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6427_), .C(AES_CORE_DATAPATH__abc_15863_new_n6422_), .Y(AES_CORE_DATAPATH__0col_1__31_0__21_));
OAI21X1 OAI21X1_1205 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6434_), .C(AES_CORE_DATAPATH__abc_15863_new_n6429_), .Y(AES_CORE_DATAPATH__0col_1__31_0__22_));
OAI21X1 OAI21X1_1206 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6441_), .C(AES_CORE_DATAPATH__abc_15863_new_n6436_), .Y(AES_CORE_DATAPATH__0col_1__31_0__23_));
OAI21X1 OAI21X1_1207 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6448_), .C(AES_CORE_DATAPATH__abc_15863_new_n6443_), .Y(AES_CORE_DATAPATH__0col_1__31_0__24_));
OAI21X1 OAI21X1_1208 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6455_), .C(AES_CORE_DATAPATH__abc_15863_new_n6450_), .Y(AES_CORE_DATAPATH__0col_1__31_0__25_));
OAI21X1 OAI21X1_1209 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6462_), .C(AES_CORE_DATAPATH__abc_15863_new_n6457_), .Y(AES_CORE_DATAPATH__0col_1__31_0__26_));
OAI21X1 OAI21X1_121 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2702_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2708_), .Y(\iv_out[31] ));
OAI21X1 OAI21X1_1210 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6469_), .C(AES_CORE_DATAPATH__abc_15863_new_n6464_), .Y(AES_CORE_DATAPATH__0col_1__31_0__27_));
OAI21X1 OAI21X1_1211 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6476_), .C(AES_CORE_DATAPATH__abc_15863_new_n6471_), .Y(AES_CORE_DATAPATH__0col_1__31_0__28_));
OAI21X1 OAI21X1_1212 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6483_), .C(AES_CORE_DATAPATH__abc_15863_new_n6478_), .Y(AES_CORE_DATAPATH__0col_1__31_0__29_));
OAI21X1 OAI21X1_1213 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6490_), .C(AES_CORE_DATAPATH__abc_15863_new_n6485_), .Y(AES_CORE_DATAPATH__0col_1__31_0__30_));
OAI21X1 OAI21X1_1214 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2474_), .B(AES_CORE_DATAPATH__abc_15863_new_n6497_), .C(AES_CORE_DATAPATH__abc_15863_new_n6492_), .Y(AES_CORE_DATAPATH__0col_1__31_0__31_));
OAI21X1 OAI21X1_1215 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6505_), .C(AES_CORE_DATAPATH__abc_15863_new_n6500_), .Y(AES_CORE_DATAPATH__0col_2__31_0__0_));
OAI21X1 OAI21X1_1216 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3116_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6511_), .Y(AES_CORE_DATAPATH__0col_2__31_0__1_));
OAI21X1 OAI21X1_1217 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6518_), .C(AES_CORE_DATAPATH__abc_15863_new_n6513_), .Y(AES_CORE_DATAPATH__0col_2__31_0__2_));
OAI21X1 OAI21X1_1218 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3161_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6524_), .Y(AES_CORE_DATAPATH__0col_2__31_0__3_));
OAI21X1 OAI21X1_1219 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6531_), .C(AES_CORE_DATAPATH__abc_15863_new_n6526_), .Y(AES_CORE_DATAPATH__0col_2__31_0__4_));
OAI21X1 OAI21X1_122 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH__abc_15863_new_n2713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2714_));
OAI21X1 OAI21X1_1220 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6538_), .C(AES_CORE_DATAPATH__abc_15863_new_n6533_), .Y(AES_CORE_DATAPATH__0col_2__31_0__5_));
OAI21X1 OAI21X1_1221 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6545_), .C(AES_CORE_DATAPATH__abc_15863_new_n6540_), .Y(AES_CORE_DATAPATH__0col_2__31_0__6_));
OAI21X1 OAI21X1_1222 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3250_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6551_), .Y(AES_CORE_DATAPATH__0col_2__31_0__7_));
OAI21X1 OAI21X1_1223 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6558_), .C(AES_CORE_DATAPATH__abc_15863_new_n6553_), .Y(AES_CORE_DATAPATH__0col_2__31_0__8_));
OAI21X1 OAI21X1_1224 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3294_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6564_), .Y(AES_CORE_DATAPATH__0col_2__31_0__9_));
OAI21X1 OAI21X1_1225 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6571_), .C(AES_CORE_DATAPATH__abc_15863_new_n6566_), .Y(AES_CORE_DATAPATH__0col_2__31_0__10_));
OAI21X1 OAI21X1_1226 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3338_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6577_), .Y(AES_CORE_DATAPATH__0col_2__31_0__11_));
OAI21X1 OAI21X1_1227 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6584_), .C(AES_CORE_DATAPATH__abc_15863_new_n6579_), .Y(AES_CORE_DATAPATH__0col_2__31_0__12_));
OAI21X1 OAI21X1_1228 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3382_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6590_), .Y(AES_CORE_DATAPATH__0col_2__31_0__13_));
OAI21X1 OAI21X1_1229 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6597_), .C(AES_CORE_DATAPATH__abc_15863_new_n6592_), .Y(AES_CORE_DATAPATH__0col_2__31_0__14_));
OAI21X1 OAI21X1_123 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH__abc_15863_new_n2722_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2723_));
OAI21X1 OAI21X1_1230 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3426_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6603_), .Y(AES_CORE_DATAPATH__0col_2__31_0__15_));
OAI21X1 OAI21X1_1231 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6610_), .C(AES_CORE_DATAPATH__abc_15863_new_n6605_), .Y(AES_CORE_DATAPATH__0col_2__31_0__16_));
OAI21X1 OAI21X1_1232 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3470_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6616_), .Y(AES_CORE_DATAPATH__0col_2__31_0__17_));
OAI21X1 OAI21X1_1233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3492_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6622_), .Y(AES_CORE_DATAPATH__0col_2__31_0__18_));
OAI21X1 OAI21X1_1234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3514_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6628_), .Y(AES_CORE_DATAPATH__0col_2__31_0__19_));
OAI21X1 OAI21X1_1235 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6635_), .C(AES_CORE_DATAPATH__abc_15863_new_n6630_), .Y(AES_CORE_DATAPATH__0col_2__31_0__20_));
OAI21X1 OAI21X1_1236 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3558_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6641_), .Y(AES_CORE_DATAPATH__0col_2__31_0__21_));
OAI21X1 OAI21X1_1237 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6648_), .C(AES_CORE_DATAPATH__abc_15863_new_n6643_), .Y(AES_CORE_DATAPATH__0col_2__31_0__22_));
OAI21X1 OAI21X1_1238 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3602_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6654_), .Y(AES_CORE_DATAPATH__0col_2__31_0__23_));
OAI21X1 OAI21X1_1239 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6661_), .C(AES_CORE_DATAPATH__abc_15863_new_n6656_), .Y(AES_CORE_DATAPATH__0col_2__31_0__24_));
OAI21X1 OAI21X1_124 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2732_));
OAI21X1 OAI21X1_1240 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3646_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6667_), .Y(AES_CORE_DATAPATH__0col_2__31_0__25_));
OAI21X1 OAI21X1_1241 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3668_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6673_), .Y(AES_CORE_DATAPATH__0col_2__31_0__26_));
OAI21X1 OAI21X1_1242 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6680_), .C(AES_CORE_DATAPATH__abc_15863_new_n6675_), .Y(AES_CORE_DATAPATH__0col_2__31_0__27_));
OAI21X1 OAI21X1_1243 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3712_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6686_), .Y(AES_CORE_DATAPATH__0col_2__31_0__28_));
OAI21X1 OAI21X1_1244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6693_), .C(AES_CORE_DATAPATH__abc_15863_new_n6688_), .Y(AES_CORE_DATAPATH__0col_2__31_0__29_));
OAI21X1 OAI21X1_1245 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6499_), .B(AES_CORE_DATAPATH__abc_15863_new_n6700_), .C(AES_CORE_DATAPATH__abc_15863_new_n6695_), .Y(AES_CORE_DATAPATH__0col_2__31_0__30_));
OAI21X1 OAI21X1_1246 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3778_), .B(AES_CORE_DATAPATH__abc_15863_new_n2466_), .C(AES_CORE_DATAPATH__abc_15863_new_n6706_), .Y(AES_CORE_DATAPATH__0col_2__31_0__31_));
OAI21X1 OAI21X1_1247 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n6708_), .C(AES_CORE_DATAPATH__abc_15863_new_n2716_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6709_));
OAI21X1 OAI21X1_1248 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4631_), .C(AES_CORE_DATAPATH__abc_15863_new_n6714_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__0_));
OAI21X1 OAI21X1_1249 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4670_), .C(AES_CORE_DATAPATH__abc_15863_new_n6716_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__1_));
OAI21X1 OAI21X1_125 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2717_), .B(AES_CORE_DATAPATH__abc_15863_new_n2710_), .C(AES_CORE_DATAPATH__abc_15863_new_n2732_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2733_));
OAI21X1 OAI21X1_1250 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4709_), .C(AES_CORE_DATAPATH__abc_15863_new_n6718_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__2_));
OAI21X1 OAI21X1_1251 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4749_), .C(AES_CORE_DATAPATH__abc_15863_new_n6720_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__3_));
OAI21X1 OAI21X1_1252 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4785_), .C(AES_CORE_DATAPATH__abc_15863_new_n6722_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__4_));
OAI21X1 OAI21X1_1253 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4824_), .C(AES_CORE_DATAPATH__abc_15863_new_n6724_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__5_));
OAI21X1 OAI21X1_1254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4859_), .C(AES_CORE_DATAPATH__abc_15863_new_n6726_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__6_));
OAI21X1 OAI21X1_1255 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4898_), .C(AES_CORE_DATAPATH__abc_15863_new_n6728_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__7_));
OAI21X1 OAI21X1_1256 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4933_), .C(AES_CORE_DATAPATH__abc_15863_new_n6730_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__8_));
OAI21X1 OAI21X1_1257 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n4972_), .C(AES_CORE_DATAPATH__abc_15863_new_n6732_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__9_));
OAI21X1 OAI21X1_1258 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5011_), .C(AES_CORE_DATAPATH__abc_15863_new_n6734_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__10_));
OAI21X1 OAI21X1_1259 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5050_), .C(AES_CORE_DATAPATH__abc_15863_new_n6736_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__11_));
OAI21X1 OAI21X1_126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2738_));
OAI21X1 OAI21X1_1260 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5089_), .C(AES_CORE_DATAPATH__abc_15863_new_n6738_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__12_));
OAI21X1 OAI21X1_1261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5128_), .C(AES_CORE_DATAPATH__abc_15863_new_n6740_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__13_));
OAI21X1 OAI21X1_1262 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5164_), .C(AES_CORE_DATAPATH__abc_15863_new_n6742_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__14_));
OAI21X1 OAI21X1_1263 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5203_), .C(AES_CORE_DATAPATH__abc_15863_new_n6744_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__15_));
OAI21X1 OAI21X1_1264 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5242_), .C(AES_CORE_DATAPATH__abc_15863_new_n6746_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__16_));
OAI21X1 OAI21X1_1265 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5281_), .C(AES_CORE_DATAPATH__abc_15863_new_n6748_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__17_));
OAI21X1 OAI21X1_1266 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5320_), .C(AES_CORE_DATAPATH__abc_15863_new_n6750_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__18_));
OAI21X1 OAI21X1_1267 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5359_), .C(AES_CORE_DATAPATH__abc_15863_new_n6752_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__19_));
OAI21X1 OAI21X1_1268 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5398_), .C(AES_CORE_DATAPATH__abc_15863_new_n6754_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__20_));
OAI21X1 OAI21X1_1269 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5437_), .C(AES_CORE_DATAPATH__abc_15863_new_n6756_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__21_));
OAI21X1 OAI21X1_127 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2742_));
OAI21X1 OAI21X1_1270 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5473_), .C(AES_CORE_DATAPATH__abc_15863_new_n6758_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__22_));
OAI21X1 OAI21X1_1271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5512_), .C(AES_CORE_DATAPATH__abc_15863_new_n6760_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__23_));
OAI21X1 OAI21X1_1272 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5551_), .C(AES_CORE_DATAPATH__abc_15863_new_n6762_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__24_));
OAI21X1 OAI21X1_1273 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5590_), .C(AES_CORE_DATAPATH__abc_15863_new_n6764_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__25_));
OAI21X1 OAI21X1_1274 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5629_), .C(AES_CORE_DATAPATH__abc_15863_new_n6766_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__26_));
OAI21X1 OAI21X1_1275 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5668_), .C(AES_CORE_DATAPATH__abc_15863_new_n6768_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__27_));
OAI21X1 OAI21X1_1276 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5707_), .C(AES_CORE_DATAPATH__abc_15863_new_n6770_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__28_));
OAI21X1 OAI21X1_1277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5743_), .C(AES_CORE_DATAPATH__abc_15863_new_n6772_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__29_));
OAI21X1 OAI21X1_1278 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5782_), .C(AES_CORE_DATAPATH__abc_15863_new_n6774_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__30_));
OAI21X1 OAI21X1_1279 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6713_), .B(AES_CORE_DATAPATH__abc_15863_new_n5821_), .C(AES_CORE_DATAPATH__abc_15863_new_n6776_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__31_));
OAI21X1 OAI21X1_128 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2741_), .C(AES_CORE_DATAPATH__abc_15863_new_n2742_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__0_));
OAI21X1 OAI21X1_1280 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4630_), .C(AES_CORE_DATAPATH__abc_15863_new_n6780_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6781_));
OAI21X1 OAI21X1_1281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4669_), .C(AES_CORE_DATAPATH__abc_15863_new_n6786_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6787_));
OAI21X1 OAI21X1_1282 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4708_), .C(AES_CORE_DATAPATH__abc_15863_new_n6792_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6793_));
OAI21X1 OAI21X1_1283 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4748_), .C(AES_CORE_DATAPATH__abc_15863_new_n6798_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6799_));
OAI21X1 OAI21X1_1284 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4784_), .C(AES_CORE_DATAPATH__abc_15863_new_n6805_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6806_));
OAI21X1 OAI21X1_1285 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4823_), .C(AES_CORE_DATAPATH__abc_15863_new_n6811_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6812_));
OAI21X1 OAI21X1_1286 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4858_), .C(AES_CORE_DATAPATH__abc_15863_new_n6818_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6819_));
OAI21X1 OAI21X1_1287 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4897_), .C(AES_CORE_DATAPATH__abc_15863_new_n6824_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6825_));
OAI21X1 OAI21X1_1288 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4932_), .C(AES_CORE_DATAPATH__abc_15863_new_n6831_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6832_));
OAI21X1 OAI21X1_1289 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n4971_), .C(AES_CORE_DATAPATH__abc_15863_new_n6837_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6838_));
OAI21X1 OAI21X1_129 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2744_));
OAI21X1 OAI21X1_1290 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5010_), .C(AES_CORE_DATAPATH__abc_15863_new_n6843_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6844_));
OAI21X1 OAI21X1_1291 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5049_), .C(AES_CORE_DATAPATH__abc_15863_new_n6849_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6850_));
OAI21X1 OAI21X1_1292 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5088_), .C(AES_CORE_DATAPATH__abc_15863_new_n6855_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6856_));
OAI21X1 OAI21X1_1293 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5127_), .C(AES_CORE_DATAPATH__abc_15863_new_n6861_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6862_));
OAI21X1 OAI21X1_1294 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5163_), .C(AES_CORE_DATAPATH__abc_15863_new_n6868_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6869_));
OAI21X1 OAI21X1_1295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5202_), .C(AES_CORE_DATAPATH__abc_15863_new_n6874_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6875_));
OAI21X1 OAI21X1_1296 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5241_), .C(AES_CORE_DATAPATH__abc_15863_new_n6880_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6881_));
OAI21X1 OAI21X1_1297 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5280_), .C(AES_CORE_DATAPATH__abc_15863_new_n6886_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6887_));
OAI21X1 OAI21X1_1298 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5319_), .C(AES_CORE_DATAPATH__abc_15863_new_n6892_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6893_));
OAI21X1 OAI21X1_1299 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5358_), .C(AES_CORE_DATAPATH__abc_15863_new_n6898_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6899_));
OAI21X1 OAI21X1_13 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT_state_13_), .C(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n151_));
OAI21X1 OAI21X1_130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2747_));
OAI21X1 OAI21X1_1300 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5397_), .C(AES_CORE_DATAPATH__abc_15863_new_n6904_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6905_));
OAI21X1 OAI21X1_1301 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5436_), .C(AES_CORE_DATAPATH__abc_15863_new_n6910_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6911_));
OAI21X1 OAI21X1_1302 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5472_), .C(AES_CORE_DATAPATH__abc_15863_new_n6917_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6918_));
OAI21X1 OAI21X1_1303 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5511_), .C(AES_CORE_DATAPATH__abc_15863_new_n6923_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6924_));
OAI21X1 OAI21X1_1304 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5550_), .C(AES_CORE_DATAPATH__abc_15863_new_n6929_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6930_));
OAI21X1 OAI21X1_1305 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5589_), .C(AES_CORE_DATAPATH__abc_15863_new_n6935_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6936_));
OAI21X1 OAI21X1_1306 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5628_), .C(AES_CORE_DATAPATH__abc_15863_new_n6941_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6942_));
OAI21X1 OAI21X1_1307 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5667_), .C(AES_CORE_DATAPATH__abc_15863_new_n6947_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6948_));
OAI21X1 OAI21X1_1308 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5706_), .C(AES_CORE_DATAPATH__abc_15863_new_n6953_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6954_));
OAI21X1 OAI21X1_1309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5742_), .C(AES_CORE_DATAPATH__abc_15863_new_n6960_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6961_));
OAI21X1 OAI21X1_131 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2754_), .B(AES_CORE_DATAPATH__abc_15863_new_n2751_), .C(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2756_));
OAI21X1 OAI21X1_1310 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5781_), .C(AES_CORE_DATAPATH__abc_15863_new_n6966_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6967_));
OAI21X1 OAI21X1_1311 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n5820_), .C(AES_CORE_DATAPATH__abc_15863_new_n6972_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6973_));
OAI21X1 OAI21X1_1312 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n6979_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6980_));
OAI21X1 OAI21X1_1313 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6979_), .B(AES_CORE_DATAPATH__abc_15863_new_n6988_), .C(AES_CORE_DATAPATH__abc_15863_new_n6985_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6989_));
OAI21X1 OAI21X1_1314 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2457_), .B(AES_CORE_DATAPATH__abc_15863_new_n2716_), .C(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_15863_new_n6990_));
OAI21X1 OAI21X1_1315 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(\iv_en[3] ), .C(AES_CORE_DATAPATH__abc_15863_new_n6990_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6991_));
OAI21X1 OAI21X1_1316 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6979_), .B(AES_CORE_DATAPATH__abc_15863_new_n6993_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6994_));
OAI21X1 OAI21X1_1317 ( .A(\bus_in[2] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6996_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6997_));
OAI21X1 OAI21X1_1318 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6979_), .B(AES_CORE_DATAPATH__abc_15863_new_n6995_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6999_));
OAI21X1 OAI21X1_1319 ( .A(\bus_in[3] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n7004_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7005_));
OAI21X1 OAI21X1_132 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2756_), .B(AES_CORE_DATAPATH__abc_15863_new_n2753_), .C(AES_CORE_DATAPATH__abc_15863_new_n2744_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__1_));
OAI21X1 OAI21X1_1320 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6979_), .B(AES_CORE_DATAPATH__abc_15863_new_n7003_), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7007_));
OAI21X1 OAI21X1_1321 ( .A(\bus_in[4] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n7010_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7011_));
OAI21X1 OAI21X1_1322 ( .A(\bus_in[5] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7017_));
OAI21X1 OAI21X1_1323 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6979_), .B(AES_CORE_DATAPATH__abc_15863_new_n7016_), .C(AES_CORE_DATAPATH__abc_15863_new_n7018_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7019_));
OAI21X1 OAI21X1_1324 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2514_), .B(AES_CORE_DATAPATH__abc_15863_new_n6978_), .C(AES_CORE_DATAPATH__abc_15863_new_n7019_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__5_));
OAI21X1 OAI21X1_1325 ( .A(\bus_in[6] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7021_));
OAI21X1 OAI21X1_1326 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6979_), .B(AES_CORE_DATAPATH__abc_15863_new_n7023_), .C(AES_CORE_DATAPATH__abc_15863_new_n7022_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7024_));
OAI21X1 OAI21X1_1327 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2520_), .B(AES_CORE_DATAPATH__abc_15863_new_n6978_), .C(AES_CORE_DATAPATH__abc_15863_new_n7024_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__6_));
OAI21X1 OAI21X1_1328 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6980_), .B(AES_CORE_DATAPATH__abc_15863_new_n7030_), .C(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7032_));
OAI21X1 OAI21X1_1329 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6977_), .B(AES_CORE_DATAPATH__abc_15863_new_n7031_), .C(AES_CORE_DATAPATH__abc_15863_new_n7032_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__7_));
OAI21X1 OAI21X1_133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2760_));
OAI21X1 OAI21X1_1330 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6980_), .B(AES_CORE_DATAPATH__abc_15863_new_n7035_), .C(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7037_));
OAI21X1 OAI21X1_1331 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6977_), .B(AES_CORE_DATAPATH__abc_15863_new_n7036_), .C(AES_CORE_DATAPATH__abc_15863_new_n7037_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__8_));
OAI21X1 OAI21X1_1332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6982_), .B(AES_CORE_DATAPATH__abc_15863_new_n7042_), .C(AES_CORE_DATAPATH__abc_15863_new_n7040_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7043_));
OAI21X1 OAI21X1_1333 ( .A(AES_CORE_DATAPATH_iv_3__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n7034_), .C(AES_CORE_DATAPATH__abc_15863_new_n7043_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7044_));
OAI21X1 OAI21X1_1334 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6982_), .B(AES_CORE_DATAPATH__abc_15863_new_n7049_), .C(AES_CORE_DATAPATH__abc_15863_new_n7047_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7050_));
OAI21X1 OAI21X1_1335 ( .A(AES_CORE_DATAPATH_iv_3__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n7042_), .C(AES_CORE_DATAPATH__abc_15863_new_n7050_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7051_));
OAI21X1 OAI21X1_1336 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6982_), .B(AES_CORE_DATAPATH__abc_15863_new_n7055_), .C(AES_CORE_DATAPATH__abc_15863_new_n7054_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7056_));
OAI21X1 OAI21X1_1337 ( .A(AES_CORE_DATAPATH_iv_3__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n7049_), .C(AES_CORE_DATAPATH__abc_15863_new_n7056_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7057_));
OAI21X1 OAI21X1_1338 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2560_), .B(AES_CORE_DATAPATH__abc_15863_new_n7048_), .C(AES_CORE_DATAPATH__abc_15863_new_n2568_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7061_));
OAI21X1 OAI21X1_1339 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4279_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7063_));
OAI21X1 OAI21X1_134 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2766_));
OAI21X1 OAI21X1_1340 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2574_), .B(AES_CORE_DATAPATH__abc_15863_new_n7060_), .C(AES_CORE_DATAPATH__abc_15863_new_n7066_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7067_));
OAI21X1 OAI21X1_1341 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4284_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7068_));
OAI21X1 OAI21X1_1342 ( .A(AES_CORE_DATAPATH_iv_3__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n7071_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7073_));
OAI21X1 OAI21X1_1343 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4289_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7075_));
OAI21X1 OAI21X1_1344 ( .A(AES_CORE_DATAPATH_iv_3__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n7072_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7079_));
OAI21X1 OAI21X1_1345 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4294_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7081_));
OAI21X1 OAI21X1_1346 ( .A(AES_CORE_DATAPATH_iv_3__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n7078_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7086_));
OAI21X1 OAI21X1_1347 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4299_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7088_));
OAI21X1 OAI21X1_1348 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2602_), .B(AES_CORE_DATAPATH__abc_15863_new_n7084_), .C(AES_CORE_DATAPATH__abc_15863_new_n7091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7092_));
OAI21X1 OAI21X1_1349 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4304_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7093_));
OAI21X1 OAI21X1_135 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2765_), .C(AES_CORE_DATAPATH__abc_15863_new_n2766_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__2_));
OAI21X1 OAI21X1_1350 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2602_), .B(AES_CORE_DATAPATH__abc_15863_new_n7084_), .C(AES_CORE_DATAPATH__abc_15863_new_n2610_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7096_));
OAI21X1 OAI21X1_1351 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4309_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7099_));
OAI21X1 OAI21X1_1352 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2618_), .B(AES_CORE_DATAPATH__abc_15863_new_n7097_), .C(AES_CORE_DATAPATH__abc_15863_new_n7102_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7103_));
OAI21X1 OAI21X1_1353 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4314_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7104_));
OAI21X1 OAI21X1_1354 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7116_), .B(AES_CORE_DATAPATH__abc_15863_new_n7118_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7119_));
OAI21X1 OAI21X1_1355 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4319_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7120_));
OAI21X1 OAI21X1_1356 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7124_), .B(AES_CORE_DATAPATH__abc_15863_new_n7125_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7126_));
OAI21X1 OAI21X1_1357 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4324_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7127_));
OAI21X1 OAI21X1_1358 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7132_), .B(AES_CORE_DATAPATH__abc_15863_new_n7133_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7134_));
OAI21X1 OAI21X1_1359 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4329_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7135_));
OAI21X1 OAI21X1_136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2772_));
OAI21X1 OAI21X1_1360 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7138_), .B(AES_CORE_DATAPATH__abc_15863_new_n7140_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7141_));
OAI21X1 OAI21X1_1361 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4334_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7142_));
OAI21X1 OAI21X1_1362 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7151_), .B(AES_CORE_DATAPATH__abc_15863_new_n7150_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7152_));
OAI21X1 OAI21X1_1363 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4339_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7153_));
OAI21X1 OAI21X1_1364 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7157_), .B(AES_CORE_DATAPATH__abc_15863_new_n7158_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7159_));
OAI21X1 OAI21X1_1365 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4344_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7160_));
OAI21X1 OAI21X1_1366 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7167_), .B(AES_CORE_DATAPATH__abc_15863_new_n7166_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7168_));
OAI21X1 OAI21X1_1367 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4349_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7169_));
OAI21X1 OAI21X1_1368 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7172_), .B(AES_CORE_DATAPATH__abc_15863_new_n7174_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7175_));
OAI21X1 OAI21X1_1369 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4354_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7176_));
OAI21X1 OAI21X1_137 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2776_));
OAI21X1 OAI21X1_1370 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7181_), .B(AES_CORE_DATAPATH__abc_15863_new_n7183_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7184_));
OAI21X1 OAI21X1_1371 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4359_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7185_));
OAI21X1 OAI21X1_1372 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7188_), .B(AES_CORE_DATAPATH__abc_15863_new_n7190_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7191_));
OAI21X1 OAI21X1_1373 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4364_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7192_));
OAI21X1 OAI21X1_1374 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7197_), .B(AES_CORE_DATAPATH__abc_15863_new_n7198_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7199_));
OAI21X1 OAI21X1_1375 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4369_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7200_));
OAI21X1 OAI21X1_1376 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7203_), .B(AES_CORE_DATAPATH__abc_15863_new_n7205_), .C(AES_CORE_DATAPATH__abc_15863_new_n6981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7206_));
OAI21X1 OAI21X1_1377 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4023_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n6978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7207_));
OAI21X1 OAI21X1_1378 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2481_), .C(AES_CORE_DATAPATH__abc_15863_new_n7210_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__0_));
OAI21X1 OAI21X1_1379 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2490_), .C(AES_CORE_DATAPATH__abc_15863_new_n7212_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__1_));
OAI21X1 OAI21X1_138 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2775_), .C(AES_CORE_DATAPATH__abc_15863_new_n2776_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__3_));
OAI21X1 OAI21X1_1380 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2504_), .C(AES_CORE_DATAPATH__abc_15863_new_n7216_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__3_));
OAI21X1 OAI21X1_1381 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2524_), .C(AES_CORE_DATAPATH__abc_15863_new_n7222_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__6_));
OAI21X1 OAI21X1_1382 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2532_), .C(AES_CORE_DATAPATH__abc_15863_new_n7224_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__7_));
OAI21X1 OAI21X1_1383 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2540_), .C(AES_CORE_DATAPATH__abc_15863_new_n7226_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__8_));
OAI21X1 OAI21X1_1384 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2548_), .C(AES_CORE_DATAPATH__abc_15863_new_n7228_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__9_));
OAI21X1 OAI21X1_1385 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2556_), .C(AES_CORE_DATAPATH__abc_15863_new_n7230_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__10_));
OAI21X1 OAI21X1_1386 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2564_), .C(AES_CORE_DATAPATH__abc_15863_new_n7232_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__11_));
OAI21X1 OAI21X1_1387 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2578_), .C(AES_CORE_DATAPATH__abc_15863_new_n7236_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__13_));
OAI21X1 OAI21X1_1388 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2592_), .C(AES_CORE_DATAPATH__abc_15863_new_n7240_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__15_));
OAI21X1 OAI21X1_1389 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2606_), .C(AES_CORE_DATAPATH__abc_15863_new_n7244_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__17_));
OAI21X1 OAI21X1_139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2782_));
OAI21X1 OAI21X1_1390 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2614_), .C(AES_CORE_DATAPATH__abc_15863_new_n7246_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__18_));
OAI21X1 OAI21X1_1391 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2622_), .C(AES_CORE_DATAPATH__abc_15863_new_n7248_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__19_));
OAI21X1 OAI21X1_1392 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2636_), .C(AES_CORE_DATAPATH__abc_15863_new_n7252_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__21_));
OAI21X1 OAI21X1_1393 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2650_), .C(AES_CORE_DATAPATH__abc_15863_new_n7256_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__23_));
OAI21X1 OAI21X1_1394 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2664_), .C(AES_CORE_DATAPATH__abc_15863_new_n7260_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__25_));
OAI21X1 OAI21X1_1395 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2672_), .C(AES_CORE_DATAPATH__abc_15863_new_n7262_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__26_));
OAI21X1 OAI21X1_1396 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2686_), .C(AES_CORE_DATAPATH__abc_15863_new_n7266_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__28_));
OAI21X1 OAI21X1_1397 ( .A(\iv_en[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2706_), .C(AES_CORE_DATAPATH__abc_15863_new_n7272_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__31_));
OAI21X1 OAI21X1_1398 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6280_), .C(AES_CORE_DATAPATH__abc_15863_new_n7275_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__0_));
OAI21X1 OAI21X1_1399 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6287_), .C(AES_CORE_DATAPATH__abc_15863_new_n7277_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__1_));
OAI21X1 OAI21X1_14 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n151_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n152_));
OAI21X1 OAI21X1_140 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2786_));
OAI21X1 OAI21X1_1400 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6294_), .C(AES_CORE_DATAPATH__abc_15863_new_n7279_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__2_));
OAI21X1 OAI21X1_1401 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6301_), .C(AES_CORE_DATAPATH__abc_15863_new_n7281_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__3_));
OAI21X1 OAI21X1_1402 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6308_), .C(AES_CORE_DATAPATH__abc_15863_new_n7283_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__4_));
OAI21X1 OAI21X1_1403 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6315_), .C(AES_CORE_DATAPATH__abc_15863_new_n7285_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__5_));
OAI21X1 OAI21X1_1404 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6322_), .C(AES_CORE_DATAPATH__abc_15863_new_n7287_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__6_));
OAI21X1 OAI21X1_1405 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6329_), .C(AES_CORE_DATAPATH__abc_15863_new_n7289_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__7_));
OAI21X1 OAI21X1_1406 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6336_), .C(AES_CORE_DATAPATH__abc_15863_new_n7291_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__8_));
OAI21X1 OAI21X1_1407 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6343_), .C(AES_CORE_DATAPATH__abc_15863_new_n7293_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__9_));
OAI21X1 OAI21X1_1408 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6350_), .C(AES_CORE_DATAPATH__abc_15863_new_n7295_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__10_));
OAI21X1 OAI21X1_1409 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6357_), .C(AES_CORE_DATAPATH__abc_15863_new_n7297_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__11_));
OAI21X1 OAI21X1_141 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2785_), .C(AES_CORE_DATAPATH__abc_15863_new_n2786_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__4_));
OAI21X1 OAI21X1_1410 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6364_), .C(AES_CORE_DATAPATH__abc_15863_new_n7299_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__12_));
OAI21X1 OAI21X1_1411 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6371_), .C(AES_CORE_DATAPATH__abc_15863_new_n7301_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__13_));
OAI21X1 OAI21X1_1412 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6378_), .C(AES_CORE_DATAPATH__abc_15863_new_n7303_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__14_));
OAI21X1 OAI21X1_1413 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6385_), .C(AES_CORE_DATAPATH__abc_15863_new_n7305_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__15_));
OAI21X1 OAI21X1_1414 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6392_), .C(AES_CORE_DATAPATH__abc_15863_new_n7307_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__16_));
OAI21X1 OAI21X1_1415 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6399_), .C(AES_CORE_DATAPATH__abc_15863_new_n7309_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__17_));
OAI21X1 OAI21X1_1416 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6406_), .C(AES_CORE_DATAPATH__abc_15863_new_n7311_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__18_));
OAI21X1 OAI21X1_1417 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6413_), .C(AES_CORE_DATAPATH__abc_15863_new_n7313_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__19_));
OAI21X1 OAI21X1_1418 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6420_), .C(AES_CORE_DATAPATH__abc_15863_new_n7315_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__20_));
OAI21X1 OAI21X1_1419 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6427_), .C(AES_CORE_DATAPATH__abc_15863_new_n7317_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__21_));
OAI21X1 OAI21X1_142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2790_));
OAI21X1 OAI21X1_1420 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6434_), .C(AES_CORE_DATAPATH__abc_15863_new_n7319_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__22_));
OAI21X1 OAI21X1_1421 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6441_), .C(AES_CORE_DATAPATH__abc_15863_new_n7321_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__23_));
OAI21X1 OAI21X1_1422 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6448_), .C(AES_CORE_DATAPATH__abc_15863_new_n7323_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__24_));
OAI21X1 OAI21X1_1423 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6455_), .C(AES_CORE_DATAPATH__abc_15863_new_n7325_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__25_));
OAI21X1 OAI21X1_1424 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6462_), .C(AES_CORE_DATAPATH__abc_15863_new_n7327_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__26_));
OAI21X1 OAI21X1_1425 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6469_), .C(AES_CORE_DATAPATH__abc_15863_new_n7329_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__27_));
OAI21X1 OAI21X1_1426 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6476_), .C(AES_CORE_DATAPATH__abc_15863_new_n7331_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__28_));
OAI21X1 OAI21X1_1427 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6483_), .C(AES_CORE_DATAPATH__abc_15863_new_n7333_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__29_));
OAI21X1 OAI21X1_1428 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6490_), .C(AES_CORE_DATAPATH__abc_15863_new_n7335_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__30_));
OAI21X1 OAI21X1_1429 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7274_), .B(AES_CORE_DATAPATH__abc_15863_new_n6497_), .C(AES_CORE_DATAPATH__abc_15863_new_n7337_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__31_));
OAI21X1 OAI21X1_143 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2796_));
OAI21X1 OAI21X1_1430 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6279_), .C(AES_CORE_DATAPATH__abc_15863_new_n7340_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7341_));
OAI21X1 OAI21X1_1431 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6286_), .C(AES_CORE_DATAPATH__abc_15863_new_n7345_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7346_));
OAI21X1 OAI21X1_1432 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6293_), .C(AES_CORE_DATAPATH__abc_15863_new_n7350_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7351_));
OAI21X1 OAI21X1_1433 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6300_), .C(AES_CORE_DATAPATH__abc_15863_new_n7355_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7356_));
OAI21X1 OAI21X1_1434 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6307_), .C(AES_CORE_DATAPATH__abc_15863_new_n7360_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7361_));
OAI21X1 OAI21X1_1435 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6314_), .C(AES_CORE_DATAPATH__abc_15863_new_n7365_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7366_));
OAI21X1 OAI21X1_1436 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6321_), .C(AES_CORE_DATAPATH__abc_15863_new_n7370_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7371_));
OAI21X1 OAI21X1_1437 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6328_), .C(AES_CORE_DATAPATH__abc_15863_new_n7375_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7376_));
OAI21X1 OAI21X1_1438 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6335_), .C(AES_CORE_DATAPATH__abc_15863_new_n7380_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7381_));
OAI21X1 OAI21X1_1439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6342_), .C(AES_CORE_DATAPATH__abc_15863_new_n7385_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7386_));
OAI21X1 OAI21X1_144 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2795_), .C(AES_CORE_DATAPATH__abc_15863_new_n2796_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__5_));
OAI21X1 OAI21X1_1440 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6349_), .C(AES_CORE_DATAPATH__abc_15863_new_n7390_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7391_));
OAI21X1 OAI21X1_1441 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6356_), .C(AES_CORE_DATAPATH__abc_15863_new_n7395_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7396_));
OAI21X1 OAI21X1_1442 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6363_), .C(AES_CORE_DATAPATH__abc_15863_new_n7400_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7401_));
OAI21X1 OAI21X1_1443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6370_), .C(AES_CORE_DATAPATH__abc_15863_new_n7405_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7406_));
OAI21X1 OAI21X1_1444 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6377_), .C(AES_CORE_DATAPATH__abc_15863_new_n7410_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7411_));
OAI21X1 OAI21X1_1445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6384_), .C(AES_CORE_DATAPATH__abc_15863_new_n7415_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7416_));
OAI21X1 OAI21X1_1446 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6391_), .C(AES_CORE_DATAPATH__abc_15863_new_n7420_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7421_));
OAI21X1 OAI21X1_1447 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6398_), .C(AES_CORE_DATAPATH__abc_15863_new_n7425_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7426_));
OAI21X1 OAI21X1_1448 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6405_), .C(AES_CORE_DATAPATH__abc_15863_new_n7430_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7431_));
OAI21X1 OAI21X1_1449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6412_), .C(AES_CORE_DATAPATH__abc_15863_new_n7435_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7436_));
OAI21X1 OAI21X1_145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2802_));
OAI21X1 OAI21X1_1450 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6419_), .C(AES_CORE_DATAPATH__abc_15863_new_n7440_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7441_));
OAI21X1 OAI21X1_1451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6426_), .C(AES_CORE_DATAPATH__abc_15863_new_n7445_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7446_));
OAI21X1 OAI21X1_1452 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6433_), .C(AES_CORE_DATAPATH__abc_15863_new_n7450_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7451_));
OAI21X1 OAI21X1_1453 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6440_), .C(AES_CORE_DATAPATH__abc_15863_new_n7455_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7456_));
OAI21X1 OAI21X1_1454 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6447_), .C(AES_CORE_DATAPATH__abc_15863_new_n7460_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7461_));
OAI21X1 OAI21X1_1455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6454_), .C(AES_CORE_DATAPATH__abc_15863_new_n7465_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7466_));
OAI21X1 OAI21X1_1456 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6461_), .C(AES_CORE_DATAPATH__abc_15863_new_n7470_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7471_));
OAI21X1 OAI21X1_1457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6468_), .C(AES_CORE_DATAPATH__abc_15863_new_n7475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7476_));
OAI21X1 OAI21X1_1458 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6475_), .C(AES_CORE_DATAPATH__abc_15863_new_n7480_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7481_));
OAI21X1 OAI21X1_1459 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6482_), .C(AES_CORE_DATAPATH__abc_15863_new_n7485_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7486_));
OAI21X1 OAI21X1_146 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2806_));
OAI21X1 OAI21X1_1460 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6489_), .C(AES_CORE_DATAPATH__abc_15863_new_n7490_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7491_));
OAI21X1 OAI21X1_1461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6496_), .C(AES_CORE_DATAPATH__abc_15863_new_n7495_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7496_));
OAI21X1 OAI21X1_1462 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2469_), .C(AES_CORE_DATAPATH__abc_15863_new_n7499_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__0_));
OAI21X1 OAI21X1_1463 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2521_), .C(AES_CORE_DATAPATH__abc_15863_new_n7511_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__6_));
OAI21X1 OAI21X1_1464 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2529_), .C(AES_CORE_DATAPATH__abc_15863_new_n7513_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__7_));
OAI21X1 OAI21X1_1465 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2537_), .C(AES_CORE_DATAPATH__abc_15863_new_n7515_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__8_));
OAI21X1 OAI21X1_1466 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2545_), .C(AES_CORE_DATAPATH__abc_15863_new_n7517_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__9_));
OAI21X1 OAI21X1_1467 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2553_), .C(AES_CORE_DATAPATH__abc_15863_new_n7519_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__10_));
OAI21X1 OAI21X1_1468 ( .A(\iv_en[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2561_), .C(AES_CORE_DATAPATH__abc_15863_new_n7521_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__11_));
OAI21X1 OAI21X1_1469 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6505_), .C(AES_CORE_DATAPATH__abc_15863_new_n7564_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__0_));
OAI21X1 OAI21X1_147 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2805_), .C(AES_CORE_DATAPATH__abc_15863_new_n2806_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__6_));
OAI21X1 OAI21X1_1470 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6518_), .C(AES_CORE_DATAPATH__abc_15863_new_n7569_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__2_));
OAI21X1 OAI21X1_1471 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6531_), .C(AES_CORE_DATAPATH__abc_15863_new_n7574_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__4_));
OAI21X1 OAI21X1_1472 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6538_), .C(AES_CORE_DATAPATH__abc_15863_new_n7576_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__5_));
OAI21X1 OAI21X1_1473 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6545_), .C(AES_CORE_DATAPATH__abc_15863_new_n7578_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__6_));
OAI21X1 OAI21X1_1474 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6558_), .C(AES_CORE_DATAPATH__abc_15863_new_n7583_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__8_));
OAI21X1 OAI21X1_1475 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6571_), .C(AES_CORE_DATAPATH__abc_15863_new_n7588_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__10_));
OAI21X1 OAI21X1_1476 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6584_), .C(AES_CORE_DATAPATH__abc_15863_new_n7593_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__12_));
OAI21X1 OAI21X1_1477 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6597_), .C(AES_CORE_DATAPATH__abc_15863_new_n7598_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__14_));
OAI21X1 OAI21X1_1478 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6610_), .C(AES_CORE_DATAPATH__abc_15863_new_n7603_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__16_));
OAI21X1 OAI21X1_1479 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6635_), .C(AES_CORE_DATAPATH__abc_15863_new_n7614_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__20_));
OAI21X1 OAI21X1_148 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2808_));
OAI21X1 OAI21X1_1480 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6648_), .C(AES_CORE_DATAPATH__abc_15863_new_n7619_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__22_));
OAI21X1 OAI21X1_1481 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6661_), .C(AES_CORE_DATAPATH__abc_15863_new_n7624_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__24_));
OAI21X1 OAI21X1_1482 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6680_), .C(AES_CORE_DATAPATH__abc_15863_new_n7632_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__27_));
OAI21X1 OAI21X1_1483 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6693_), .C(AES_CORE_DATAPATH__abc_15863_new_n7637_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__29_));
OAI21X1 OAI21X1_1484 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7563_), .B(AES_CORE_DATAPATH__abc_15863_new_n6700_), .C(AES_CORE_DATAPATH__abc_15863_new_n7639_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__30_));
OAI21X1 OAI21X1_1485 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6504_), .C(AES_CORE_DATAPATH__abc_15863_new_n7646_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7647_));
OAI21X1 OAI21X1_1486 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6510_), .C(AES_CORE_DATAPATH__abc_15863_new_n7651_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7652_));
OAI21X1 OAI21X1_1487 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6517_), .C(AES_CORE_DATAPATH__abc_15863_new_n7657_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7658_));
OAI21X1 OAI21X1_1488 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6523_), .C(AES_CORE_DATAPATH__abc_15863_new_n7662_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7663_));
OAI21X1 OAI21X1_1489 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6530_), .C(AES_CORE_DATAPATH__abc_15863_new_n7668_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7669_));
OAI21X1 OAI21X1_149 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2811_));
OAI21X1 OAI21X1_1490 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6537_), .C(AES_CORE_DATAPATH__abc_15863_new_n7674_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7675_));
OAI21X1 OAI21X1_1491 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6544_), .C(AES_CORE_DATAPATH__abc_15863_new_n7680_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7681_));
OAI21X1 OAI21X1_1492 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6550_), .C(AES_CORE_DATAPATH__abc_15863_new_n7685_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7686_));
OAI21X1 OAI21X1_1493 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6557_), .C(AES_CORE_DATAPATH__abc_15863_new_n7691_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7692_));
OAI21X1 OAI21X1_1494 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6563_), .C(AES_CORE_DATAPATH__abc_15863_new_n7696_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7697_));
OAI21X1 OAI21X1_1495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6570_), .C(AES_CORE_DATAPATH__abc_15863_new_n7702_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7703_));
OAI21X1 OAI21X1_1496 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6576_), .C(AES_CORE_DATAPATH__abc_15863_new_n7707_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7708_));
OAI21X1 OAI21X1_1497 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6583_), .C(AES_CORE_DATAPATH__abc_15863_new_n7713_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7714_));
OAI21X1 OAI21X1_1498 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6589_), .C(AES_CORE_DATAPATH__abc_15863_new_n7718_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7719_));
OAI21X1 OAI21X1_1499 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6596_), .C(AES_CORE_DATAPATH__abc_15863_new_n7724_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7725_));
OAI21X1 OAI21X1_15 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n154_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n155_));
OAI21X1 OAI21X1_150 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2818_), .B(AES_CORE_DATAPATH__abc_15863_new_n2815_), .C(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2819_));
OAI21X1 OAI21X1_1500 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6602_), .C(AES_CORE_DATAPATH__abc_15863_new_n7729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7730_));
OAI21X1 OAI21X1_1501 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6609_), .C(AES_CORE_DATAPATH__abc_15863_new_n7735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7736_));
OAI21X1 OAI21X1_1502 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6615_), .C(AES_CORE_DATAPATH__abc_15863_new_n7740_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7741_));
OAI21X1 OAI21X1_1503 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6621_), .C(AES_CORE_DATAPATH__abc_15863_new_n7745_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7746_));
OAI21X1 OAI21X1_1504 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6627_), .C(AES_CORE_DATAPATH__abc_15863_new_n7750_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7751_));
OAI21X1 OAI21X1_1505 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6634_), .C(AES_CORE_DATAPATH__abc_15863_new_n7756_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7757_));
OAI21X1 OAI21X1_1506 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6640_), .C(AES_CORE_DATAPATH__abc_15863_new_n7761_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7762_));
OAI21X1 OAI21X1_1507 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6647_), .C(AES_CORE_DATAPATH__abc_15863_new_n7767_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7768_));
OAI21X1 OAI21X1_1508 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6653_), .C(AES_CORE_DATAPATH__abc_15863_new_n7772_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7773_));
OAI21X1 OAI21X1_1509 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6660_), .C(AES_CORE_DATAPATH__abc_15863_new_n7778_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7779_));
OAI21X1 OAI21X1_151 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2819_), .B(AES_CORE_DATAPATH__abc_15863_new_n2817_), .C(AES_CORE_DATAPATH__abc_15863_new_n2808_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__7_));
OAI21X1 OAI21X1_1510 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6666_), .C(AES_CORE_DATAPATH__abc_15863_new_n7783_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7784_));
OAI21X1 OAI21X1_1511 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6672_), .C(AES_CORE_DATAPATH__abc_15863_new_n7788_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7789_));
OAI21X1 OAI21X1_1512 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6679_), .C(AES_CORE_DATAPATH__abc_15863_new_n7794_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7795_));
OAI21X1 OAI21X1_1513 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6685_), .C(AES_CORE_DATAPATH__abc_15863_new_n7799_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7800_));
OAI21X1 OAI21X1_1514 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6692_), .C(AES_CORE_DATAPATH__abc_15863_new_n7805_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7806_));
OAI21X1 OAI21X1_1515 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6699_), .C(AES_CORE_DATAPATH__abc_15863_new_n7811_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7812_));
OAI21X1 OAI21X1_1516 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6705_), .C(AES_CORE_DATAPATH__abc_15863_new_n7816_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7817_));
OAI21X1 OAI21X1_1517 ( .A(\iv_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n7832_), .C(AES_CORE_DATAPATH__abc_15863_new_n7833_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__6_));
OAI21X1 OAI21X1_1518 ( .A(\iv_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n7835_), .C(AES_CORE_DATAPATH__abc_15863_new_n7836_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__7_));
OAI21X1 OAI21X1_1519 ( .A(\iv_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n7838_), .C(AES_CORE_DATAPATH__abc_15863_new_n7839_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__8_));
OAI21X1 OAI21X1_152 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2821_));
OAI21X1 OAI21X1_1520 ( .A(\iv_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n7841_), .C(AES_CORE_DATAPATH__abc_15863_new_n7842_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__9_));
OAI21X1 OAI21X1_1521 ( .A(\iv_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n7844_), .C(AES_CORE_DATAPATH__abc_15863_new_n7845_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__10_));
OAI21X1 OAI21X1_1522 ( .A(\iv_en[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n7847_), .C(AES_CORE_DATAPATH__abc_15863_new_n7848_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__11_));
OAI21X1 OAI21X1_1523 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6056_), .C(AES_CORE_DATAPATH__abc_15863_new_n7891_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__0_));
OAI21X1 OAI21X1_1524 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6063_), .C(AES_CORE_DATAPATH__abc_15863_new_n7893_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__1_));
OAI21X1 OAI21X1_1525 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6070_), .C(AES_CORE_DATAPATH__abc_15863_new_n7895_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__2_));
OAI21X1 OAI21X1_1526 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6077_), .C(AES_CORE_DATAPATH__abc_15863_new_n7897_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__3_));
OAI21X1 OAI21X1_1527 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6084_), .C(AES_CORE_DATAPATH__abc_15863_new_n7899_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__4_));
OAI21X1 OAI21X1_1528 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6091_), .C(AES_CORE_DATAPATH__abc_15863_new_n7901_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__5_));
OAI21X1 OAI21X1_1529 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6098_), .C(AES_CORE_DATAPATH__abc_15863_new_n7903_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__6_));
OAI21X1 OAI21X1_153 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2824_));
OAI21X1 OAI21X1_1530 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6105_), .C(AES_CORE_DATAPATH__abc_15863_new_n7905_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__7_));
OAI21X1 OAI21X1_1531 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6112_), .C(AES_CORE_DATAPATH__abc_15863_new_n7907_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__8_));
OAI21X1 OAI21X1_1532 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6119_), .C(AES_CORE_DATAPATH__abc_15863_new_n7909_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__9_));
OAI21X1 OAI21X1_1533 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6126_), .C(AES_CORE_DATAPATH__abc_15863_new_n7911_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__10_));
OAI21X1 OAI21X1_1534 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6133_), .C(AES_CORE_DATAPATH__abc_15863_new_n7913_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__11_));
OAI21X1 OAI21X1_1535 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6140_), .C(AES_CORE_DATAPATH__abc_15863_new_n7915_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__12_));
OAI21X1 OAI21X1_1536 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6147_), .C(AES_CORE_DATAPATH__abc_15863_new_n7917_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__13_));
OAI21X1 OAI21X1_1537 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6154_), .C(AES_CORE_DATAPATH__abc_15863_new_n7919_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__14_));
OAI21X1 OAI21X1_1538 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6161_), .C(AES_CORE_DATAPATH__abc_15863_new_n7921_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__15_));
OAI21X1 OAI21X1_1539 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6168_), .C(AES_CORE_DATAPATH__abc_15863_new_n7923_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__16_));
OAI21X1 OAI21X1_154 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2831_), .B(AES_CORE_DATAPATH__abc_15863_new_n2828_), .C(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2832_));
OAI21X1 OAI21X1_1540 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6175_), .C(AES_CORE_DATAPATH__abc_15863_new_n7925_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__17_));
OAI21X1 OAI21X1_1541 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6182_), .C(AES_CORE_DATAPATH__abc_15863_new_n7927_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__18_));
OAI21X1 OAI21X1_1542 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6189_), .C(AES_CORE_DATAPATH__abc_15863_new_n7929_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__19_));
OAI21X1 OAI21X1_1543 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6196_), .C(AES_CORE_DATAPATH__abc_15863_new_n7931_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__20_));
OAI21X1 OAI21X1_1544 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6203_), .C(AES_CORE_DATAPATH__abc_15863_new_n7933_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__21_));
OAI21X1 OAI21X1_1545 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6210_), .C(AES_CORE_DATAPATH__abc_15863_new_n7935_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__22_));
OAI21X1 OAI21X1_1546 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6217_), .C(AES_CORE_DATAPATH__abc_15863_new_n7937_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__23_));
OAI21X1 OAI21X1_1547 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6224_), .C(AES_CORE_DATAPATH__abc_15863_new_n7939_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__24_));
OAI21X1 OAI21X1_1548 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6231_), .C(AES_CORE_DATAPATH__abc_15863_new_n7941_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__25_));
OAI21X1 OAI21X1_1549 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6238_), .C(AES_CORE_DATAPATH__abc_15863_new_n7943_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__26_));
OAI21X1 OAI21X1_155 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2832_), .B(AES_CORE_DATAPATH__abc_15863_new_n2830_), .C(AES_CORE_DATAPATH__abc_15863_new_n2821_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__8_));
OAI21X1 OAI21X1_1550 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6245_), .C(AES_CORE_DATAPATH__abc_15863_new_n7945_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__27_));
OAI21X1 OAI21X1_1551 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6252_), .C(AES_CORE_DATAPATH__abc_15863_new_n7947_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__28_));
OAI21X1 OAI21X1_1552 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6259_), .C(AES_CORE_DATAPATH__abc_15863_new_n7949_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__29_));
OAI21X1 OAI21X1_1553 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6266_), .C(AES_CORE_DATAPATH__abc_15863_new_n7951_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__30_));
OAI21X1 OAI21X1_1554 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7890_), .B(AES_CORE_DATAPATH__abc_15863_new_n6273_), .C(AES_CORE_DATAPATH__abc_15863_new_n7953_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__31_));
OAI21X1 OAI21X1_1555 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6055_), .C(AES_CORE_DATAPATH__abc_15863_new_n7957_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7958_));
OAI21X1 OAI21X1_1556 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6062_), .C(AES_CORE_DATAPATH__abc_15863_new_n7963_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7964_));
OAI21X1 OAI21X1_1557 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6069_), .C(AES_CORE_DATAPATH__abc_15863_new_n7969_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7970_));
OAI21X1 OAI21X1_1558 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6076_), .C(AES_CORE_DATAPATH__abc_15863_new_n7975_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7976_));
OAI21X1 OAI21X1_1559 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6083_), .C(AES_CORE_DATAPATH__abc_15863_new_n7981_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7982_));
OAI21X1 OAI21X1_156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2836_));
OAI21X1 OAI21X1_1560 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6090_), .C(AES_CORE_DATAPATH__abc_15863_new_n7987_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7988_));
OAI21X1 OAI21X1_1561 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6097_), .C(AES_CORE_DATAPATH__abc_15863_new_n7993_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7994_));
OAI21X1 OAI21X1_1562 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6104_), .C(AES_CORE_DATAPATH__abc_15863_new_n7999_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8000_));
OAI21X1 OAI21X1_1563 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6111_), .C(AES_CORE_DATAPATH__abc_15863_new_n8005_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8006_));
OAI21X1 OAI21X1_1564 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6118_), .C(AES_CORE_DATAPATH__abc_15863_new_n8011_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8012_));
OAI21X1 OAI21X1_1565 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6125_), .C(AES_CORE_DATAPATH__abc_15863_new_n8017_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8018_));
OAI21X1 OAI21X1_1566 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6132_), .C(AES_CORE_DATAPATH__abc_15863_new_n8023_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8024_));
OAI21X1 OAI21X1_1567 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6139_), .C(AES_CORE_DATAPATH__abc_15863_new_n8029_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8030_));
OAI21X1 OAI21X1_1568 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6146_), .C(AES_CORE_DATAPATH__abc_15863_new_n8035_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8036_));
OAI21X1 OAI21X1_1569 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6153_), .C(AES_CORE_DATAPATH__abc_15863_new_n8041_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8042_));
OAI21X1 OAI21X1_157 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2842_));
OAI21X1 OAI21X1_1570 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6160_), .C(AES_CORE_DATAPATH__abc_15863_new_n8047_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8048_));
OAI21X1 OAI21X1_1571 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6167_), .C(AES_CORE_DATAPATH__abc_15863_new_n8053_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8054_));
OAI21X1 OAI21X1_1572 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6174_), .C(AES_CORE_DATAPATH__abc_15863_new_n8059_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8060_));
OAI21X1 OAI21X1_1573 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6181_), .C(AES_CORE_DATAPATH__abc_15863_new_n8065_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8066_));
OAI21X1 OAI21X1_1574 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6188_), .C(AES_CORE_DATAPATH__abc_15863_new_n8071_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8072_));
OAI21X1 OAI21X1_1575 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6195_), .C(AES_CORE_DATAPATH__abc_15863_new_n8077_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8078_));
OAI21X1 OAI21X1_1576 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6202_), .C(AES_CORE_DATAPATH__abc_15863_new_n8083_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8084_));
OAI21X1 OAI21X1_1577 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6209_), .C(AES_CORE_DATAPATH__abc_15863_new_n8089_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8090_));
OAI21X1 OAI21X1_1578 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6216_), .C(AES_CORE_DATAPATH__abc_15863_new_n8095_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8096_));
OAI21X1 OAI21X1_1579 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6223_), .C(AES_CORE_DATAPATH__abc_15863_new_n8101_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8102_));
OAI21X1 OAI21X1_158 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2841_), .C(AES_CORE_DATAPATH__abc_15863_new_n2842_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__9_));
OAI21X1 OAI21X1_1580 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6230_), .C(AES_CORE_DATAPATH__abc_15863_new_n8107_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8108_));
OAI21X1 OAI21X1_1581 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6237_), .C(AES_CORE_DATAPATH__abc_15863_new_n8113_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8114_));
OAI21X1 OAI21X1_1582 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6244_), .C(AES_CORE_DATAPATH__abc_15863_new_n8119_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8120_));
OAI21X1 OAI21X1_1583 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6251_), .C(AES_CORE_DATAPATH__abc_15863_new_n8125_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8126_));
OAI21X1 OAI21X1_1584 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6258_), .C(AES_CORE_DATAPATH__abc_15863_new_n8131_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8132_));
OAI21X1 OAI21X1_1585 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6265_), .C(AES_CORE_DATAPATH__abc_15863_new_n8137_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8138_));
OAI21X1 OAI21X1_1586 ( .A(AES_CORE_DATAPATH__abc_15863_new_n6778_), .B(AES_CORE_DATAPATH__abc_15863_new_n6272_), .C(AES_CORE_DATAPATH__abc_15863_new_n8143_), .Y(AES_CORE_DATAPATH__abc_15863_new_n8144_));
OAI21X1 OAI21X1_1587 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n8147_), .C(AES_CORE_DATAPATH__abc_15863_new_n8148_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__0_));
OAI21X1 OAI21X1_1588 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n8150_), .C(AES_CORE_DATAPATH__abc_15863_new_n8151_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__1_));
OAI21X1 OAI21X1_1589 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n8153_), .C(AES_CORE_DATAPATH__abc_15863_new_n8154_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__2_));
OAI21X1 OAI21X1_159 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2844_));
OAI21X1 OAI21X1_1590 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2458_), .B(AES_CORE_DATAPATH__abc_15863_new_n8156_), .C(AES_CORE_DATAPATH__abc_15863_new_n8157_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__3_));
OAI21X1 OAI21X1_1591 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH__abc_15863_new_n4030_), .C(AES_CORE_DATAPATH__abc_15863_new_n8159_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__0_));
OAI21X1 OAI21X1_1592 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH__abc_15863_new_n8161_), .C(AES_CORE_DATAPATH__abc_15863_new_n8162_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__1_));
OAI21X1 OAI21X1_1593 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH__abc_15863_new_n8164_), .C(AES_CORE_DATAPATH__abc_15863_new_n8165_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__2_));
OAI21X1 OAI21X1_1594 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_DATAPATH__abc_15863_new_n8167_), .C(AES_CORE_DATAPATH__abc_15863_new_n8168_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__3_));
OAI21X1 OAI21X1_1595 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n8147_), .C(AES_CORE_DATAPATH__abc_15863_new_n8170_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__0_));
OAI21X1 OAI21X1_1596 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n8150_), .C(AES_CORE_DATAPATH__abc_15863_new_n8172_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__1_));
OAI21X1 OAI21X1_1597 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n8153_), .C(AES_CORE_DATAPATH__abc_15863_new_n8174_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__2_));
OAI21X1 OAI21X1_1598 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n8156_), .C(AES_CORE_DATAPATH__abc_15863_new_n8176_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__3_));
OAI21X1 OAI21X1_1599 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n416_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n415_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n413_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n417_));
OAI21X1 OAI21X1_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n126_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n171_));
OAI21X1 OAI21X1_160 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2847_));
OAI21X1 OAI21X1_1600 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n418_));
OAI21X1 OAI21X1_1601 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n423_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n426_));
OAI21X1 OAI21X1_1602 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n422_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n426_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n419_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n427_));
OAI21X1 OAI21X1_1603 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n405_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n445_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n446_));
OAI21X1 OAI21X1_1604 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n444_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n446_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n438_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n447_));
OAI21X1 OAI21X1_1605 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n426_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n465_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n463_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n466_));
OAI21X1 OAI21X1_1606 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n482_));
OAI21X1 OAI21X1_1607 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n482_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n483_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n484_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n485_));
OAI21X1 OAI21X1_1608 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n439_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n441_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n477_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n497_));
OAI21X1 OAI21X1_1609 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n483_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n446_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n496_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n499_));
OAI21X1 OAI21X1_161 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2852_), .C(AES_CORE_DATAPATH__abc_15863_new_n2844_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__10_));
OAI21X1 OAI21X1_1610 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n509_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n510_));
OAI21X1 OAI21X1_1611 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n511_));
OAI21X1 OAI21X1_1612 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n465_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n510_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n514_));
OAI21X1 OAI21X1_1613 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n519_));
OAI21X1 OAI21X1_1614 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n509_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n520_));
OAI21X1 OAI21X1_1615 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n444_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n520_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n523_));
OAI21X1 OAI21X1_1616 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n528_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n529_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_));
OAI21X1 OAI21X1_1617 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n532_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n533_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_));
OAI21X1 OAI21X1_1618 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n536_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n537_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_));
OAI21X1 OAI21X1_1619 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n540_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n541_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_));
OAI21X1 OAI21X1_162 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2856_));
OAI21X1 OAI21X1_1620 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n544_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n545_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_));
OAI21X1 OAI21X1_1621 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n548_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n549_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_));
OAI21X1 OAI21X1_1622 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n552_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n553_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_));
OAI21X1 OAI21X1_1623 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n556_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n557_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_));
OAI21X1 OAI21X1_1624 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n560_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n561_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_));
OAI21X1 OAI21X1_1625 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n564_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n565_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_));
OAI21X1 OAI21X1_1626 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n568_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n569_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_));
OAI21X1 OAI21X1_1627 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n572_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n573_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_));
OAI21X1 OAI21X1_1628 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n576_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n577_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_));
OAI21X1 OAI21X1_1629 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n580_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n581_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_));
OAI21X1 OAI21X1_163 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2862_));
OAI21X1 OAI21X1_1630 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n584_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n585_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_));
OAI21X1 OAI21X1_1631 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n588_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n589_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_));
OAI21X1 OAI21X1_1632 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n592_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n593_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_));
OAI21X1 OAI21X1_1633 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n596_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n597_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_));
OAI21X1 OAI21X1_1634 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n600_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n601_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_));
OAI21X1 OAI21X1_1635 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n604_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n605_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_));
OAI21X1 OAI21X1_1636 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n608_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n609_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_));
OAI21X1 OAI21X1_1637 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n612_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n613_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_));
OAI21X1 OAI21X1_1638 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n616_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n617_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_));
OAI21X1 OAI21X1_1639 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n620_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n621_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_));
OAI21X1 OAI21X1_164 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2861_), .C(AES_CORE_DATAPATH__abc_15863_new_n2862_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__11_));
OAI21X1 OAI21X1_1640 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n624_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n625_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_));
OAI21X1 OAI21X1_1641 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n628_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n629_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_));
OAI21X1 OAI21X1_1642 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n632_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n633_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_));
OAI21X1 OAI21X1_1643 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n636_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n637_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_));
OAI21X1 OAI21X1_1644 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n640_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n641_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_));
OAI21X1 OAI21X1_1645 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n644_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n645_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_));
OAI21X1 OAI21X1_1646 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n648_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n649_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_));
OAI21X1 OAI21X1_1647 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n403_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n652_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n653_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_));
OAI21X1 OAI21X1_1648 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n108_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n109_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n110_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n111_));
OAI21X1 OAI21X1_1649 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n115_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n117_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n119_));
OAI21X1 OAI21X1_165 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2866_));
OAI21X1 OAI21X1_1650 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n152_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n151_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n153_));
OAI21X1 OAI21X1_1651 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n152_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n151_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n138_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n155_));
OAI21X1 OAI21X1_1652 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n176_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n182_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n138_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n183_));
OAI21X1 OAI21X1_1653 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n184_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n185_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n186_));
OAI21X1 OAI21X1_1654 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n176_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n182_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n191_));
OAI21X1 OAI21X1_1655 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n184_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n185_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n138_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n192_));
OAI21X1 OAI21X1_1656 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n218_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n220_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n221_));
OAI21X1 OAI21X1_1657 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n132_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n137_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n240_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n241_));
OAI21X1 OAI21X1_1658 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n149_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n148_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n242_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n243_));
OAI21X1 OAI21X1_1659 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n213_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n215_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n245_));
OAI21X1 OAI21X1_166 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2872_));
OAI21X1 OAI21X1_1660 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n218_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n220_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n144_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n246_));
OAI21X1 OAI21X1_1661 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n258_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n260_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n261_));
OAI21X1 OAI21X1_1662 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n263_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n265_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n259_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n266_));
OAI21X1 OAI21X1_1663 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n132_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n137_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n242_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n278_));
OAI21X1 OAI21X1_1664 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n149_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n148_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n240_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n279_));
OAI21X1 OAI21X1_1665 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n258_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n260_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n112_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n282_));
OAI21X1 OAI21X1_1666 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n176_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n182_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n299_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n300_));
OAI21X1 OAI21X1_1667 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n184_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n185_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n301_));
OAI21X1 OAI21X1_1668 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n251_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n252_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n303_));
OAI21X1 OAI21X1_1669 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n139_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n140_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n304_));
OAI21X1 OAI21X1_167 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2871_), .C(AES_CORE_DATAPATH__abc_15863_new_n2872_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__12_));
OAI21X1 OAI21X1_1670 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n139_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n140_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n306_));
OAI21X1 OAI21X1_1671 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n251_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n252_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n307_));
OAI21X1 OAI21X1_1672 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n305_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n308_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n244_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n309_));
OAI21X1 OAI21X1_1673 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n305_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n308_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n280_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n314_));
OAI21X1 OAI21X1_1674 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n318_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n319_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n320_));
OAI21X1 OAI21X1_1675 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n366_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n365_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n363_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n367_));
OAI21X1 OAI21X1_1676 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n386_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n387_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n388_));
OAI21X1 OAI21X1_1677 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n318_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n319_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n472_));
OAI21X1 OAI21X1_1678 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n366_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n365_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n492_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n493_));
OAI21X1 OAI21X1_1679 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n386_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n387_), .C(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n505_));
OAI21X1 OAI21X1_168 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2878_));
OAI21X1 OAI21X1_1680 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n102_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n107_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_));
OAI21X1 OAI21X1_1681 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n121_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n123_));
OAI21X1 OAI21X1_1682 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n76_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n123_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_));
OAI21X1 OAI21X1_1683 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n97_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n125_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_));
OAI21X1 OAI21X1_1684 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n127_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n133_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_));
OAI21X1 OAI21X1_1685 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n141_));
OAI21X1 OAI21X1_1686 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n146_));
OAI21X1 OAI21X1_1687 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n150_));
OAI21X1 OAI21X1_1688 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n171_));
OAI21X1 OAI21X1_1689 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n170_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_));
OAI21X1 OAI21X1_169 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2882_));
OAI21X1 OAI21X1_1690 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n187_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n188_));
OAI21X1 OAI21X1_1691 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n178_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n200_));
OAI21X1 OAI21X1_1692 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_));
OAI21X1 OAI21X1_1693 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n209_));
OAI21X1 OAI21X1_1694 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n213_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n221_));
OAI21X1 OAI21X1_1695 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n260_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n261_));
OAI21X1 OAI21X1_1696 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n275_));
OAI21X1 OAI21X1_1697 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n280_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n285_));
OAI21X1 OAI21X1_1698 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n290_));
OAI21X1 OAI21X1_1699 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n291_));
OAI21X1 OAI21X1_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n180_), .Y(AES_CORE_CONTROL_UNIT_col_en_3_));
OAI21X1 OAI21X1_170 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2881_), .C(AES_CORE_DATAPATH__abc_15863_new_n2882_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__13_));
OAI21X1 OAI21X1_1700 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n304_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n305_));
OAI21X1 OAI21X1_1701 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n316_));
OAI21X1 OAI21X1_1702 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n331_));
OAI21X1 OAI21X1_1703 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n332_));
OAI21X1 OAI21X1_1704 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n371_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n372_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n376_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n377_));
OAI21X1 OAI21X1_1705 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n387_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n117_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n388_));
OAI21X1 OAI21X1_1706 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n92_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n390_));
OAI21X1 OAI21X1_1707 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n396_));
OAI21X1 OAI21X1_1708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n399_));
OAI21X1 OAI21X1_1709 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n400_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n401_));
OAI21X1 OAI21X1_171 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2886_));
OAI21X1 OAI21X1_1710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n393_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n399_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n402_));
OAI21X1 OAI21X1_1711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n404_));
OAI21X1 OAI21X1_1712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n405_));
OAI21X1 OAI21X1_1713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n415_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n403_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n417_));
OAI21X1 OAI21X1_1714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n419_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n421_));
OAI21X1 OAI21X1_1715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n430_));
OAI21X1 OAI21X1_1716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n432_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n106_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n433_));
OAI21X1 OAI21X1_1717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n434_));
OAI21X1 OAI21X1_1718 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n78_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n440_));
OAI21X1 OAI21X1_1719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n446_));
OAI21X1 OAI21X1_172 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2892_));
OAI21X1 OAI21X1_1720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n448_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n439_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n449_));
OAI21X1 OAI21X1_1721 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n81_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n458_));
OAI21X1 OAI21X1_1722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n459_));
OAI21X1 OAI21X1_1723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n461_));
OAI21X1 OAI21X1_1724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n462_));
OAI21X1 OAI21X1_1725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n432_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n477_));
OAI21X1 OAI21X1_1726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n478_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n479_));
OAI21X1 OAI21X1_1727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n484_));
OAI21X1 OAI21X1_1728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n496_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n339_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n497_));
OAI21X1 OAI21X1_1729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n102_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n107_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_));
OAI21X1 OAI21X1_173 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2891_), .C(AES_CORE_DATAPATH__abc_15863_new_n2892_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__14_));
OAI21X1 OAI21X1_1730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n121_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n123_));
OAI21X1 OAI21X1_1731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n76_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n123_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_));
OAI21X1 OAI21X1_1732 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n97_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n125_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_));
OAI21X1 OAI21X1_1733 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n127_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n133_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_));
OAI21X1 OAI21X1_1734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n141_));
OAI21X1 OAI21X1_1735 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n146_));
OAI21X1 OAI21X1_1736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n150_));
OAI21X1 OAI21X1_1737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n171_));
OAI21X1 OAI21X1_1738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n170_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_));
OAI21X1 OAI21X1_1739 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n187_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n188_));
OAI21X1 OAI21X1_174 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2898_));
OAI21X1 OAI21X1_1740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n178_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n200_));
OAI21X1 OAI21X1_1741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_));
OAI21X1 OAI21X1_1742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n209_));
OAI21X1 OAI21X1_1743 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n213_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n221_));
OAI21X1 OAI21X1_1744 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n260_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n261_));
OAI21X1 OAI21X1_1745 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n275_));
OAI21X1 OAI21X1_1746 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n280_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n285_));
OAI21X1 OAI21X1_1747 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n290_));
OAI21X1 OAI21X1_1748 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n291_));
OAI21X1 OAI21X1_1749 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n304_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n305_));
OAI21X1 OAI21X1_175 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2902_));
OAI21X1 OAI21X1_1750 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n316_));
OAI21X1 OAI21X1_1751 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n331_));
OAI21X1 OAI21X1_1752 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n332_));
OAI21X1 OAI21X1_1753 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n371_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n372_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n376_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n377_));
OAI21X1 OAI21X1_1754 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n387_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n117_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n388_));
OAI21X1 OAI21X1_1755 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n92_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n390_));
OAI21X1 OAI21X1_1756 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n396_));
OAI21X1 OAI21X1_1757 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n399_));
OAI21X1 OAI21X1_1758 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n400_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n401_));
OAI21X1 OAI21X1_1759 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n393_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n399_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n402_));
OAI21X1 OAI21X1_176 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2901_), .C(AES_CORE_DATAPATH__abc_15863_new_n2902_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__15_));
OAI21X1 OAI21X1_1760 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n404_));
OAI21X1 OAI21X1_1761 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n405_));
OAI21X1 OAI21X1_1762 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n415_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n403_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n417_));
OAI21X1 OAI21X1_1763 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n419_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n421_));
OAI21X1 OAI21X1_1764 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n430_));
OAI21X1 OAI21X1_1765 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n432_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n106_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n433_));
OAI21X1 OAI21X1_1766 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n434_));
OAI21X1 OAI21X1_1767 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n78_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n440_));
OAI21X1 OAI21X1_1768 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n446_));
OAI21X1 OAI21X1_1769 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n448_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n439_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n449_));
OAI21X1 OAI21X1_177 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2904_));
OAI21X1 OAI21X1_1770 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n81_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n458_));
OAI21X1 OAI21X1_1771 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n459_));
OAI21X1 OAI21X1_1772 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n461_));
OAI21X1 OAI21X1_1773 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n462_));
OAI21X1 OAI21X1_1774 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n432_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n477_));
OAI21X1 OAI21X1_1775 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n478_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n479_));
OAI21X1 OAI21X1_1776 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n484_));
OAI21X1 OAI21X1_1777 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n496_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n339_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n497_));
OAI21X1 OAI21X1_1778 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n102_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n107_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_));
OAI21X1 OAI21X1_1779 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n121_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n123_));
OAI21X1 OAI21X1_178 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2909_));
OAI21X1 OAI21X1_1780 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n76_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n123_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_));
OAI21X1 OAI21X1_1781 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n97_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n125_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_));
OAI21X1 OAI21X1_1782 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n127_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n133_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_));
OAI21X1 OAI21X1_1783 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n141_));
OAI21X1 OAI21X1_1784 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n146_));
OAI21X1 OAI21X1_1785 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n150_));
OAI21X1 OAI21X1_1786 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n171_));
OAI21X1 OAI21X1_1787 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n170_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_));
OAI21X1 OAI21X1_1788 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n187_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n188_));
OAI21X1 OAI21X1_1789 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n178_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n200_));
OAI21X1 OAI21X1_179 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2912_), .C(AES_CORE_DATAPATH__abc_15863_new_n2904_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__16_));
OAI21X1 OAI21X1_1790 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_));
OAI21X1 OAI21X1_1791 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n209_));
OAI21X1 OAI21X1_1792 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n213_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n221_));
OAI21X1 OAI21X1_1793 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n260_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n261_));
OAI21X1 OAI21X1_1794 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n275_));
OAI21X1 OAI21X1_1795 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n280_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n285_));
OAI21X1 OAI21X1_1796 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n290_));
OAI21X1 OAI21X1_1797 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n291_));
OAI21X1 OAI21X1_1798 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n304_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n305_));
OAI21X1 OAI21X1_1799 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n316_));
OAI21X1 OAI21X1_18 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n168_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n161_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n185_));
OAI21X1 OAI21X1_180 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2918_));
OAI21X1 OAI21X1_1800 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n331_));
OAI21X1 OAI21X1_1801 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n332_));
OAI21X1 OAI21X1_1802 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n371_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n372_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n376_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n377_));
OAI21X1 OAI21X1_1803 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n387_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n117_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n388_));
OAI21X1 OAI21X1_1804 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n92_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n390_));
OAI21X1 OAI21X1_1805 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n396_));
OAI21X1 OAI21X1_1806 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n399_));
OAI21X1 OAI21X1_1807 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n400_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n401_));
OAI21X1 OAI21X1_1808 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n393_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n399_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n402_));
OAI21X1 OAI21X1_1809 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n404_));
OAI21X1 OAI21X1_181 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2922_));
OAI21X1 OAI21X1_1810 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n405_));
OAI21X1 OAI21X1_1811 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n415_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n403_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n417_));
OAI21X1 OAI21X1_1812 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n419_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n421_));
OAI21X1 OAI21X1_1813 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n430_));
OAI21X1 OAI21X1_1814 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n432_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n106_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n433_));
OAI21X1 OAI21X1_1815 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n434_));
OAI21X1 OAI21X1_1816 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n78_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n440_));
OAI21X1 OAI21X1_1817 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n446_));
OAI21X1 OAI21X1_1818 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n448_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n439_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n449_));
OAI21X1 OAI21X1_1819 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n81_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n458_));
OAI21X1 OAI21X1_182 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2921_), .C(AES_CORE_DATAPATH__abc_15863_new_n2922_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__17_));
OAI21X1 OAI21X1_1820 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n459_));
OAI21X1 OAI21X1_1821 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n461_));
OAI21X1 OAI21X1_1822 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n462_));
OAI21X1 OAI21X1_1823 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n432_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n477_));
OAI21X1 OAI21X1_1824 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n478_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n479_));
OAI21X1 OAI21X1_1825 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n484_));
OAI21X1 OAI21X1_1826 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n496_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n339_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n497_));
OAI21X1 OAI21X1_1827 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n102_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n107_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_));
OAI21X1 OAI21X1_1828 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n121_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n123_));
OAI21X1 OAI21X1_1829 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n76_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n123_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_));
OAI21X1 OAI21X1_183 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2928_));
OAI21X1 OAI21X1_1830 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n97_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n125_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_));
OAI21X1 OAI21X1_1831 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n127_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n133_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_));
OAI21X1 OAI21X1_1832 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n141_));
OAI21X1 OAI21X1_1833 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n146_));
OAI21X1 OAI21X1_1834 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n136_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n150_));
OAI21X1 OAI21X1_1835 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n135_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n140_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n171_));
OAI21X1 OAI21X1_1836 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n170_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_));
OAI21X1 OAI21X1_1837 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n187_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n188_));
OAI21X1 OAI21X1_1838 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n178_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n200_));
OAI21X1 OAI21X1_1839 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_));
OAI21X1 OAI21X1_184 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2932_));
OAI21X1 OAI21X1_1840 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n209_));
OAI21X1 OAI21X1_1841 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n213_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n221_));
OAI21X1 OAI21X1_1842 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n214_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n260_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n261_));
OAI21X1 OAI21X1_1843 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n275_));
OAI21X1 OAI21X1_1844 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n280_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n285_));
OAI21X1 OAI21X1_1845 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n278_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n290_));
OAI21X1 OAI21X1_1846 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n286_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n291_));
OAI21X1 OAI21X1_1847 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n304_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n305_));
OAI21X1 OAI21X1_1848 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n270_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n271_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n316_));
OAI21X1 OAI21X1_1849 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n206_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n331_));
OAI21X1 OAI21X1_185 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2931_), .C(AES_CORE_DATAPATH__abc_15863_new_n2932_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__18_));
OAI21X1 OAI21X1_1850 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n332_));
OAI21X1 OAI21X1_1851 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n371_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n372_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n376_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n377_));
OAI21X1 OAI21X1_1852 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n387_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n117_), .C(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n388_));
OAI21X1 OAI21X1_1853 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n92_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n390_));
OAI21X1 OAI21X1_1854 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n396_));
OAI21X1 OAI21X1_1855 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n398_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n399_));
OAI21X1 OAI21X1_1856 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n400_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n401_));
OAI21X1 OAI21X1_1857 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n393_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n399_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n402_));
OAI21X1 OAI21X1_1858 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n404_));
OAI21X1 OAI21X1_1859 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n405_));
OAI21X1 OAI21X1_186 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2938_));
OAI21X1 OAI21X1_1860 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n415_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n403_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n417_));
OAI21X1 OAI21X1_1861 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n419_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n402_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n421_));
OAI21X1 OAI21X1_1862 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n430_));
OAI21X1 OAI21X1_1863 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n432_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n106_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n433_));
OAI21X1 OAI21X1_1864 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n434_));
OAI21X1 OAI21X1_1865 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n78_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n440_));
OAI21X1 OAI21X1_1866 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n385_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n446_));
OAI21X1 OAI21X1_1867 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n448_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n439_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n449_));
OAI21X1 OAI21X1_1868 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n81_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n428_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n458_));
OAI21X1 OAI21X1_1869 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n394_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n395_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n459_));
OAI21X1 OAI21X1_187 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2942_));
OAI21X1 OAI21X1_1870 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n95_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n407_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n461_));
OAI21X1 OAI21X1_1871 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n89_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n94_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n462_));
OAI21X1 OAI21X1_1872 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n432_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n477_));
OAI21X1 OAI21X1_1873 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n478_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n479_));
OAI21X1 OAI21X1_1874 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n425_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n456_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n484_));
OAI21X1 OAI21X1_1875 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n496_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n339_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n497_));
OAI21X1 OAI21X1_188 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2941_), .C(AES_CORE_DATAPATH__abc_15863_new_n2942_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__19_));
OAI21X1 OAI21X1_189 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2944_));
OAI21X1 OAI21X1_19 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n184_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n185_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n183_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n186_));
OAI21X1 OAI21X1_190 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2949_));
OAI21X1 OAI21X1_191 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2954_), .B(AES_CORE_DATAPATH__abc_15863_new_n2951_), .C(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2955_));
OAI21X1 OAI21X1_192 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2955_), .B(AES_CORE_DATAPATH__abc_15863_new_n2953_), .C(AES_CORE_DATAPATH__abc_15863_new_n2944_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__20_));
OAI21X1 OAI21X1_193 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2961_));
OAI21X1 OAI21X1_194 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2965_));
OAI21X1 OAI21X1_195 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2964_), .C(AES_CORE_DATAPATH__abc_15863_new_n2965_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__21_));
OAI21X1 OAI21X1_196 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2971_));
OAI21X1 OAI21X1_197 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2975_));
OAI21X1 OAI21X1_198 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n2974_), .C(AES_CORE_DATAPATH__abc_15863_new_n2975_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__22_));
OAI21X1 OAI21X1_199 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2977_));
OAI21X1 OAI21X1_2 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .C(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n88_));
OAI21X1 OAI21X1_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n123_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n187_));
OAI21X1 OAI21X1_200 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2982_));
OAI21X1 OAI21X1_201 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2987_), .B(AES_CORE_DATAPATH__abc_15863_new_n2984_), .C(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2988_));
OAI21X1 OAI21X1_202 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2988_), .B(AES_CORE_DATAPATH__abc_15863_new_n2986_), .C(AES_CORE_DATAPATH__abc_15863_new_n2977_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__23_));
OAI21X1 OAI21X1_203 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2990_));
OAI21X1 OAI21X1_204 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2993_));
OAI21X1 OAI21X1_205 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3000_), .B(AES_CORE_DATAPATH__abc_15863_new_n2997_), .C(AES_CORE_DATAPATH__abc_15863_new_n2755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3001_));
OAI21X1 OAI21X1_206 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3001_), .B(AES_CORE_DATAPATH__abc_15863_new_n2999_), .C(AES_CORE_DATAPATH__abc_15863_new_n2990_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__24_));
OAI21X1 OAI21X1_207 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3005_));
OAI21X1 OAI21X1_208 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3011_));
OAI21X1 OAI21X1_209 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3010_), .C(AES_CORE_DATAPATH__abc_15863_new_n3011_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__25_));
OAI21X1 OAI21X1_21 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n124_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n196_), .Y(AES_CORE_CONTROL_UNIT_key_sel));
OAI21X1 OAI21X1_210 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3015_));
OAI21X1 OAI21X1_211 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3021_));
OAI21X1 OAI21X1_212 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3020_), .C(AES_CORE_DATAPATH__abc_15863_new_n3021_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__26_));
OAI21X1 OAI21X1_213 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3025_));
OAI21X1 OAI21X1_214 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3031_));
OAI21X1 OAI21X1_215 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3030_), .C(AES_CORE_DATAPATH__abc_15863_new_n3031_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__27_));
OAI21X1 OAI21X1_216 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3033_));
OAI21X1 OAI21X1_217 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3036_));
OAI21X1 OAI21X1_218 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3041_), .C(AES_CORE_DATAPATH__abc_15863_new_n3033_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__28_));
OAI21X1 OAI21X1_219 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3043_));
OAI21X1 OAI21X1_22 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n199_), .Y(AES_CORE_CONTROL_UNIT_key_en_1_));
OAI21X1 OAI21X1_220 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3046_));
OAI21X1 OAI21X1_221 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3051_), .C(AES_CORE_DATAPATH__abc_15863_new_n3043_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__29_));
OAI21X1 OAI21X1_222 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3053_));
OAI21X1 OAI21X1_223 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3056_));
OAI21X1 OAI21X1_224 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3061_), .C(AES_CORE_DATAPATH__abc_15863_new_n3053_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__30_));
OAI21X1 OAI21X1_225 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH__abc_15863_new_n2735_), .C(AES_CORE_DATAPATH__abc_15863_new_n2737_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3067_));
OAI21X1 OAI21X1_226 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3071_));
OAI21X1 OAI21X1_227 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2710_), .B(AES_CORE_DATAPATH__abc_15863_new_n3070_), .C(AES_CORE_DATAPATH__abc_15863_new_n3071_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__31_));
OAI21X1 OAI21X1_228 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n3074_), .C(AES_CORE_DATAPATH__abc_15863_new_n3075_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3076_));
OAI21X1 OAI21X1_229 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n3077_), .C(AES_CORE_DATAPATH__abc_15863_new_n3078_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3079_));
OAI21X1 OAI21X1_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n108_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n201_));
OAI21X1 OAI21X1_230 ( .A(AES_CORE_DATAPATH_col_sel_host_1_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_1_), .C(AES_CORE_DATAPATH__abc_15863_new_n3083_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3084_));
OAI21X1 OAI21X1_231 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3081_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3090_));
OAI21X1 OAI21X1_232 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3096_), .B(AES_CORE_DATAPATH__abc_15863_new_n3090_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3097_));
OAI21X1 OAI21X1_233 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3107_), .B(AES_CORE_DATAPATH_last_round_pp2), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3109_));
OAI21X1 OAI21X1_234 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3112_), .C(AES_CORE_DATAPATH__abc_15863_new_n3113_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_));
OAI21X1 OAI21X1_235 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3122_), .B(AES_CORE_DATAPATH__abc_15863_new_n3118_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3124_));
OAI21X1 OAI21X1_236 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3131_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3132_));
OAI21X1 OAI21X1_237 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3135_), .C(AES_CORE_DATAPATH__abc_15863_new_n3136_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_));
OAI21X1 OAI21X1_238 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3138_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3139_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3140_));
OAI21X1 OAI21X1_239 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3144_), .B(AES_CORE_DATAPATH__abc_15863_new_n3140_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3146_));
OAI21X1 OAI21X1_24 ( .A(AES_CORE_CONTROL_UNIT_state_1_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n201_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_));
OAI21X1 OAI21X1_240 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3153_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3154_));
OAI21X1 OAI21X1_241 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3157_), .C(AES_CORE_DATAPATH__abc_15863_new_n3158_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_));
OAI21X1 OAI21X1_242 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3166_), .B(AES_CORE_DATAPATH__abc_15863_new_n3162_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3169_));
OAI21X1 OAI21X1_243 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3176_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3177_));
OAI21X1 OAI21X1_244 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3180_), .C(AES_CORE_DATAPATH__abc_15863_new_n3181_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_));
OAI21X1 OAI21X1_245 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3183_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3184_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3185_));
OAI21X1 OAI21X1_246 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3189_), .B(AES_CORE_DATAPATH__abc_15863_new_n3185_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3191_));
OAI21X1 OAI21X1_247 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3198_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3199_));
OAI21X1 OAI21X1_248 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3202_), .C(AES_CORE_DATAPATH__abc_15863_new_n3203_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_));
OAI21X1 OAI21X1_249 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3205_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3206_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3207_));
OAI21X1 OAI21X1_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n119_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n204_), .Y(AES_CORE_CONTROL_UNIT_key_en_3_));
OAI21X1 OAI21X1_250 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3211_), .B(AES_CORE_DATAPATH__abc_15863_new_n3207_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3213_));
OAI21X1 OAI21X1_251 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3220_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3221_));
OAI21X1 OAI21X1_252 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3224_), .C(AES_CORE_DATAPATH__abc_15863_new_n3225_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_));
OAI21X1 OAI21X1_253 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3227_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3228_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3229_));
OAI21X1 OAI21X1_254 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3233_), .B(AES_CORE_DATAPATH__abc_15863_new_n3229_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3235_));
OAI21X1 OAI21X1_255 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3242_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3243_));
OAI21X1 OAI21X1_256 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3246_), .C(AES_CORE_DATAPATH__abc_15863_new_n3247_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_));
OAI21X1 OAI21X1_257 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3255_), .B(AES_CORE_DATAPATH__abc_15863_new_n3251_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3257_));
OAI21X1 OAI21X1_258 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3264_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3265_));
OAI21X1 OAI21X1_259 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3268_), .C(AES_CORE_DATAPATH__abc_15863_new_n3269_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_));
OAI21X1 OAI21X1_26 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2479_));
OAI21X1 OAI21X1_260 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3271_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3272_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3273_));
OAI21X1 OAI21X1_261 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3277_), .B(AES_CORE_DATAPATH__abc_15863_new_n3273_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3279_));
OAI21X1 OAI21X1_262 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3286_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3287_));
OAI21X1 OAI21X1_263 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3290_), .C(AES_CORE_DATAPATH__abc_15863_new_n3291_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_));
OAI21X1 OAI21X1_264 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3299_), .B(AES_CORE_DATAPATH__abc_15863_new_n3295_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3301_));
OAI21X1 OAI21X1_265 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3308_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3309_));
OAI21X1 OAI21X1_266 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3312_), .C(AES_CORE_DATAPATH__abc_15863_new_n3313_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_));
OAI21X1 OAI21X1_267 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3315_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3316_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3317_));
OAI21X1 OAI21X1_268 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3321_), .B(AES_CORE_DATAPATH__abc_15863_new_n3317_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3323_));
OAI21X1 OAI21X1_269 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3330_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3331_));
OAI21X1 OAI21X1_27 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2480_), .C(AES_CORE_DATAPATH__abc_15863_new_n2483_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2484_));
OAI21X1 OAI21X1_270 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3334_), .C(AES_CORE_DATAPATH__abc_15863_new_n3335_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_));
OAI21X1 OAI21X1_271 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3343_), .B(AES_CORE_DATAPATH__abc_15863_new_n3339_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3345_));
OAI21X1 OAI21X1_272 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3352_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3353_));
OAI21X1 OAI21X1_273 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3356_), .C(AES_CORE_DATAPATH__abc_15863_new_n3357_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_));
OAI21X1 OAI21X1_274 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3359_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3360_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3361_));
OAI21X1 OAI21X1_275 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3365_), .B(AES_CORE_DATAPATH__abc_15863_new_n3361_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3367_));
OAI21X1 OAI21X1_276 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3374_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3375_));
OAI21X1 OAI21X1_277 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3378_), .C(AES_CORE_DATAPATH__abc_15863_new_n3379_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_));
OAI21X1 OAI21X1_278 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3387_), .B(AES_CORE_DATAPATH__abc_15863_new_n3383_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3389_));
OAI21X1 OAI21X1_279 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3396_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3397_));
OAI21X1 OAI21X1_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2457_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2484_), .Y(\iv_out[0] ));
OAI21X1 OAI21X1_280 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3400_), .C(AES_CORE_DATAPATH__abc_15863_new_n3401_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_));
OAI21X1 OAI21X1_281 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3403_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3404_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3405_));
OAI21X1 OAI21X1_282 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3409_), .B(AES_CORE_DATAPATH__abc_15863_new_n3405_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3411_));
OAI21X1 OAI21X1_283 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3418_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3419_));
OAI21X1 OAI21X1_284 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3422_), .C(AES_CORE_DATAPATH__abc_15863_new_n3423_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_));
OAI21X1 OAI21X1_285 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3431_), .B(AES_CORE_DATAPATH__abc_15863_new_n3427_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3433_));
OAI21X1 OAI21X1_286 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3440_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3441_));
OAI21X1 OAI21X1_287 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3444_), .C(AES_CORE_DATAPATH__abc_15863_new_n3445_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_));
OAI21X1 OAI21X1_288 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3447_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3448_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3449_));
OAI21X1 OAI21X1_289 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3453_), .B(AES_CORE_DATAPATH__abc_15863_new_n3449_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3455_));
OAI21X1 OAI21X1_29 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2487_));
OAI21X1 OAI21X1_290 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3462_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3463_));
OAI21X1 OAI21X1_291 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3466_), .C(AES_CORE_DATAPATH__abc_15863_new_n3467_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_));
OAI21X1 OAI21X1_292 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3475_), .B(AES_CORE_DATAPATH__abc_15863_new_n3471_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3477_));
OAI21X1 OAI21X1_293 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3484_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3485_));
OAI21X1 OAI21X1_294 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3488_), .C(AES_CORE_DATAPATH__abc_15863_new_n3489_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_));
OAI21X1 OAI21X1_295 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3497_), .B(AES_CORE_DATAPATH__abc_15863_new_n3493_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3499_));
OAI21X1 OAI21X1_296 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3506_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3507_));
OAI21X1 OAI21X1_297 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3510_), .C(AES_CORE_DATAPATH__abc_15863_new_n3511_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_));
OAI21X1 OAI21X1_298 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3519_), .B(AES_CORE_DATAPATH__abc_15863_new_n3515_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3521_));
OAI21X1 OAI21X1_299 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3528_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3529_));
OAI21X1 OAI21X1_3 ( .A(\aes_mode[0] ), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_), .C(\op_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_));
OAI21X1 OAI21X1_30 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2487_), .C(AES_CORE_DATAPATH__abc_15863_new_n2488_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2489_));
OAI21X1 OAI21X1_300 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3532_), .C(AES_CORE_DATAPATH__abc_15863_new_n3533_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_));
OAI21X1 OAI21X1_301 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3535_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3536_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3537_));
OAI21X1 OAI21X1_302 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3541_), .B(AES_CORE_DATAPATH__abc_15863_new_n3537_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3543_));
OAI21X1 OAI21X1_303 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3550_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3551_));
OAI21X1 OAI21X1_304 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3554_), .C(AES_CORE_DATAPATH__abc_15863_new_n3555_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_));
OAI21X1 OAI21X1_305 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3563_), .B(AES_CORE_DATAPATH__abc_15863_new_n3559_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3565_));
OAI21X1 OAI21X1_306 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3572_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3573_));
OAI21X1 OAI21X1_307 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3576_), .C(AES_CORE_DATAPATH__abc_15863_new_n3577_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_));
OAI21X1 OAI21X1_308 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3579_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3580_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3581_));
OAI21X1 OAI21X1_309 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3585_), .B(AES_CORE_DATAPATH__abc_15863_new_n3581_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3587_));
OAI21X1 OAI21X1_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2486_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2492_), .Y(\iv_out[1] ));
OAI21X1 OAI21X1_310 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3594_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3595_));
OAI21X1 OAI21X1_311 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3598_), .C(AES_CORE_DATAPATH__abc_15863_new_n3599_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_));
OAI21X1 OAI21X1_312 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3607_), .B(AES_CORE_DATAPATH__abc_15863_new_n3603_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3609_));
OAI21X1 OAI21X1_313 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3616_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3617_));
OAI21X1 OAI21X1_314 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3620_), .C(AES_CORE_DATAPATH__abc_15863_new_n3621_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_));
OAI21X1 OAI21X1_315 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3623_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3624_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3625_));
OAI21X1 OAI21X1_316 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3629_), .B(AES_CORE_DATAPATH__abc_15863_new_n3625_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3631_));
OAI21X1 OAI21X1_317 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3638_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3639_));
OAI21X1 OAI21X1_318 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3642_), .C(AES_CORE_DATAPATH__abc_15863_new_n3643_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_));
OAI21X1 OAI21X1_319 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3651_), .B(AES_CORE_DATAPATH__abc_15863_new_n3647_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3653_));
OAI21X1 OAI21X1_32 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2495_));
OAI21X1 OAI21X1_320 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3660_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3661_));
OAI21X1 OAI21X1_321 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3664_), .C(AES_CORE_DATAPATH__abc_15863_new_n3665_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_));
OAI21X1 OAI21X1_322 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3673_), .B(AES_CORE_DATAPATH__abc_15863_new_n3669_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3675_));
OAI21X1 OAI21X1_323 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3682_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3683_));
OAI21X1 OAI21X1_324 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3686_), .C(AES_CORE_DATAPATH__abc_15863_new_n3687_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_));
OAI21X1 OAI21X1_325 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3689_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3690_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3691_));
OAI21X1 OAI21X1_326 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3695_), .B(AES_CORE_DATAPATH__abc_15863_new_n3691_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3697_));
OAI21X1 OAI21X1_327 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3704_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3705_));
OAI21X1 OAI21X1_328 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3708_), .C(AES_CORE_DATAPATH__abc_15863_new_n3709_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_));
OAI21X1 OAI21X1_329 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3717_), .B(AES_CORE_DATAPATH__abc_15863_new_n3713_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3719_));
OAI21X1 OAI21X1_33 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2495_), .C(AES_CORE_DATAPATH__abc_15863_new_n2496_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2497_));
OAI21X1 OAI21X1_330 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3726_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3727_));
OAI21X1 OAI21X1_331 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3730_), .C(AES_CORE_DATAPATH__abc_15863_new_n3731_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_));
OAI21X1 OAI21X1_332 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3733_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3734_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3735_));
OAI21X1 OAI21X1_333 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3739_), .B(AES_CORE_DATAPATH__abc_15863_new_n3735_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3741_));
OAI21X1 OAI21X1_334 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3748_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3749_));
OAI21X1 OAI21X1_335 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3752_), .C(AES_CORE_DATAPATH__abc_15863_new_n3753_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_));
OAI21X1 OAI21X1_336 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3755_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3756_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3757_));
OAI21X1 OAI21X1_337 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3761_), .B(AES_CORE_DATAPATH__abc_15863_new_n3757_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3763_));
OAI21X1 OAI21X1_338 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3770_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3771_));
OAI21X1 OAI21X1_339 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3774_), .C(AES_CORE_DATAPATH__abc_15863_new_n3775_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_));
OAI21X1 OAI21X1_34 ( .A(AES_CORE_DATAPATH_iv_2__2_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2497_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2498_));
OAI21X1 OAI21X1_340 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3783_), .B(AES_CORE_DATAPATH__abc_15863_new_n3779_), .C(AES_CORE_DATAPATH__abc_15863_new_n3080_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3785_));
OAI21X1 OAI21X1_341 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH__abc_15863_new_n3792_), .C(AES_CORE_DATAPATH__abc_15863_new_n3108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3793_));
OAI21X1 OAI21X1_342 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2715_), .B(AES_CORE_DATAPATH__abc_15863_new_n3796_), .C(AES_CORE_DATAPATH__abc_15863_new_n3797_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_));
OAI21X1 OAI21X1_343 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3112_), .C(AES_CORE_DATAPATH__abc_15863_new_n3799_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_));
OAI21X1 OAI21X1_344 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3135_), .C(AES_CORE_DATAPATH__abc_15863_new_n3801_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_));
OAI21X1 OAI21X1_345 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3157_), .C(AES_CORE_DATAPATH__abc_15863_new_n3803_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_));
OAI21X1 OAI21X1_346 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3180_), .C(AES_CORE_DATAPATH__abc_15863_new_n3805_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_));
OAI21X1 OAI21X1_347 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3202_), .C(AES_CORE_DATAPATH__abc_15863_new_n3807_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_));
OAI21X1 OAI21X1_348 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3224_), .C(AES_CORE_DATAPATH__abc_15863_new_n3809_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_));
OAI21X1 OAI21X1_349 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3246_), .C(AES_CORE_DATAPATH__abc_15863_new_n3811_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_));
OAI21X1 OAI21X1_35 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2501_));
OAI21X1 OAI21X1_350 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3268_), .C(AES_CORE_DATAPATH__abc_15863_new_n3813_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_));
OAI21X1 OAI21X1_351 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3290_), .C(AES_CORE_DATAPATH__abc_15863_new_n3815_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_));
OAI21X1 OAI21X1_352 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3312_), .C(AES_CORE_DATAPATH__abc_15863_new_n3817_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_));
OAI21X1 OAI21X1_353 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3334_), .C(AES_CORE_DATAPATH__abc_15863_new_n3819_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_));
OAI21X1 OAI21X1_354 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3356_), .C(AES_CORE_DATAPATH__abc_15863_new_n3821_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_));
OAI21X1 OAI21X1_355 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3378_), .C(AES_CORE_DATAPATH__abc_15863_new_n3823_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_));
OAI21X1 OAI21X1_356 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3400_), .C(AES_CORE_DATAPATH__abc_15863_new_n3825_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_));
OAI21X1 OAI21X1_357 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3422_), .C(AES_CORE_DATAPATH__abc_15863_new_n3827_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_));
OAI21X1 OAI21X1_358 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3444_), .C(AES_CORE_DATAPATH__abc_15863_new_n3829_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_));
OAI21X1 OAI21X1_359 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3466_), .C(AES_CORE_DATAPATH__abc_15863_new_n3831_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_));
OAI21X1 OAI21X1_36 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2501_), .C(AES_CORE_DATAPATH__abc_15863_new_n2502_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2503_));
OAI21X1 OAI21X1_360 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3488_), .C(AES_CORE_DATAPATH__abc_15863_new_n3833_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_));
OAI21X1 OAI21X1_361 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3510_), .C(AES_CORE_DATAPATH__abc_15863_new_n3835_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_));
OAI21X1 OAI21X1_362 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3532_), .C(AES_CORE_DATAPATH__abc_15863_new_n3837_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_));
OAI21X1 OAI21X1_363 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3554_), .C(AES_CORE_DATAPATH__abc_15863_new_n3839_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_));
OAI21X1 OAI21X1_364 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3576_), .C(AES_CORE_DATAPATH__abc_15863_new_n3841_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_));
OAI21X1 OAI21X1_365 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3598_), .C(AES_CORE_DATAPATH__abc_15863_new_n3843_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_));
OAI21X1 OAI21X1_366 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3620_), .C(AES_CORE_DATAPATH__abc_15863_new_n3845_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_));
OAI21X1 OAI21X1_367 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3642_), .C(AES_CORE_DATAPATH__abc_15863_new_n3847_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_));
OAI21X1 OAI21X1_368 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3664_), .C(AES_CORE_DATAPATH__abc_15863_new_n3849_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_));
OAI21X1 OAI21X1_369 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3686_), .C(AES_CORE_DATAPATH__abc_15863_new_n3851_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_));
OAI21X1 OAI21X1_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2500_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2506_), .Y(\iv_out[3] ));
OAI21X1 OAI21X1_370 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3708_), .C(AES_CORE_DATAPATH__abc_15863_new_n3853_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_));
OAI21X1 OAI21X1_371 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3730_), .C(AES_CORE_DATAPATH__abc_15863_new_n3855_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_));
OAI21X1 OAI21X1_372 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3752_), .C(AES_CORE_DATAPATH__abc_15863_new_n3857_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_));
OAI21X1 OAI21X1_373 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3774_), .C(AES_CORE_DATAPATH__abc_15863_new_n3859_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_));
OAI21X1 OAI21X1_374 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH__abc_15863_new_n3796_), .C(AES_CORE_DATAPATH__abc_15863_new_n3861_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_));
OAI21X1 OAI21X1_375 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3869_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3870_));
OAI21X1 OAI21X1_376 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3870_), .C(AES_CORE_DATAPATH__abc_15863_new_n3871_), .Y(AES_CORE_DATAPATH__0key_1__31_0__0_));
OAI21X1 OAI21X1_377 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3874_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3875_));
OAI21X1 OAI21X1_378 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3875_), .C(AES_CORE_DATAPATH__abc_15863_new_n3876_), .Y(AES_CORE_DATAPATH__0key_1__31_0__1_));
OAI21X1 OAI21X1_379 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3879_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3880_));
OAI21X1 OAI21X1_38 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2509_));
OAI21X1 OAI21X1_380 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3880_), .C(AES_CORE_DATAPATH__abc_15863_new_n3881_), .Y(AES_CORE_DATAPATH__0key_1__31_0__2_));
OAI21X1 OAI21X1_381 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3884_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3885_));
OAI21X1 OAI21X1_382 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3885_), .C(AES_CORE_DATAPATH__abc_15863_new_n3886_), .Y(AES_CORE_DATAPATH__0key_1__31_0__3_));
OAI21X1 OAI21X1_383 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3889_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3890_));
OAI21X1 OAI21X1_384 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3890_), .C(AES_CORE_DATAPATH__abc_15863_new_n3891_), .Y(AES_CORE_DATAPATH__0key_1__31_0__4_));
OAI21X1 OAI21X1_385 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3894_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3895_));
OAI21X1 OAI21X1_386 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3895_), .C(AES_CORE_DATAPATH__abc_15863_new_n3896_), .Y(AES_CORE_DATAPATH__0key_1__31_0__5_));
OAI21X1 OAI21X1_387 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3899_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3900_));
OAI21X1 OAI21X1_388 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3900_), .C(AES_CORE_DATAPATH__abc_15863_new_n3901_), .Y(AES_CORE_DATAPATH__0key_1__31_0__6_));
OAI21X1 OAI21X1_389 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3904_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3905_));
OAI21X1 OAI21X1_39 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2509_), .C(AES_CORE_DATAPATH__abc_15863_new_n2510_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2511_));
OAI21X1 OAI21X1_390 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3905_), .C(AES_CORE_DATAPATH__abc_15863_new_n3906_), .Y(AES_CORE_DATAPATH__0key_1__31_0__7_));
OAI21X1 OAI21X1_391 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3909_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3910_));
OAI21X1 OAI21X1_392 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3910_), .C(AES_CORE_DATAPATH__abc_15863_new_n3911_), .Y(AES_CORE_DATAPATH__0key_1__31_0__8_));
OAI21X1 OAI21X1_393 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3914_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3915_));
OAI21X1 OAI21X1_394 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3915_), .C(AES_CORE_DATAPATH__abc_15863_new_n3916_), .Y(AES_CORE_DATAPATH__0key_1__31_0__9_));
OAI21X1 OAI21X1_395 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3919_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3920_));
OAI21X1 OAI21X1_396 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3920_), .C(AES_CORE_DATAPATH__abc_15863_new_n3921_), .Y(AES_CORE_DATAPATH__0key_1__31_0__10_));
OAI21X1 OAI21X1_397 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3924_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3925_));
OAI21X1 OAI21X1_398 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3925_), .C(AES_CORE_DATAPATH__abc_15863_new_n3926_), .Y(AES_CORE_DATAPATH__0key_1__31_0__11_));
OAI21X1 OAI21X1_399 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3929_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3930_));
OAI21X1 OAI21X1_4 ( .A(\op_mode[1] ), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n95_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n96_));
OAI21X1 OAI21X1_40 ( .A(AES_CORE_DATAPATH_iv_2__4_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2511_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2512_));
OAI21X1 OAI21X1_400 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3930_), .C(AES_CORE_DATAPATH__abc_15863_new_n3931_), .Y(AES_CORE_DATAPATH__0key_1__31_0__12_));
OAI21X1 OAI21X1_401 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3934_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3935_));
OAI21X1 OAI21X1_402 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3935_), .C(AES_CORE_DATAPATH__abc_15863_new_n3936_), .Y(AES_CORE_DATAPATH__0key_1__31_0__13_));
OAI21X1 OAI21X1_403 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3939_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3940_));
OAI21X1 OAI21X1_404 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3940_), .C(AES_CORE_DATAPATH__abc_15863_new_n3941_), .Y(AES_CORE_DATAPATH__0key_1__31_0__14_));
OAI21X1 OAI21X1_405 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3944_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3945_));
OAI21X1 OAI21X1_406 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3945_), .C(AES_CORE_DATAPATH__abc_15863_new_n3946_), .Y(AES_CORE_DATAPATH__0key_1__31_0__15_));
OAI21X1 OAI21X1_407 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3949_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3950_));
OAI21X1 OAI21X1_408 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3950_), .C(AES_CORE_DATAPATH__abc_15863_new_n3951_), .Y(AES_CORE_DATAPATH__0key_1__31_0__16_));
OAI21X1 OAI21X1_409 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3954_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3955_));
OAI21X1 OAI21X1_41 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2515_));
OAI21X1 OAI21X1_410 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3955_), .C(AES_CORE_DATAPATH__abc_15863_new_n3956_), .Y(AES_CORE_DATAPATH__0key_1__31_0__17_));
OAI21X1 OAI21X1_411 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3959_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3960_));
OAI21X1 OAI21X1_412 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3960_), .C(AES_CORE_DATAPATH__abc_15863_new_n3961_), .Y(AES_CORE_DATAPATH__0key_1__31_0__18_));
OAI21X1 OAI21X1_413 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3964_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3965_));
OAI21X1 OAI21X1_414 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3965_), .C(AES_CORE_DATAPATH__abc_15863_new_n3966_), .Y(AES_CORE_DATAPATH__0key_1__31_0__19_));
OAI21X1 OAI21X1_415 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3969_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3970_));
OAI21X1 OAI21X1_416 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3970_), .C(AES_CORE_DATAPATH__abc_15863_new_n3971_), .Y(AES_CORE_DATAPATH__0key_1__31_0__20_));
OAI21X1 OAI21X1_417 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3974_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3975_));
OAI21X1 OAI21X1_418 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3975_), .C(AES_CORE_DATAPATH__abc_15863_new_n3976_), .Y(AES_CORE_DATAPATH__0key_1__31_0__21_));
OAI21X1 OAI21X1_419 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3979_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3980_));
OAI21X1 OAI21X1_42 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2515_), .C(AES_CORE_DATAPATH__abc_15863_new_n2516_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2517_));
OAI21X1 OAI21X1_420 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3980_), .C(AES_CORE_DATAPATH__abc_15863_new_n3981_), .Y(AES_CORE_DATAPATH__0key_1__31_0__22_));
OAI21X1 OAI21X1_421 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3984_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3985_));
OAI21X1 OAI21X1_422 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3985_), .C(AES_CORE_DATAPATH__abc_15863_new_n3986_), .Y(AES_CORE_DATAPATH__0key_1__31_0__23_));
OAI21X1 OAI21X1_423 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3989_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3990_));
OAI21X1 OAI21X1_424 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3990_), .C(AES_CORE_DATAPATH__abc_15863_new_n3991_), .Y(AES_CORE_DATAPATH__0key_1__31_0__24_));
OAI21X1 OAI21X1_425 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3994_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3995_));
OAI21X1 OAI21X1_426 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n3995_), .C(AES_CORE_DATAPATH__abc_15863_new_n3996_), .Y(AES_CORE_DATAPATH__0key_1__31_0__25_));
OAI21X1 OAI21X1_427 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n3999_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4000_));
OAI21X1 OAI21X1_428 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4000_), .C(AES_CORE_DATAPATH__abc_15863_new_n4001_), .Y(AES_CORE_DATAPATH__0key_1__31_0__26_));
OAI21X1 OAI21X1_429 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4004_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4005_));
OAI21X1 OAI21X1_43 ( .A(AES_CORE_DATAPATH_iv_2__5_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2517_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2518_));
OAI21X1 OAI21X1_430 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4005_), .C(AES_CORE_DATAPATH__abc_15863_new_n4006_), .Y(AES_CORE_DATAPATH__0key_1__31_0__27_));
OAI21X1 OAI21X1_431 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4009_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4010_));
OAI21X1 OAI21X1_432 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4010_), .C(AES_CORE_DATAPATH__abc_15863_new_n4011_), .Y(AES_CORE_DATAPATH__0key_1__31_0__28_));
OAI21X1 OAI21X1_433 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4014_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4015_));
OAI21X1 OAI21X1_434 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4015_), .C(AES_CORE_DATAPATH__abc_15863_new_n4016_), .Y(AES_CORE_DATAPATH__0key_1__31_0__29_));
OAI21X1 OAI21X1_435 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4019_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4020_));
OAI21X1 OAI21X1_436 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4020_), .C(AES_CORE_DATAPATH__abc_15863_new_n4021_), .Y(AES_CORE_DATAPATH__0key_1__31_0__30_));
OAI21X1 OAI21X1_437 ( .A(\key_en[1] ), .B(AES_CORE_DATAPATH_key_host_1__31_), .C(AES_CORE_DATAPATH__abc_15863_new_n4024_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4025_));
OAI21X1 OAI21X1_438 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4026_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4027_));
OAI21X1 OAI21X1_439 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4027_), .C(AES_CORE_DATAPATH__abc_15863_new_n4028_), .Y(AES_CORE_DATAPATH__0key_1__31_0__31_));
OAI21X1 OAI21X1_44 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2522_));
OAI21X1 OAI21X1_440 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2712_), .B(AES_CORE_DATAPATH__abc_15863_new_n4030_), .C(AES_CORE_DATAPATH__abc_15863_new_n4031_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4032_));
OAI21X1 OAI21X1_441 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4037_), .C(AES_CORE_DATAPATH__abc_15863_new_n4038_), .Y(AES_CORE_DATAPATH__0key_0__31_0__0_));
OAI21X1 OAI21X1_442 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4041_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4042_));
OAI21X1 OAI21X1_443 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4042_), .C(AES_CORE_DATAPATH__abc_15863_new_n4043_), .Y(AES_CORE_DATAPATH__0key_0__31_0__1_));
OAI21X1 OAI21X1_444 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4046_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4047_));
OAI21X1 OAI21X1_445 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4047_), .C(AES_CORE_DATAPATH__abc_15863_new_n4048_), .Y(AES_CORE_DATAPATH__0key_0__31_0__2_));
OAI21X1 OAI21X1_446 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4051_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4052_));
OAI21X1 OAI21X1_447 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4052_), .C(AES_CORE_DATAPATH__abc_15863_new_n4053_), .Y(AES_CORE_DATAPATH__0key_0__31_0__3_));
OAI21X1 OAI21X1_448 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4056_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4057_));
OAI21X1 OAI21X1_449 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4057_), .C(AES_CORE_DATAPATH__abc_15863_new_n4058_), .Y(AES_CORE_DATAPATH__0key_0__31_0__4_));
OAI21X1 OAI21X1_45 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2523_), .C(AES_CORE_DATAPATH__abc_15863_new_n2525_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2526_));
OAI21X1 OAI21X1_450 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4061_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4062_));
OAI21X1 OAI21X1_451 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4062_), .C(AES_CORE_DATAPATH__abc_15863_new_n4063_), .Y(AES_CORE_DATAPATH__0key_0__31_0__5_));
OAI21X1 OAI21X1_452 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4066_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4067_));
OAI21X1 OAI21X1_453 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4067_), .C(AES_CORE_DATAPATH__abc_15863_new_n4068_), .Y(AES_CORE_DATAPATH__0key_0__31_0__6_));
OAI21X1 OAI21X1_454 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4071_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4072_));
OAI21X1 OAI21X1_455 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4072_), .C(AES_CORE_DATAPATH__abc_15863_new_n4073_), .Y(AES_CORE_DATAPATH__0key_0__31_0__7_));
OAI21X1 OAI21X1_456 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4076_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4077_));
OAI21X1 OAI21X1_457 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4077_), .C(AES_CORE_DATAPATH__abc_15863_new_n4078_), .Y(AES_CORE_DATAPATH__0key_0__31_0__8_));
OAI21X1 OAI21X1_458 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4081_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4082_));
OAI21X1 OAI21X1_459 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4082_), .C(AES_CORE_DATAPATH__abc_15863_new_n4083_), .Y(AES_CORE_DATAPATH__0key_0__31_0__9_));
OAI21X1 OAI21X1_46 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2520_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2526_), .Y(\iv_out[6] ));
OAI21X1 OAI21X1_460 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4087_));
OAI21X1 OAI21X1_461 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4087_), .C(AES_CORE_DATAPATH__abc_15863_new_n4088_), .Y(AES_CORE_DATAPATH__0key_0__31_0__10_));
OAI21X1 OAI21X1_462 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4091_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4092_));
OAI21X1 OAI21X1_463 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4092_), .C(AES_CORE_DATAPATH__abc_15863_new_n4093_), .Y(AES_CORE_DATAPATH__0key_0__31_0__11_));
OAI21X1 OAI21X1_464 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4096_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4097_));
OAI21X1 OAI21X1_465 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4097_), .C(AES_CORE_DATAPATH__abc_15863_new_n4098_), .Y(AES_CORE_DATAPATH__0key_0__31_0__12_));
OAI21X1 OAI21X1_466 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4101_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4102_));
OAI21X1 OAI21X1_467 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4102_), .C(AES_CORE_DATAPATH__abc_15863_new_n4103_), .Y(AES_CORE_DATAPATH__0key_0__31_0__13_));
OAI21X1 OAI21X1_468 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4106_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4107_));
OAI21X1 OAI21X1_469 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4107_), .C(AES_CORE_DATAPATH__abc_15863_new_n4108_), .Y(AES_CORE_DATAPATH__0key_0__31_0__14_));
OAI21X1 OAI21X1_47 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2530_));
OAI21X1 OAI21X1_470 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4111_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4112_));
OAI21X1 OAI21X1_471 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4112_), .C(AES_CORE_DATAPATH__abc_15863_new_n4113_), .Y(AES_CORE_DATAPATH__0key_0__31_0__15_));
OAI21X1 OAI21X1_472 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4116_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4117_));
OAI21X1 OAI21X1_473 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4117_), .C(AES_CORE_DATAPATH__abc_15863_new_n4118_), .Y(AES_CORE_DATAPATH__0key_0__31_0__16_));
OAI21X1 OAI21X1_474 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4121_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4122_));
OAI21X1 OAI21X1_475 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4122_), .C(AES_CORE_DATAPATH__abc_15863_new_n4123_), .Y(AES_CORE_DATAPATH__0key_0__31_0__17_));
OAI21X1 OAI21X1_476 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4126_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4127_));
OAI21X1 OAI21X1_477 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4127_), .C(AES_CORE_DATAPATH__abc_15863_new_n4128_), .Y(AES_CORE_DATAPATH__0key_0__31_0__18_));
OAI21X1 OAI21X1_478 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4131_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4132_));
OAI21X1 OAI21X1_479 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4132_), .C(AES_CORE_DATAPATH__abc_15863_new_n4133_), .Y(AES_CORE_DATAPATH__0key_0__31_0__19_));
OAI21X1 OAI21X1_48 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2531_), .C(AES_CORE_DATAPATH__abc_15863_new_n2533_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2534_));
OAI21X1 OAI21X1_480 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4136_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4137_));
OAI21X1 OAI21X1_481 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4137_), .C(AES_CORE_DATAPATH__abc_15863_new_n4138_), .Y(AES_CORE_DATAPATH__0key_0__31_0__20_));
OAI21X1 OAI21X1_482 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4141_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4142_));
OAI21X1 OAI21X1_483 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4142_), .C(AES_CORE_DATAPATH__abc_15863_new_n4143_), .Y(AES_CORE_DATAPATH__0key_0__31_0__21_));
OAI21X1 OAI21X1_484 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4146_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4147_));
OAI21X1 OAI21X1_485 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4147_), .C(AES_CORE_DATAPATH__abc_15863_new_n4148_), .Y(AES_CORE_DATAPATH__0key_0__31_0__22_));
OAI21X1 OAI21X1_486 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4151_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4152_));
OAI21X1 OAI21X1_487 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4152_), .C(AES_CORE_DATAPATH__abc_15863_new_n4153_), .Y(AES_CORE_DATAPATH__0key_0__31_0__23_));
OAI21X1 OAI21X1_488 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4156_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4157_));
OAI21X1 OAI21X1_489 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4157_), .C(AES_CORE_DATAPATH__abc_15863_new_n4158_), .Y(AES_CORE_DATAPATH__0key_0__31_0__24_));
OAI21X1 OAI21X1_49 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2528_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2534_), .Y(\iv_out[7] ));
OAI21X1 OAI21X1_490 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4161_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4162_));
OAI21X1 OAI21X1_491 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4162_), .C(AES_CORE_DATAPATH__abc_15863_new_n4163_), .Y(AES_CORE_DATAPATH__0key_0__31_0__25_));
OAI21X1 OAI21X1_492 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4166_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4167_));
OAI21X1 OAI21X1_493 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4167_), .C(AES_CORE_DATAPATH__abc_15863_new_n4168_), .Y(AES_CORE_DATAPATH__0key_0__31_0__26_));
OAI21X1 OAI21X1_494 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4171_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4172_));
OAI21X1 OAI21X1_495 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4172_), .C(AES_CORE_DATAPATH__abc_15863_new_n4173_), .Y(AES_CORE_DATAPATH__0key_0__31_0__27_));
OAI21X1 OAI21X1_496 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4176_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4177_));
OAI21X1 OAI21X1_497 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4177_), .C(AES_CORE_DATAPATH__abc_15863_new_n4178_), .Y(AES_CORE_DATAPATH__0key_0__31_0__28_));
OAI21X1 OAI21X1_498 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4181_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4182_));
OAI21X1 OAI21X1_499 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4182_), .C(AES_CORE_DATAPATH__abc_15863_new_n4183_), .Y(AES_CORE_DATAPATH__0key_0__31_0__29_));
OAI21X1 OAI21X1_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n105_));
OAI21X1 OAI21X1_50 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2538_));
OAI21X1 OAI21X1_500 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4186_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4187_));
OAI21X1 OAI21X1_501 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4187_), .C(AES_CORE_DATAPATH__abc_15863_new_n4188_), .Y(AES_CORE_DATAPATH__0key_0__31_0__30_));
OAI21X1 OAI21X1_502 ( .A(\key_en[0] ), .B(AES_CORE_DATAPATH_key_host_0__31_), .C(AES_CORE_DATAPATH__abc_15863_new_n4190_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4191_));
OAI21X1 OAI21X1_503 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4192_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4193_));
OAI21X1 OAI21X1_504 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4034_), .B(AES_CORE_DATAPATH__abc_15863_new_n4193_), .C(AES_CORE_DATAPATH__abc_15863_new_n4194_), .Y(AES_CORE_DATAPATH__0key_0__31_0__31_));
OAI21X1 OAI21X1_505 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .B(AES_CORE_DATAPATH__abc_15863_new_n4035_), .C(AES_CORE_DATAPATH__abc_15863_new_n4196_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__0_));
OAI21X1 OAI21X1_506 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__0_), .C(AES_CORE_DATAPATH__abc_15863_new_n4232_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4233_));
OAI21X1 OAI21X1_507 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .B(AES_CORE_DATAPATH__abc_15863_new_n4233_), .C(AES_CORE_DATAPATH__abc_15863_new_n4230_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__0_));
OAI21X1 OAI21X1_508 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__1_), .C(AES_CORE_DATAPATH__abc_15863_new_n4237_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4238_));
OAI21X1 OAI21X1_509 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__2_), .C(AES_CORE_DATAPATH__abc_15863_new_n4242_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4243_));
OAI21X1 OAI21X1_51 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2539_), .C(AES_CORE_DATAPATH__abc_15863_new_n2541_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2542_));
OAI21X1 OAI21X1_510 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__3_), .C(AES_CORE_DATAPATH__abc_15863_new_n4247_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4248_));
OAI21X1 OAI21X1_511 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__4_), .C(AES_CORE_DATAPATH__abc_15863_new_n4252_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4253_));
OAI21X1 OAI21X1_512 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__5_), .C(AES_CORE_DATAPATH__abc_15863_new_n4257_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4258_));
OAI21X1 OAI21X1_513 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__12_), .C(AES_CORE_DATAPATH__abc_15863_new_n4280_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4281_));
OAI21X1 OAI21X1_514 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__13_), .C(AES_CORE_DATAPATH__abc_15863_new_n4285_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4286_));
OAI21X1 OAI21X1_515 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__14_), .C(AES_CORE_DATAPATH__abc_15863_new_n4290_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4291_));
OAI21X1 OAI21X1_516 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__15_), .C(AES_CORE_DATAPATH__abc_15863_new_n4295_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4296_));
OAI21X1 OAI21X1_517 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__16_), .C(AES_CORE_DATAPATH__abc_15863_new_n4300_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4301_));
OAI21X1 OAI21X1_518 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__17_), .C(AES_CORE_DATAPATH__abc_15863_new_n4305_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4306_));
OAI21X1 OAI21X1_519 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__18_), .C(AES_CORE_DATAPATH__abc_15863_new_n4310_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4311_));
OAI21X1 OAI21X1_52 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2536_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2542_), .Y(\iv_out[8] ));
OAI21X1 OAI21X1_520 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__19_), .C(AES_CORE_DATAPATH__abc_15863_new_n4315_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4316_));
OAI21X1 OAI21X1_521 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__20_), .C(AES_CORE_DATAPATH__abc_15863_new_n4320_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4321_));
OAI21X1 OAI21X1_522 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__21_), .C(AES_CORE_DATAPATH__abc_15863_new_n4325_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4326_));
OAI21X1 OAI21X1_523 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__22_), .C(AES_CORE_DATAPATH__abc_15863_new_n4330_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4331_));
OAI21X1 OAI21X1_524 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__23_), .C(AES_CORE_DATAPATH__abc_15863_new_n4335_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4336_));
OAI21X1 OAI21X1_525 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__24_), .C(AES_CORE_DATAPATH__abc_15863_new_n4340_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4341_));
OAI21X1 OAI21X1_526 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__25_), .C(AES_CORE_DATAPATH__abc_15863_new_n4345_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4346_));
OAI21X1 OAI21X1_527 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__26_), .C(AES_CORE_DATAPATH__abc_15863_new_n4350_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4351_));
OAI21X1 OAI21X1_528 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__27_), .C(AES_CORE_DATAPATH__abc_15863_new_n4355_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4356_));
OAI21X1 OAI21X1_529 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__28_), .C(AES_CORE_DATAPATH__abc_15863_new_n4360_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4361_));
OAI21X1 OAI21X1_53 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2546_));
OAI21X1 OAI21X1_530 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__29_), .C(AES_CORE_DATAPATH__abc_15863_new_n4365_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4366_));
OAI21X1 OAI21X1_531 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__30_), .C(AES_CORE_DATAPATH__abc_15863_new_n4370_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4371_));
OAI21X1 OAI21X1_532 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .B(AES_CORE_DATAPATH__abc_15863_new_n3868_), .C(AES_CORE_DATAPATH__abc_15863_new_n4376_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__0_));
OAI21X1 OAI21X1_533 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4443_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4444_));
OAI21X1 OAI21X1_534 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4444_), .C(AES_CORE_DATAPATH__abc_15863_new_n4445_), .Y(AES_CORE_DATAPATH__0key_2__31_0__0_));
OAI21X1 OAI21X1_535 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4447_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4448_));
OAI21X1 OAI21X1_536 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4448_), .C(AES_CORE_DATAPATH__abc_15863_new_n4449_), .Y(AES_CORE_DATAPATH__0key_2__31_0__1_));
OAI21X1 OAI21X1_537 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4451_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4452_));
OAI21X1 OAI21X1_538 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4452_), .C(AES_CORE_DATAPATH__abc_15863_new_n4453_), .Y(AES_CORE_DATAPATH__0key_2__31_0__2_));
OAI21X1 OAI21X1_539 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4455_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4456_));
OAI21X1 OAI21X1_54 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2547_), .C(AES_CORE_DATAPATH__abc_15863_new_n2549_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2550_));
OAI21X1 OAI21X1_540 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4456_), .C(AES_CORE_DATAPATH__abc_15863_new_n4457_), .Y(AES_CORE_DATAPATH__0key_2__31_0__3_));
OAI21X1 OAI21X1_541 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4459_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4460_));
OAI21X1 OAI21X1_542 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4460_), .C(AES_CORE_DATAPATH__abc_15863_new_n4461_), .Y(AES_CORE_DATAPATH__0key_2__31_0__4_));
OAI21X1 OAI21X1_543 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4463_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4464_));
OAI21X1 OAI21X1_544 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4464_), .C(AES_CORE_DATAPATH__abc_15863_new_n4465_), .Y(AES_CORE_DATAPATH__0key_2__31_0__5_));
OAI21X1 OAI21X1_545 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4467_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4468_));
OAI21X1 OAI21X1_546 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4468_), .C(AES_CORE_DATAPATH__abc_15863_new_n4469_), .Y(AES_CORE_DATAPATH__0key_2__31_0__6_));
OAI21X1 OAI21X1_547 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4471_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4472_));
OAI21X1 OAI21X1_548 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4472_), .C(AES_CORE_DATAPATH__abc_15863_new_n4473_), .Y(AES_CORE_DATAPATH__0key_2__31_0__7_));
OAI21X1 OAI21X1_549 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4475_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4476_));
OAI21X1 OAI21X1_55 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2544_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2550_), .Y(\iv_out[9] ));
OAI21X1 OAI21X1_550 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4476_), .C(AES_CORE_DATAPATH__abc_15863_new_n4477_), .Y(AES_CORE_DATAPATH__0key_2__31_0__8_));
OAI21X1 OAI21X1_551 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4479_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4480_));
OAI21X1 OAI21X1_552 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4480_), .C(AES_CORE_DATAPATH__abc_15863_new_n4481_), .Y(AES_CORE_DATAPATH__0key_2__31_0__9_));
OAI21X1 OAI21X1_553 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4483_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4484_));
OAI21X1 OAI21X1_554 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4484_), .C(AES_CORE_DATAPATH__abc_15863_new_n4485_), .Y(AES_CORE_DATAPATH__0key_2__31_0__10_));
OAI21X1 OAI21X1_555 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4487_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4488_));
OAI21X1 OAI21X1_556 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4488_), .C(AES_CORE_DATAPATH__abc_15863_new_n4489_), .Y(AES_CORE_DATAPATH__0key_2__31_0__11_));
OAI21X1 OAI21X1_557 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4491_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4492_));
OAI21X1 OAI21X1_558 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4492_), .C(AES_CORE_DATAPATH__abc_15863_new_n4493_), .Y(AES_CORE_DATAPATH__0key_2__31_0__12_));
OAI21X1 OAI21X1_559 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4495_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4496_));
OAI21X1 OAI21X1_56 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2554_));
OAI21X1 OAI21X1_560 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4496_), .C(AES_CORE_DATAPATH__abc_15863_new_n4497_), .Y(AES_CORE_DATAPATH__0key_2__31_0__13_));
OAI21X1 OAI21X1_561 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4500_));
OAI21X1 OAI21X1_562 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4500_), .C(AES_CORE_DATAPATH__abc_15863_new_n4501_), .Y(AES_CORE_DATAPATH__0key_2__31_0__14_));
OAI21X1 OAI21X1_563 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4503_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4504_));
OAI21X1 OAI21X1_564 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4504_), .C(AES_CORE_DATAPATH__abc_15863_new_n4505_), .Y(AES_CORE_DATAPATH__0key_2__31_0__15_));
OAI21X1 OAI21X1_565 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4507_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4508_));
OAI21X1 OAI21X1_566 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4508_), .C(AES_CORE_DATAPATH__abc_15863_new_n4509_), .Y(AES_CORE_DATAPATH__0key_2__31_0__16_));
OAI21X1 OAI21X1_567 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4511_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4512_));
OAI21X1 OAI21X1_568 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4512_), .C(AES_CORE_DATAPATH__abc_15863_new_n4513_), .Y(AES_CORE_DATAPATH__0key_2__31_0__17_));
OAI21X1 OAI21X1_569 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4515_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4516_));
OAI21X1 OAI21X1_57 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2555_), .C(AES_CORE_DATAPATH__abc_15863_new_n2557_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2558_));
OAI21X1 OAI21X1_570 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4516_), .C(AES_CORE_DATAPATH__abc_15863_new_n4517_), .Y(AES_CORE_DATAPATH__0key_2__31_0__18_));
OAI21X1 OAI21X1_571 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4519_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4520_));
OAI21X1 OAI21X1_572 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4520_), .C(AES_CORE_DATAPATH__abc_15863_new_n4521_), .Y(AES_CORE_DATAPATH__0key_2__31_0__19_));
OAI21X1 OAI21X1_573 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4523_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4524_));
OAI21X1 OAI21X1_574 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4524_), .C(AES_CORE_DATAPATH__abc_15863_new_n4525_), .Y(AES_CORE_DATAPATH__0key_2__31_0__20_));
OAI21X1 OAI21X1_575 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4527_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4528_));
OAI21X1 OAI21X1_576 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4528_), .C(AES_CORE_DATAPATH__abc_15863_new_n4529_), .Y(AES_CORE_DATAPATH__0key_2__31_0__21_));
OAI21X1 OAI21X1_577 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4531_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4532_));
OAI21X1 OAI21X1_578 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4532_), .C(AES_CORE_DATAPATH__abc_15863_new_n4533_), .Y(AES_CORE_DATAPATH__0key_2__31_0__22_));
OAI21X1 OAI21X1_579 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4535_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4536_));
OAI21X1 OAI21X1_58 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2552_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2558_), .Y(\iv_out[10] ));
OAI21X1 OAI21X1_580 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4536_), .C(AES_CORE_DATAPATH__abc_15863_new_n4537_), .Y(AES_CORE_DATAPATH__0key_2__31_0__23_));
OAI21X1 OAI21X1_581 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4539_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4540_));
OAI21X1 OAI21X1_582 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4540_), .C(AES_CORE_DATAPATH__abc_15863_new_n4541_), .Y(AES_CORE_DATAPATH__0key_2__31_0__24_));
OAI21X1 OAI21X1_583 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4543_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4544_));
OAI21X1 OAI21X1_584 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4544_), .C(AES_CORE_DATAPATH__abc_15863_new_n4545_), .Y(AES_CORE_DATAPATH__0key_2__31_0__25_));
OAI21X1 OAI21X1_585 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4547_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4548_));
OAI21X1 OAI21X1_586 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4548_), .C(AES_CORE_DATAPATH__abc_15863_new_n4549_), .Y(AES_CORE_DATAPATH__0key_2__31_0__26_));
OAI21X1 OAI21X1_587 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4551_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4552_));
OAI21X1 OAI21X1_588 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4552_), .C(AES_CORE_DATAPATH__abc_15863_new_n4553_), .Y(AES_CORE_DATAPATH__0key_2__31_0__27_));
OAI21X1 OAI21X1_589 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4555_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4556_));
OAI21X1 OAI21X1_59 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2562_));
OAI21X1 OAI21X1_590 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4556_), .C(AES_CORE_DATAPATH__abc_15863_new_n4557_), .Y(AES_CORE_DATAPATH__0key_2__31_0__28_));
OAI21X1 OAI21X1_591 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4559_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4560_));
OAI21X1 OAI21X1_592 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4560_), .C(AES_CORE_DATAPATH__abc_15863_new_n4561_), .Y(AES_CORE_DATAPATH__0key_2__31_0__29_));
OAI21X1 OAI21X1_593 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4563_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4564_));
OAI21X1 OAI21X1_594 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4564_), .C(AES_CORE_DATAPATH__abc_15863_new_n4565_), .Y(AES_CORE_DATAPATH__0key_2__31_0__30_));
OAI21X1 OAI21X1_595 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_), .B(AES_CORE_DATAPATH__abc_15863_new_n3867_), .C(AES_CORE_DATAPATH__abc_15863_new_n4567_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4568_));
OAI21X1 OAI21X1_596 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4442_), .B(AES_CORE_DATAPATH__abc_15863_new_n4568_), .C(AES_CORE_DATAPATH__abc_15863_new_n4569_), .Y(AES_CORE_DATAPATH__0key_2__31_0__31_));
OAI21X1 OAI21X1_597 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n4573_), .C(AES_CORE_DATAPATH__abc_15863_new_n4574_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4575_));
OAI21X1 OAI21X1_598 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH__abc_15863_new_n4576_), .C(AES_CORE_DATAPATH__abc_15863_new_n4577_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4578_));
OAI21X1 OAI21X1_599 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2740_), .B(AES_CORE_DATAPATH__abc_15863_new_n3104_), .C(AES_CORE_DATAPATH__abc_15863_new_n4589_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4590_));
OAI21X1 OAI21X1_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_));
OAI21X1 OAI21X1_60 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2468_), .B(AES_CORE_DATAPATH__abc_15863_new_n2563_), .C(AES_CORE_DATAPATH__abc_15863_new_n2565_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2566_));
OAI21X1 OAI21X1_600 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4600_));
OAI21X1 OAI21X1_601 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4601_));
OAI21X1 OAI21X1_602 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4601_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4600_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4602_));
OAI21X1 OAI21X1_603 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4599_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4603_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4604_));
OAI21X1 OAI21X1_604 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4605_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4606_));
OAI21X1 OAI21X1_605 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4604_), .C(AES_CORE_DATAPATH__abc_15863_new_n4606_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4607_));
OAI21X1 OAI21X1_606 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4607_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4608_));
OAI21X1 OAI21X1_607 ( .A(\iv_out[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4608_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4609_));
OAI21X1 OAI21X1_608 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3110_), .B(AES_CORE_DATAPATH__abc_15863_new_n3106_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4611_));
OAI21X1 OAI21X1_609 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4607_), .C(AES_CORE_DATAPATH__abc_15863_new_n4614_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4615_));
OAI21X1 OAI21X1_61 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2560_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2566_), .Y(\iv_out[11] ));
OAI21X1 OAI21X1_610 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[0] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4619_));
OAI21X1 OAI21X1_611 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4625_));
OAI21X1 OAI21X1_612 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4625_), .B(AES_CORE_DATAPATH__abc_15863_new_n4622_), .C(AES_CORE_DATAPATH__abc_15863_new_n4627_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4628_));
OAI21X1 OAI21X1_613 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4620_), .B(AES_CORE_DATAPATH__abc_15863_new_n4628_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4629_));
OAI21X1 OAI21X1_614 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4631_), .C(AES_CORE_DATAPATH__abc_15863_new_n4572_), .Y(AES_CORE_DATAPATH__0col_0__31_0__0_));
OAI21X1 OAI21X1_615 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3133_), .B(AES_CORE_DATAPATH__abc_15863_new_n3130_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4637_));
OAI21X1 OAI21X1_616 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4641_));
OAI21X1 OAI21X1_617 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4642_));
OAI21X1 OAI21X1_618 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4642_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4641_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4643_));
OAI21X1 OAI21X1_619 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4640_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4644_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4645_));
OAI21X1 OAI21X1_62 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2569_));
OAI21X1 OAI21X1_620 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4646_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4647_));
OAI21X1 OAI21X1_621 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4645_), .C(AES_CORE_DATAPATH__abc_15863_new_n4647_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4648_));
OAI21X1 OAI21X1_622 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4648_), .C(AES_CORE_DATAPATH__abc_15863_new_n4649_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4650_));
OAI21X1 OAI21X1_623 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4648_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4657_));
OAI21X1 OAI21X1_624 ( .A(\iv_out[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4657_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4658_));
OAI21X1 OAI21X1_625 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4638_), .B(AES_CORE_DATAPATH__abc_15863_new_n4656_), .C(AES_CORE_DATAPATH__abc_15863_new_n4658_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4659_));
OAI21X1 OAI21X1_626 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[1] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4661_));
OAI21X1 OAI21X1_627 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4664_));
OAI21X1 OAI21X1_628 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4664_), .B(AES_CORE_DATAPATH__abc_15863_new_n4663_), .C(AES_CORE_DATAPATH__abc_15863_new_n4665_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4666_));
OAI21X1 OAI21X1_629 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4662_), .B(AES_CORE_DATAPATH__abc_15863_new_n4666_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4667_));
OAI21X1 OAI21X1_63 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2569_), .C(AES_CORE_DATAPATH__abc_15863_new_n2570_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2571_));
OAI21X1 OAI21X1_630 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4670_), .C(AES_CORE_DATAPATH__abc_15863_new_n4633_), .Y(AES_CORE_DATAPATH__0col_0__31_0__1_));
OAI21X1 OAI21X1_631 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2764_), .B(AES_CORE_DATAPATH__abc_15863_new_n3150_), .C(AES_CORE_DATAPATH__abc_15863_new_n4676_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4677_));
OAI21X1 OAI21X1_632 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4682_));
OAI21X1 OAI21X1_633 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4683_));
OAI21X1 OAI21X1_634 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4683_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4682_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4684_));
OAI21X1 OAI21X1_635 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4681_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4685_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4686_));
OAI21X1 OAI21X1_636 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4687_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4688_));
OAI21X1 OAI21X1_637 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4686_), .C(AES_CORE_DATAPATH__abc_15863_new_n4688_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4689_));
OAI21X1 OAI21X1_638 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4689_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4690_));
OAI21X1 OAI21X1_639 ( .A(\iv_out[2] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4690_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4691_));
OAI21X1 OAI21X1_64 ( .A(AES_CORE_DATAPATH_iv_2__12_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2572_));
OAI21X1 OAI21X1_640 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3155_), .B(AES_CORE_DATAPATH__abc_15863_new_n3152_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4693_));
OAI21X1 OAI21X1_641 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4689_), .C(AES_CORE_DATAPATH__abc_15863_new_n4696_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4697_));
OAI21X1 OAI21X1_642 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[2] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4700_));
OAI21X1 OAI21X1_643 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4703_));
OAI21X1 OAI21X1_644 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4703_), .B(AES_CORE_DATAPATH__abc_15863_new_n4702_), .C(AES_CORE_DATAPATH__abc_15863_new_n4704_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4705_));
OAI21X1 OAI21X1_645 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4701_), .B(AES_CORE_DATAPATH__abc_15863_new_n4705_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4706_));
OAI21X1 OAI21X1_646 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4709_), .C(AES_CORE_DATAPATH__abc_15863_new_n4672_), .Y(AES_CORE_DATAPATH__0col_0__31_0__2_));
OAI21X1 OAI21X1_647 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3178_), .B(AES_CORE_DATAPATH__abc_15863_new_n4717_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4718_));
OAI21X1 OAI21X1_648 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4722_));
OAI21X1 OAI21X1_649 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4723_));
OAI21X1 OAI21X1_65 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2575_));
OAI21X1 OAI21X1_650 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4723_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4722_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4724_));
OAI21X1 OAI21X1_651 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4721_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4725_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4726_));
OAI21X1 OAI21X1_652 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4727_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4728_));
OAI21X1 OAI21X1_653 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4726_), .C(AES_CORE_DATAPATH__abc_15863_new_n4728_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4729_));
OAI21X1 OAI21X1_654 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4729_), .C(AES_CORE_DATAPATH__abc_15863_new_n4730_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4731_));
OAI21X1 OAI21X1_655 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4729_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4734_));
OAI21X1 OAI21X1_656 ( .A(\iv_out[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4734_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4735_));
OAI21X1 OAI21X1_657 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4719_), .B(AES_CORE_DATAPATH__abc_15863_new_n4733_), .C(AES_CORE_DATAPATH__abc_15863_new_n4735_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4736_));
OAI21X1 OAI21X1_658 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[3] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4738_));
OAI21X1 OAI21X1_659 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4741_));
OAI21X1 OAI21X1_66 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2575_), .C(AES_CORE_DATAPATH__abc_15863_new_n2576_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2577_));
OAI21X1 OAI21X1_660 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4741_), .B(AES_CORE_DATAPATH__abc_15863_new_n4740_), .C(AES_CORE_DATAPATH__abc_15863_new_n4742_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4743_));
OAI21X1 OAI21X1_661 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4739_), .B(AES_CORE_DATAPATH__abc_15863_new_n4743_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4744_));
OAI21X1 OAI21X1_662 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4749_), .C(AES_CORE_DATAPATH__abc_15863_new_n4711_), .Y(AES_CORE_DATAPATH__0col_0__31_0__3_));
OAI21X1 OAI21X1_663 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2784_), .B(AES_CORE_DATAPATH__abc_15863_new_n3195_), .C(AES_CORE_DATAPATH__abc_15863_new_n4755_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4756_));
OAI21X1 OAI21X1_664 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4760_));
OAI21X1 OAI21X1_665 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n4760_), .C(AES_CORE_DATAPATH__abc_15863_new_n4761_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4762_));
OAI21X1 OAI21X1_666 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4765_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4766_));
OAI21X1 OAI21X1_667 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4598_), .B(\iv_out[4] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4766_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4767_));
OAI21X1 OAI21X1_668 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3200_), .B(AES_CORE_DATAPATH__abc_15863_new_n3197_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4769_));
OAI21X1 OAI21X1_669 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4765_), .C(AES_CORE_DATAPATH__abc_15863_new_n4772_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4773_));
OAI21X1 OAI21X1_67 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2574_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2580_), .Y(\iv_out[13] ));
OAI21X1 OAI21X1_670 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[4] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4776_));
OAI21X1 OAI21X1_671 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4779_));
OAI21X1 OAI21X1_672 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4779_), .B(AES_CORE_DATAPATH__abc_15863_new_n4778_), .C(AES_CORE_DATAPATH__abc_15863_new_n4780_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4781_));
OAI21X1 OAI21X1_673 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4777_), .B(AES_CORE_DATAPATH__abc_15863_new_n4781_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4782_));
OAI21X1 OAI21X1_674 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4785_), .C(AES_CORE_DATAPATH__abc_15863_new_n4751_), .Y(AES_CORE_DATAPATH__0col_0__31_0__4_));
OAI21X1 OAI21X1_675 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2794_), .B(AES_CORE_DATAPATH__abc_15863_new_n3217_), .C(AES_CORE_DATAPATH__abc_15863_new_n4791_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4792_));
OAI21X1 OAI21X1_676 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4797_));
OAI21X1 OAI21X1_677 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4798_));
OAI21X1 OAI21X1_678 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4798_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4797_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4799_));
OAI21X1 OAI21X1_679 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4796_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4800_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4801_));
OAI21X1 OAI21X1_68 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2583_));
OAI21X1 OAI21X1_680 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4802_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4803_));
OAI21X1 OAI21X1_681 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4801_), .C(AES_CORE_DATAPATH__abc_15863_new_n4803_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4804_));
OAI21X1 OAI21X1_682 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4804_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4805_));
OAI21X1 OAI21X1_683 ( .A(\iv_out[5] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4805_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4806_));
OAI21X1 OAI21X1_684 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3222_), .B(AES_CORE_DATAPATH__abc_15863_new_n3219_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4808_));
OAI21X1 OAI21X1_685 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4804_), .C(AES_CORE_DATAPATH__abc_15863_new_n4811_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4812_));
OAI21X1 OAI21X1_686 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[5] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4815_));
OAI21X1 OAI21X1_687 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4818_));
OAI21X1 OAI21X1_688 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4818_), .B(AES_CORE_DATAPATH__abc_15863_new_n4817_), .C(AES_CORE_DATAPATH__abc_15863_new_n4819_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4820_));
OAI21X1 OAI21X1_689 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4816_), .B(AES_CORE_DATAPATH__abc_15863_new_n4820_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4821_));
OAI21X1 OAI21X1_69 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2583_), .C(AES_CORE_DATAPATH__abc_15863_new_n2584_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2585_));
OAI21X1 OAI21X1_690 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4824_), .C(AES_CORE_DATAPATH__abc_15863_new_n4787_), .Y(AES_CORE_DATAPATH__0col_0__31_0__5_));
OAI21X1 OAI21X1_691 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2804_), .B(AES_CORE_DATAPATH__abc_15863_new_n3239_), .C(AES_CORE_DATAPATH__abc_15863_new_n4830_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4831_));
OAI21X1 OAI21X1_692 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4835_));
OAI21X1 OAI21X1_693 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n4835_), .C(AES_CORE_DATAPATH__abc_15863_new_n4836_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4837_));
OAI21X1 OAI21X1_694 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4840_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4841_));
OAI21X1 OAI21X1_695 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4598_), .B(\iv_out[6] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4841_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4842_));
OAI21X1 OAI21X1_696 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3244_), .B(AES_CORE_DATAPATH__abc_15863_new_n3241_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4844_));
OAI21X1 OAI21X1_697 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[6] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4850_));
OAI21X1 OAI21X1_698 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4853_));
OAI21X1 OAI21X1_699 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4853_), .B(AES_CORE_DATAPATH__abc_15863_new_n4852_), .C(AES_CORE_DATAPATH__abc_15863_new_n4854_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4855_));
OAI21X1 OAI21X1_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_), .B(start), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n112_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_0_));
OAI21X1 OAI21X1_70 ( .A(AES_CORE_DATAPATH_iv_2__14_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2585_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2586_));
OAI21X1 OAI21X1_700 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4851_), .B(AES_CORE_DATAPATH__abc_15863_new_n4855_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4856_));
OAI21X1 OAI21X1_701 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4859_), .C(AES_CORE_DATAPATH__abc_15863_new_n4826_), .Y(AES_CORE_DATAPATH__0col_0__31_0__6_));
OAI21X1 OAI21X1_702 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3266_), .B(AES_CORE_DATAPATH__abc_15863_new_n3263_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4865_));
OAI21X1 OAI21X1_703 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4869_));
OAI21X1 OAI21X1_704 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4870_));
OAI21X1 OAI21X1_705 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4870_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4869_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4871_));
OAI21X1 OAI21X1_706 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4868_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4872_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4873_));
OAI21X1 OAI21X1_707 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4874_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4875_));
OAI21X1 OAI21X1_708 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4873_), .C(AES_CORE_DATAPATH__abc_15863_new_n4875_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4876_));
OAI21X1 OAI21X1_709 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4876_), .C(AES_CORE_DATAPATH__abc_15863_new_n4877_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4878_));
OAI21X1 OAI21X1_71 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2589_));
OAI21X1 OAI21X1_710 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4876_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4885_));
OAI21X1 OAI21X1_711 ( .A(\iv_out[7] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4885_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4886_));
OAI21X1 OAI21X1_712 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4866_), .B(AES_CORE_DATAPATH__abc_15863_new_n4884_), .C(AES_CORE_DATAPATH__abc_15863_new_n4886_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4887_));
OAI21X1 OAI21X1_713 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[7] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4889_));
OAI21X1 OAI21X1_714 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4892_));
OAI21X1 OAI21X1_715 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4892_), .B(AES_CORE_DATAPATH__abc_15863_new_n4891_), .C(AES_CORE_DATAPATH__abc_15863_new_n4893_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4894_));
OAI21X1 OAI21X1_716 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4890_), .B(AES_CORE_DATAPATH__abc_15863_new_n4894_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4895_));
OAI21X1 OAI21X1_717 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4898_), .C(AES_CORE_DATAPATH__abc_15863_new_n4861_), .Y(AES_CORE_DATAPATH__0col_0__31_0__7_));
OAI21X1 OAI21X1_718 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2828_), .B(AES_CORE_DATAPATH__abc_15863_new_n3283_), .C(AES_CORE_DATAPATH__abc_15863_new_n4904_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4905_));
OAI21X1 OAI21X1_719 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__8_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4909_));
OAI21X1 OAI21X1_72 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2589_), .C(AES_CORE_DATAPATH__abc_15863_new_n2590_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2591_));
OAI21X1 OAI21X1_720 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n4909_), .C(AES_CORE_DATAPATH__abc_15863_new_n4910_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4911_));
OAI21X1 OAI21X1_721 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4914_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4915_));
OAI21X1 OAI21X1_722 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4598_), .B(\iv_out[8] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4915_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4916_));
OAI21X1 OAI21X1_723 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3288_), .B(AES_CORE_DATAPATH__abc_15863_new_n3285_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4918_));
OAI21X1 OAI21X1_724 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[8] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4924_));
OAI21X1 OAI21X1_725 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4927_));
OAI21X1 OAI21X1_726 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4927_), .B(AES_CORE_DATAPATH__abc_15863_new_n4926_), .C(AES_CORE_DATAPATH__abc_15863_new_n4928_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4929_));
OAI21X1 OAI21X1_727 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4925_), .B(AES_CORE_DATAPATH__abc_15863_new_n4929_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4930_));
OAI21X1 OAI21X1_728 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4933_), .C(AES_CORE_DATAPATH__abc_15863_new_n4900_), .Y(AES_CORE_DATAPATH__0col_0__31_0__8_));
OAI21X1 OAI21X1_729 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3310_), .B(AES_CORE_DATAPATH__abc_15863_new_n4941_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4942_));
OAI21X1 OAI21X1_73 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2588_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2594_), .Y(\iv_out[15] ));
OAI21X1 OAI21X1_730 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4946_));
OAI21X1 OAI21X1_731 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__9_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4947_));
OAI21X1 OAI21X1_732 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4947_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4946_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4948_));
OAI21X1 OAI21X1_733 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4945_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4949_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4950_));
OAI21X1 OAI21X1_734 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4951_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4952_));
OAI21X1 OAI21X1_735 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4950_), .C(AES_CORE_DATAPATH__abc_15863_new_n4952_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4953_));
OAI21X1 OAI21X1_736 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4953_), .C(AES_CORE_DATAPATH__abc_15863_new_n4954_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4955_));
OAI21X1 OAI21X1_737 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4953_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4958_));
OAI21X1 OAI21X1_738 ( .A(\iv_out[9] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4958_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4959_));
OAI21X1 OAI21X1_739 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4943_), .B(AES_CORE_DATAPATH__abc_15863_new_n4957_), .C(AES_CORE_DATAPATH__abc_15863_new_n4959_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4960_));
OAI21X1 OAI21X1_74 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2597_));
OAI21X1 OAI21X1_740 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[9] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4962_));
OAI21X1 OAI21X1_741 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n4965_));
OAI21X1 OAI21X1_742 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4965_), .B(AES_CORE_DATAPATH__abc_15863_new_n4964_), .C(AES_CORE_DATAPATH__abc_15863_new_n4966_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4967_));
OAI21X1 OAI21X1_743 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4963_), .B(AES_CORE_DATAPATH__abc_15863_new_n4967_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4968_));
OAI21X1 OAI21X1_744 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n4972_), .C(AES_CORE_DATAPATH__abc_15863_new_n4935_), .Y(AES_CORE_DATAPATH__0col_0__31_0__9_));
OAI21X1 OAI21X1_745 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2851_), .B(AES_CORE_DATAPATH__abc_15863_new_n3327_), .C(AES_CORE_DATAPATH__abc_15863_new_n4978_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4979_));
OAI21X1 OAI21X1_746 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4984_));
OAI21X1 OAI21X1_747 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__10_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4985_));
OAI21X1 OAI21X1_748 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4985_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n4984_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4986_));
OAI21X1 OAI21X1_749 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4983_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n4987_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4988_));
OAI21X1 OAI21X1_75 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2597_), .C(AES_CORE_DATAPATH__abc_15863_new_n2598_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2599_));
OAI21X1 OAI21X1_750 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n4989_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4990_));
OAI21X1 OAI21X1_751 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n4988_), .C(AES_CORE_DATAPATH__abc_15863_new_n4990_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4991_));
OAI21X1 OAI21X1_752 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n4991_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4992_));
OAI21X1 OAI21X1_753 ( .A(\iv_out[10] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4992_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4993_));
OAI21X1 OAI21X1_754 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3332_), .B(AES_CORE_DATAPATH__abc_15863_new_n3329_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4995_));
OAI21X1 OAI21X1_755 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n4991_), .C(AES_CORE_DATAPATH__abc_15863_new_n4998_), .Y(AES_CORE_DATAPATH__abc_15863_new_n4999_));
OAI21X1 OAI21X1_756 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[10] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5002_));
OAI21X1 OAI21X1_757 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5005_));
OAI21X1 OAI21X1_758 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5005_), .B(AES_CORE_DATAPATH__abc_15863_new_n5004_), .C(AES_CORE_DATAPATH__abc_15863_new_n5006_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5007_));
OAI21X1 OAI21X1_759 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5003_), .B(AES_CORE_DATAPATH__abc_15863_new_n5007_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5008_));
OAI21X1 OAI21X1_76 ( .A(AES_CORE_DATAPATH_iv_2__16_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2599_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2600_));
OAI21X1 OAI21X1_760 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5011_), .C(AES_CORE_DATAPATH__abc_15863_new_n4974_), .Y(AES_CORE_DATAPATH__0col_0__31_0__10_));
OAI21X1 OAI21X1_761 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3354_), .B(AES_CORE_DATAPATH__abc_15863_new_n5019_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5020_));
OAI21X1 OAI21X1_762 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5024_));
OAI21X1 OAI21X1_763 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__11_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5025_));
OAI21X1 OAI21X1_764 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5025_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5024_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5026_));
OAI21X1 OAI21X1_765 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5023_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5027_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5028_));
OAI21X1 OAI21X1_766 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5029_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5030_));
OAI21X1 OAI21X1_767 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5028_), .C(AES_CORE_DATAPATH__abc_15863_new_n5030_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5031_));
OAI21X1 OAI21X1_768 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5031_), .C(AES_CORE_DATAPATH__abc_15863_new_n5032_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5033_));
OAI21X1 OAI21X1_769 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5031_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5036_));
OAI21X1 OAI21X1_77 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2603_));
OAI21X1 OAI21X1_770 ( .A(\iv_out[11] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5036_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5037_));
OAI21X1 OAI21X1_771 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5021_), .B(AES_CORE_DATAPATH__abc_15863_new_n5035_), .C(AES_CORE_DATAPATH__abc_15863_new_n5037_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5038_));
OAI21X1 OAI21X1_772 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[11] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5040_));
OAI21X1 OAI21X1_773 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5043_));
OAI21X1 OAI21X1_774 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5043_), .B(AES_CORE_DATAPATH__abc_15863_new_n5042_), .C(AES_CORE_DATAPATH__abc_15863_new_n5044_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5045_));
OAI21X1 OAI21X1_775 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5041_), .B(AES_CORE_DATAPATH__abc_15863_new_n5045_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5046_));
OAI21X1 OAI21X1_776 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5050_), .C(AES_CORE_DATAPATH__abc_15863_new_n5013_), .Y(AES_CORE_DATAPATH__0col_0__31_0__11_));
OAI21X1 OAI21X1_777 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2870_), .B(AES_CORE_DATAPATH__abc_15863_new_n3371_), .C(AES_CORE_DATAPATH__abc_15863_new_n5056_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5057_));
OAI21X1 OAI21X1_778 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5062_));
OAI21X1 OAI21X1_779 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__12_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5063_));
OAI21X1 OAI21X1_78 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2603_), .C(AES_CORE_DATAPATH__abc_15863_new_n2604_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2605_));
OAI21X1 OAI21X1_780 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5063_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5062_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5064_));
OAI21X1 OAI21X1_781 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5061_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5065_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5066_));
OAI21X1 OAI21X1_782 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5067_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5068_));
OAI21X1 OAI21X1_783 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5066_), .C(AES_CORE_DATAPATH__abc_15863_new_n5068_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5069_));
OAI21X1 OAI21X1_784 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5069_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5070_));
OAI21X1 OAI21X1_785 ( .A(\iv_out[12] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5070_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5071_));
OAI21X1 OAI21X1_786 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3376_), .B(AES_CORE_DATAPATH__abc_15863_new_n3373_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5073_));
OAI21X1 OAI21X1_787 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5069_), .C(AES_CORE_DATAPATH__abc_15863_new_n5076_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5077_));
OAI21X1 OAI21X1_788 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[12] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5080_));
OAI21X1 OAI21X1_789 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5083_));
OAI21X1 OAI21X1_79 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2602_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2608_), .Y(\iv_out[17] ));
OAI21X1 OAI21X1_790 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5083_), .B(AES_CORE_DATAPATH__abc_15863_new_n5082_), .C(AES_CORE_DATAPATH__abc_15863_new_n5084_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5085_));
OAI21X1 OAI21X1_791 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5081_), .B(AES_CORE_DATAPATH__abc_15863_new_n5085_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5086_));
OAI21X1 OAI21X1_792 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5089_), .C(AES_CORE_DATAPATH__abc_15863_new_n5052_), .Y(AES_CORE_DATAPATH__0col_0__31_0__12_));
OAI21X1 OAI21X1_793 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3398_), .B(AES_CORE_DATAPATH__abc_15863_new_n5097_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5098_));
OAI21X1 OAI21X1_794 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5102_));
OAI21X1 OAI21X1_795 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__13_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5103_));
OAI21X1 OAI21X1_796 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5103_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5102_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5104_));
OAI21X1 OAI21X1_797 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5101_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5105_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5106_));
OAI21X1 OAI21X1_798 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5107_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5108_));
OAI21X1 OAI21X1_799 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5106_), .C(AES_CORE_DATAPATH__abc_15863_new_n5108_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5109_));
OAI21X1 OAI21X1_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .C(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n126_));
OAI21X1 OAI21X1_80 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2611_));
OAI21X1 OAI21X1_800 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5109_), .C(AES_CORE_DATAPATH__abc_15863_new_n5110_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5111_));
OAI21X1 OAI21X1_801 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5109_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5114_));
OAI21X1 OAI21X1_802 ( .A(\iv_out[13] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5114_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5115_));
OAI21X1 OAI21X1_803 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5099_), .B(AES_CORE_DATAPATH__abc_15863_new_n5113_), .C(AES_CORE_DATAPATH__abc_15863_new_n5115_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5116_));
OAI21X1 OAI21X1_804 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[13] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5118_));
OAI21X1 OAI21X1_805 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5121_));
OAI21X1 OAI21X1_806 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5121_), .B(AES_CORE_DATAPATH__abc_15863_new_n5120_), .C(AES_CORE_DATAPATH__abc_15863_new_n5122_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5123_));
OAI21X1 OAI21X1_807 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5119_), .B(AES_CORE_DATAPATH__abc_15863_new_n5123_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5124_));
OAI21X1 OAI21X1_808 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5128_), .C(AES_CORE_DATAPATH__abc_15863_new_n5091_), .Y(AES_CORE_DATAPATH__0col_0__31_0__13_));
OAI21X1 OAI21X1_809 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2890_), .B(AES_CORE_DATAPATH__abc_15863_new_n3415_), .C(AES_CORE_DATAPATH__abc_15863_new_n5134_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5135_));
OAI21X1 OAI21X1_81 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2611_), .C(AES_CORE_DATAPATH__abc_15863_new_n2612_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2613_));
OAI21X1 OAI21X1_810 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__14_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5139_));
OAI21X1 OAI21X1_811 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n5139_), .C(AES_CORE_DATAPATH__abc_15863_new_n5140_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5141_));
OAI21X1 OAI21X1_812 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5144_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5145_));
OAI21X1 OAI21X1_813 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4598_), .B(\iv_out[14] ), .C(AES_CORE_DATAPATH__abc_15863_new_n5145_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5146_));
OAI21X1 OAI21X1_814 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3420_), .B(AES_CORE_DATAPATH__abc_15863_new_n3417_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5148_));
OAI21X1 OAI21X1_815 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5144_), .C(AES_CORE_DATAPATH__abc_15863_new_n5151_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5152_));
OAI21X1 OAI21X1_816 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[14] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5155_));
OAI21X1 OAI21X1_817 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5158_));
OAI21X1 OAI21X1_818 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5158_), .B(AES_CORE_DATAPATH__abc_15863_new_n5157_), .C(AES_CORE_DATAPATH__abc_15863_new_n5159_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5160_));
OAI21X1 OAI21X1_819 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5156_), .B(AES_CORE_DATAPATH__abc_15863_new_n5160_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5161_));
OAI21X1 OAI21X1_82 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2610_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2616_), .Y(\iv_out[18] ));
OAI21X1 OAI21X1_820 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5164_), .C(AES_CORE_DATAPATH__abc_15863_new_n5130_), .Y(AES_CORE_DATAPATH__0col_0__31_0__14_));
OAI21X1 OAI21X1_821 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3442_), .B(AES_CORE_DATAPATH__abc_15863_new_n5172_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5173_));
OAI21X1 OAI21X1_822 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5177_));
OAI21X1 OAI21X1_823 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__15_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5178_));
OAI21X1 OAI21X1_824 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5178_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5177_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5179_));
OAI21X1 OAI21X1_825 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5176_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5180_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5181_));
OAI21X1 OAI21X1_826 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5182_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5183_));
OAI21X1 OAI21X1_827 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5181_), .C(AES_CORE_DATAPATH__abc_15863_new_n5183_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5184_));
OAI21X1 OAI21X1_828 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5184_), .C(AES_CORE_DATAPATH__abc_15863_new_n5185_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5186_));
OAI21X1 OAI21X1_829 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5184_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5189_));
OAI21X1 OAI21X1_83 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2619_));
OAI21X1 OAI21X1_830 ( .A(\iv_out[15] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5189_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5190_));
OAI21X1 OAI21X1_831 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5174_), .B(AES_CORE_DATAPATH__abc_15863_new_n5188_), .C(AES_CORE_DATAPATH__abc_15863_new_n5190_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5191_));
OAI21X1 OAI21X1_832 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[15] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5193_));
OAI21X1 OAI21X1_833 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5196_));
OAI21X1 OAI21X1_834 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5196_), .B(AES_CORE_DATAPATH__abc_15863_new_n5195_), .C(AES_CORE_DATAPATH__abc_15863_new_n5197_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5198_));
OAI21X1 OAI21X1_835 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5194_), .B(AES_CORE_DATAPATH__abc_15863_new_n5198_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5199_));
OAI21X1 OAI21X1_836 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5203_), .C(AES_CORE_DATAPATH__abc_15863_new_n5166_), .Y(AES_CORE_DATAPATH__0col_0__31_0__15_));
OAI21X1 OAI21X1_837 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2911_), .B(AES_CORE_DATAPATH__abc_15863_new_n3459_), .C(AES_CORE_DATAPATH__abc_15863_new_n5209_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5210_));
OAI21X1 OAI21X1_838 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5215_));
OAI21X1 OAI21X1_839 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__16_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5216_));
OAI21X1 OAI21X1_84 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2619_), .C(AES_CORE_DATAPATH__abc_15863_new_n2620_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2621_));
OAI21X1 OAI21X1_840 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5216_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5215_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5217_));
OAI21X1 OAI21X1_841 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5214_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5218_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5219_));
OAI21X1 OAI21X1_842 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5220_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5221_));
OAI21X1 OAI21X1_843 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5219_), .C(AES_CORE_DATAPATH__abc_15863_new_n5221_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5222_));
OAI21X1 OAI21X1_844 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5222_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5223_));
OAI21X1 OAI21X1_845 ( .A(\iv_out[16] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5223_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5224_));
OAI21X1 OAI21X1_846 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3464_), .B(AES_CORE_DATAPATH__abc_15863_new_n3461_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5226_));
OAI21X1 OAI21X1_847 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5222_), .C(AES_CORE_DATAPATH__abc_15863_new_n5229_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5230_));
OAI21X1 OAI21X1_848 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[16] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5233_));
OAI21X1 OAI21X1_849 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5236_));
OAI21X1 OAI21X1_85 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2618_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2624_), .Y(\iv_out[19] ));
OAI21X1 OAI21X1_850 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5236_), .B(AES_CORE_DATAPATH__abc_15863_new_n5235_), .C(AES_CORE_DATAPATH__abc_15863_new_n5237_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5238_));
OAI21X1 OAI21X1_851 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5234_), .B(AES_CORE_DATAPATH__abc_15863_new_n5238_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5239_));
OAI21X1 OAI21X1_852 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5242_), .C(AES_CORE_DATAPATH__abc_15863_new_n5205_), .Y(AES_CORE_DATAPATH__0col_0__31_0__16_));
OAI21X1 OAI21X1_853 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3486_), .B(AES_CORE_DATAPATH__abc_15863_new_n5250_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5251_));
OAI21X1 OAI21X1_854 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5255_));
OAI21X1 OAI21X1_855 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__17_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5256_));
OAI21X1 OAI21X1_856 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5256_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5255_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5257_));
OAI21X1 OAI21X1_857 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5254_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5258_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5259_));
OAI21X1 OAI21X1_858 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5260_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5261_));
OAI21X1 OAI21X1_859 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5259_), .C(AES_CORE_DATAPATH__abc_15863_new_n5261_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5262_));
OAI21X1 OAI21X1_86 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2627_));
OAI21X1 OAI21X1_860 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5262_), .C(AES_CORE_DATAPATH__abc_15863_new_n5263_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5264_));
OAI21X1 OAI21X1_861 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5262_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5267_));
OAI21X1 OAI21X1_862 ( .A(\iv_out[17] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5267_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5268_));
OAI21X1 OAI21X1_863 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5252_), .B(AES_CORE_DATAPATH__abc_15863_new_n5266_), .C(AES_CORE_DATAPATH__abc_15863_new_n5268_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5269_));
OAI21X1 OAI21X1_864 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[17] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5271_));
OAI21X1 OAI21X1_865 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5274_));
OAI21X1 OAI21X1_866 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5274_), .B(AES_CORE_DATAPATH__abc_15863_new_n5273_), .C(AES_CORE_DATAPATH__abc_15863_new_n5275_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5276_));
OAI21X1 OAI21X1_867 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5272_), .B(AES_CORE_DATAPATH__abc_15863_new_n5276_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5277_));
OAI21X1 OAI21X1_868 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5281_), .C(AES_CORE_DATAPATH__abc_15863_new_n5244_), .Y(AES_CORE_DATAPATH__0col_0__31_0__17_));
OAI21X1 OAI21X1_869 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3508_), .B(AES_CORE_DATAPATH__abc_15863_new_n5289_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5290_));
OAI21X1 OAI21X1_87 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2627_), .C(AES_CORE_DATAPATH__abc_15863_new_n2628_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2629_));
OAI21X1 OAI21X1_870 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5294_));
OAI21X1 OAI21X1_871 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__18_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5295_));
OAI21X1 OAI21X1_872 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5295_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5294_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5296_));
OAI21X1 OAI21X1_873 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5293_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5297_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5298_));
OAI21X1 OAI21X1_874 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5299_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5300_));
OAI21X1 OAI21X1_875 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5298_), .C(AES_CORE_DATAPATH__abc_15863_new_n5300_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5301_));
OAI21X1 OAI21X1_876 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5301_), .C(AES_CORE_DATAPATH__abc_15863_new_n5302_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5303_));
OAI21X1 OAI21X1_877 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5301_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5306_));
OAI21X1 OAI21X1_878 ( .A(\iv_out[18] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5306_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5307_));
OAI21X1 OAI21X1_879 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5291_), .B(AES_CORE_DATAPATH__abc_15863_new_n5305_), .C(AES_CORE_DATAPATH__abc_15863_new_n5307_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5308_));
OAI21X1 OAI21X1_88 ( .A(AES_CORE_DATAPATH_iv_2__20_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2629_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2630_));
OAI21X1 OAI21X1_880 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[18] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5310_));
OAI21X1 OAI21X1_881 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5313_));
OAI21X1 OAI21X1_882 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5313_), .B(AES_CORE_DATAPATH__abc_15863_new_n5312_), .C(AES_CORE_DATAPATH__abc_15863_new_n5314_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5315_));
OAI21X1 OAI21X1_883 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5311_), .B(AES_CORE_DATAPATH__abc_15863_new_n5315_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5316_));
OAI21X1 OAI21X1_884 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5320_), .C(AES_CORE_DATAPATH__abc_15863_new_n5283_), .Y(AES_CORE_DATAPATH__0col_0__31_0__18_));
OAI21X1 OAI21X1_885 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3530_), .B(AES_CORE_DATAPATH__abc_15863_new_n5328_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5329_));
OAI21X1 OAI21X1_886 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5333_));
OAI21X1 OAI21X1_887 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__19_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5334_));
OAI21X1 OAI21X1_888 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5334_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5333_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5335_));
OAI21X1 OAI21X1_889 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5332_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5336_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5337_));
OAI21X1 OAI21X1_89 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2633_));
OAI21X1 OAI21X1_890 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5338_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5339_));
OAI21X1 OAI21X1_891 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5337_), .C(AES_CORE_DATAPATH__abc_15863_new_n5339_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5340_));
OAI21X1 OAI21X1_892 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5340_), .C(AES_CORE_DATAPATH__abc_15863_new_n5341_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5342_));
OAI21X1 OAI21X1_893 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5340_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5345_));
OAI21X1 OAI21X1_894 ( .A(\iv_out[19] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5345_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5346_));
OAI21X1 OAI21X1_895 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5330_), .B(AES_CORE_DATAPATH__abc_15863_new_n5344_), .C(AES_CORE_DATAPATH__abc_15863_new_n5346_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5347_));
OAI21X1 OAI21X1_896 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[19] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5349_));
OAI21X1 OAI21X1_897 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5352_));
OAI21X1 OAI21X1_898 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5352_), .B(AES_CORE_DATAPATH__abc_15863_new_n5351_), .C(AES_CORE_DATAPATH__abc_15863_new_n5353_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5354_));
OAI21X1 OAI21X1_899 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5350_), .B(AES_CORE_DATAPATH__abc_15863_new_n5354_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5355_));
OAI21X1 OAI21X1_9 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n88_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n126_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n127_));
OAI21X1 OAI21X1_90 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2633_), .C(AES_CORE_DATAPATH__abc_15863_new_n2634_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2635_));
OAI21X1 OAI21X1_900 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5359_), .C(AES_CORE_DATAPATH__abc_15863_new_n5322_), .Y(AES_CORE_DATAPATH__0col_0__31_0__19_));
OAI21X1 OAI21X1_901 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2951_), .B(AES_CORE_DATAPATH__abc_15863_new_n3547_), .C(AES_CORE_DATAPATH__abc_15863_new_n5365_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5366_));
OAI21X1 OAI21X1_902 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5371_));
OAI21X1 OAI21X1_903 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__20_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5372_));
OAI21X1 OAI21X1_904 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5372_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5371_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5373_));
OAI21X1 OAI21X1_905 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5370_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5374_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5375_));
OAI21X1 OAI21X1_906 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5376_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5377_));
OAI21X1 OAI21X1_907 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5375_), .C(AES_CORE_DATAPATH__abc_15863_new_n5377_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5378_));
OAI21X1 OAI21X1_908 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5378_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5379_));
OAI21X1 OAI21X1_909 ( .A(\iv_out[20] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5379_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5380_));
OAI21X1 OAI21X1_91 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2632_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2638_), .Y(\iv_out[21] ));
OAI21X1 OAI21X1_910 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3552_), .B(AES_CORE_DATAPATH__abc_15863_new_n3549_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5382_));
OAI21X1 OAI21X1_911 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5378_), .C(AES_CORE_DATAPATH__abc_15863_new_n5385_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5386_));
OAI21X1 OAI21X1_912 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[20] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5389_));
OAI21X1 OAI21X1_913 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5392_));
OAI21X1 OAI21X1_914 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5392_), .B(AES_CORE_DATAPATH__abc_15863_new_n5391_), .C(AES_CORE_DATAPATH__abc_15863_new_n5393_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5394_));
OAI21X1 OAI21X1_915 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5390_), .B(AES_CORE_DATAPATH__abc_15863_new_n5394_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5395_));
OAI21X1 OAI21X1_916 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5398_), .C(AES_CORE_DATAPATH__abc_15863_new_n5361_), .Y(AES_CORE_DATAPATH__0col_0__31_0__20_));
OAI21X1 OAI21X1_917 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3574_), .B(AES_CORE_DATAPATH__abc_15863_new_n5406_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5407_));
OAI21X1 OAI21X1_918 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5411_));
OAI21X1 OAI21X1_919 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__21_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5412_));
OAI21X1 OAI21X1_92 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2641_));
OAI21X1 OAI21X1_920 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5412_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5411_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5413_));
OAI21X1 OAI21X1_921 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5410_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5414_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5415_));
OAI21X1 OAI21X1_922 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5416_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5417_));
OAI21X1 OAI21X1_923 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5415_), .C(AES_CORE_DATAPATH__abc_15863_new_n5417_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5418_));
OAI21X1 OAI21X1_924 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5418_), .C(AES_CORE_DATAPATH__abc_15863_new_n5419_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5420_));
OAI21X1 OAI21X1_925 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5418_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5423_));
OAI21X1 OAI21X1_926 ( .A(\iv_out[21] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5423_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5424_));
OAI21X1 OAI21X1_927 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5408_), .B(AES_CORE_DATAPATH__abc_15863_new_n5422_), .C(AES_CORE_DATAPATH__abc_15863_new_n5424_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5425_));
OAI21X1 OAI21X1_928 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[21] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5427_));
OAI21X1 OAI21X1_929 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5430_));
OAI21X1 OAI21X1_93 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2641_), .C(AES_CORE_DATAPATH__abc_15863_new_n2642_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2643_));
OAI21X1 OAI21X1_930 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5430_), .B(AES_CORE_DATAPATH__abc_15863_new_n5429_), .C(AES_CORE_DATAPATH__abc_15863_new_n5431_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5432_));
OAI21X1 OAI21X1_931 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5428_), .B(AES_CORE_DATAPATH__abc_15863_new_n5432_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5433_));
OAI21X1 OAI21X1_932 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5437_), .C(AES_CORE_DATAPATH__abc_15863_new_n5400_), .Y(AES_CORE_DATAPATH__0col_0__31_0__21_));
OAI21X1 OAI21X1_933 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2973_), .B(AES_CORE_DATAPATH__abc_15863_new_n3591_), .C(AES_CORE_DATAPATH__abc_15863_new_n5443_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5444_));
OAI21X1 OAI21X1_934 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__22_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5448_));
OAI21X1 OAI21X1_935 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n5448_), .C(AES_CORE_DATAPATH__abc_15863_new_n5449_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5450_));
OAI21X1 OAI21X1_936 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5453_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5454_));
OAI21X1 OAI21X1_937 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4598_), .B(\iv_out[22] ), .C(AES_CORE_DATAPATH__abc_15863_new_n5454_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5455_));
OAI21X1 OAI21X1_938 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3596_), .B(AES_CORE_DATAPATH__abc_15863_new_n3593_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5457_));
OAI21X1 OAI21X1_939 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5453_), .C(AES_CORE_DATAPATH__abc_15863_new_n5460_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5461_));
OAI21X1 OAI21X1_94 ( .A(AES_CORE_DATAPATH_iv_2__22_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n2643_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2644_));
OAI21X1 OAI21X1_940 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[22] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5464_));
OAI21X1 OAI21X1_941 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5467_));
OAI21X1 OAI21X1_942 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5467_), .B(AES_CORE_DATAPATH__abc_15863_new_n5466_), .C(AES_CORE_DATAPATH__abc_15863_new_n5468_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5469_));
OAI21X1 OAI21X1_943 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5465_), .B(AES_CORE_DATAPATH__abc_15863_new_n5469_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5470_));
OAI21X1 OAI21X1_944 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5473_), .C(AES_CORE_DATAPATH__abc_15863_new_n5439_), .Y(AES_CORE_DATAPATH__0col_0__31_0__22_));
OAI21X1 OAI21X1_945 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3618_), .B(AES_CORE_DATAPATH__abc_15863_new_n3615_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5479_));
OAI21X1 OAI21X1_946 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5483_));
OAI21X1 OAI21X1_947 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5484_));
OAI21X1 OAI21X1_948 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5484_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5483_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5485_));
OAI21X1 OAI21X1_949 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5482_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5486_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5487_));
OAI21X1 OAI21X1_95 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__23_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2647_));
OAI21X1 OAI21X1_950 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5488_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5489_));
OAI21X1 OAI21X1_951 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5487_), .C(AES_CORE_DATAPATH__abc_15863_new_n5489_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5490_));
OAI21X1 OAI21X1_952 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5490_), .C(AES_CORE_DATAPATH__abc_15863_new_n5491_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5492_));
OAI21X1 OAI21X1_953 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5490_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5499_));
OAI21X1 OAI21X1_954 ( .A(\iv_out[23] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5499_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5500_));
OAI21X1 OAI21X1_955 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5480_), .B(AES_CORE_DATAPATH__abc_15863_new_n5498_), .C(AES_CORE_DATAPATH__abc_15863_new_n5500_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5501_));
OAI21X1 OAI21X1_956 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[23] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5503_));
OAI21X1 OAI21X1_957 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5506_));
OAI21X1 OAI21X1_958 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5506_), .B(AES_CORE_DATAPATH__abc_15863_new_n5505_), .C(AES_CORE_DATAPATH__abc_15863_new_n5507_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5508_));
OAI21X1 OAI21X1_959 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5504_), .B(AES_CORE_DATAPATH__abc_15863_new_n5508_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5509_));
OAI21X1 OAI21X1_96 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2647_), .C(AES_CORE_DATAPATH__abc_15863_new_n2648_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2649_));
OAI21X1 OAI21X1_960 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5512_), .C(AES_CORE_DATAPATH__abc_15863_new_n5475_), .Y(AES_CORE_DATAPATH__0col_0__31_0__23_));
OAI21X1 OAI21X1_961 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2997_), .B(AES_CORE_DATAPATH__abc_15863_new_n3635_), .C(AES_CORE_DATAPATH__abc_15863_new_n5518_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5519_));
OAI21X1 OAI21X1_962 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5524_));
OAI21X1 OAI21X1_963 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5525_));
OAI21X1 OAI21X1_964 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5525_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5524_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5526_));
OAI21X1 OAI21X1_965 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5523_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5527_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5528_));
OAI21X1 OAI21X1_966 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5529_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5530_));
OAI21X1 OAI21X1_967 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5528_), .C(AES_CORE_DATAPATH__abc_15863_new_n5530_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5531_));
OAI21X1 OAI21X1_968 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5531_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5532_));
OAI21X1 OAI21X1_969 ( .A(\iv_out[24] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5532_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5533_));
OAI21X1 OAI21X1_97 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2646_), .B(AES_CORE_DATAPATH__abc_15863_new_n2463_), .C(AES_CORE_DATAPATH__abc_15863_new_n2652_), .Y(\iv_out[23] ));
OAI21X1 OAI21X1_970 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3640_), .B(AES_CORE_DATAPATH__abc_15863_new_n3637_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5535_));
OAI21X1 OAI21X1_971 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5531_), .C(AES_CORE_DATAPATH__abc_15863_new_n5538_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5539_));
OAI21X1 OAI21X1_972 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[24] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5542_));
OAI21X1 OAI21X1_973 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5545_));
OAI21X1 OAI21X1_974 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5545_), .B(AES_CORE_DATAPATH__abc_15863_new_n5544_), .C(AES_CORE_DATAPATH__abc_15863_new_n5546_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5547_));
OAI21X1 OAI21X1_975 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5543_), .B(AES_CORE_DATAPATH__abc_15863_new_n5547_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5548_));
OAI21X1 OAI21X1_976 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5551_), .C(AES_CORE_DATAPATH__abc_15863_new_n5514_), .Y(AES_CORE_DATAPATH__0col_0__31_0__24_));
OAI21X1 OAI21X1_977 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3662_), .B(AES_CORE_DATAPATH__abc_15863_new_n5559_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5560_));
OAI21X1 OAI21X1_978 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5564_));
OAI21X1 OAI21X1_979 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__25_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5565_));
OAI21X1 OAI21X1_98 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_iv_0__24_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2655_));
OAI21X1 OAI21X1_980 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5565_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5564_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5566_));
OAI21X1 OAI21X1_981 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5563_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5567_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5568_));
OAI21X1 OAI21X1_982 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5569_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5570_));
OAI21X1 OAI21X1_983 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5568_), .C(AES_CORE_DATAPATH__abc_15863_new_n5570_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5571_));
OAI21X1 OAI21X1_984 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4597_), .B(AES_CORE_DATAPATH__abc_15863_new_n5571_), .C(AES_CORE_DATAPATH__abc_15863_new_n5572_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5573_));
OAI21X1 OAI21X1_985 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH__abc_15863_new_n4596_), .C(AES_CORE_DATAPATH__abc_15863_new_n5571_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5576_));
OAI21X1 OAI21X1_986 ( .A(\iv_out[25] ), .B(AES_CORE_DATAPATH__abc_15863_new_n4598_), .C(AES_CORE_DATAPATH__abc_15863_new_n5576_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5577_));
OAI21X1 OAI21X1_987 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5561_), .B(AES_CORE_DATAPATH__abc_15863_new_n5575_), .C(AES_CORE_DATAPATH__abc_15863_new_n5577_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5578_));
OAI21X1 OAI21X1_988 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(\iv_out[25] ), .C(AES_CORE_DATAPATH__abc_15863_new_n4618_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5580_));
OAI21X1 OAI21X1_989 ( .A(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .B(AES_CORE_DATAPATH__abc_15863_new_n4624_), .C(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_15863_new_n5583_));
OAI21X1 OAI21X1_99 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2475_), .B(AES_CORE_DATAPATH__abc_15863_new_n2655_), .C(AES_CORE_DATAPATH__abc_15863_new_n2656_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2657_));
OAI21X1 OAI21X1_990 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5583_), .B(AES_CORE_DATAPATH__abc_15863_new_n5582_), .C(AES_CORE_DATAPATH__abc_15863_new_n5584_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5585_));
OAI21X1 OAI21X1_991 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5581_), .B(AES_CORE_DATAPATH__abc_15863_new_n5585_), .C(AES_CORE_DATAPATH__abc_15863_new_n4588_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5586_));
OAI21X1 OAI21X1_992 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4571_), .B(AES_CORE_DATAPATH__abc_15863_new_n5590_), .C(AES_CORE_DATAPATH__abc_15863_new_n5553_), .Y(AES_CORE_DATAPATH__0col_0__31_0__25_));
OAI21X1 OAI21X1_993 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3684_), .B(AES_CORE_DATAPATH__abc_15863_new_n5598_), .C(AES_CORE_DATAPATH__abc_15863_new_n4593_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5599_));
OAI21X1 OAI21X1_994 ( .A(\iv_sel_rd[1] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2473_), .C(AES_CORE_DATAPATH_bkp_1__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5603_));
OAI21X1 OAI21X1_995 ( .A(\iv_sel_rd[0] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2478_), .C(AES_CORE_DATAPATH_bkp_0__26_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5604_));
OAI21X1 OAI21X1_996 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5604_), .B(AES_CORE_DATAPATH__abc_15863_new_n2475_), .C(AES_CORE_DATAPATH__abc_15863_new_n5603_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5605_));
OAI21X1 OAI21X1_997 ( .A(AES_CORE_DATAPATH__abc_15863_new_n5602_), .B(AES_CORE_DATAPATH__abc_15863_new_n2467_), .C(AES_CORE_DATAPATH__abc_15863_new_n5606_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5607_));
OAI21X1 OAI21X1_998 ( .A(\iv_sel_rd[3] ), .B(AES_CORE_DATAPATH__abc_15863_new_n2462_), .C(AES_CORE_DATAPATH__abc_15863_new_n5608_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5609_));
OAI21X1 OAI21X1_999 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2482_), .B(AES_CORE_DATAPATH__abc_15863_new_n5607_), .C(AES_CORE_DATAPATH__abc_15863_new_n5609_), .Y(AES_CORE_DATAPATH__abc_15863_new_n5610_));
OAI22X1 OAI22X1_1 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n97_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n105_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n102_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_8_));
OAI22X1 OAI22X1_10 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3160_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3161_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3162_));
OAI22X1 OAI22X1_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3249_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3250_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3251_));
OAI22X1 OAI22X1_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3293_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3294_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3295_));
OAI22X1 OAI22X1_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3337_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3338_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3339_));
OAI22X1 OAI22X1_14 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3381_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3382_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3383_));
OAI22X1 OAI22X1_15 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3425_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3426_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3427_));
OAI22X1 OAI22X1_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3469_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3470_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3471_));
OAI22X1 OAI22X1_17 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3491_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3492_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3493_));
OAI22X1 OAI22X1_18 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3513_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3514_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3515_));
OAI22X1 OAI22X1_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3557_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3558_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3559_));
OAI22X1 OAI22X1_2 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n108_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_1_));
OAI22X1 OAI22X1_20 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3601_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3602_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3603_));
OAI22X1 OAI22X1_21 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3645_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3646_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3647_));
OAI22X1 OAI22X1_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3667_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3668_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3669_));
OAI22X1 OAI22X1_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3711_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3712_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3713_));
OAI22X1 OAI22X1_24 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3777_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3778_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3779_));
OAI22X1 OAI22X1_25 ( .A(\bus_in[0] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .C(AES_CORE_DATAPATH__abc_15863_new_n2457_), .D(AES_CORE_DATAPATH__abc_15863_new_n6982_), .Y(AES_CORE_DATAPATH__abc_15863_new_n6983_));
OAI22X1 OAI22X1_26 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n425_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n439_), .D(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n441_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n442_));
OAI22X1 OAI22X1_27 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n459_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n440_), .C(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n416_), .D(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n415_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n460_));
OAI22X1 OAI22X1_28 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n165_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n168_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n202_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n204_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n205_));
OAI22X1 OAI22X1_29 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n188_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n189_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n206_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n207_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n208_));
OAI22X1 OAI22X1_3 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n117_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n108_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_6_));
OAI22X1 OAI22X1_30 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n165_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n168_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n206_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n207_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n210_));
OAI22X1 OAI22X1_31 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n188_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n189_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n202_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n204_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n211_));
OAI22X1 OAI22X1_32 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n213_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n215_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n115_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n117_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n216_));
OAI22X1 OAI22X1_33 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n248_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n250_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n251_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n252_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n253_));
OAI22X1 OAI22X1_34 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n139_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n140_), .C(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n254_), .D(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n256_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n257_));
OAI22X1 OAI22X1_35 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n308_));
OAI22X1 OAI22X1_36 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n313_));
OAI22X1 OAI22X1_37 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n206_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n326_));
OAI22X1 OAI22X1_38 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n334_));
OAI22X1 OAI22X1_39 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n337_));
OAI22X1 OAI22X1_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n119_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n117_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_9_));
OAI22X1 OAI22X1_40 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n341_));
OAI22X1 OAI22X1_41 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n342_));
OAI22X1 OAI22X1_42 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n354_));
OAI22X1 OAI22X1_43 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n355_));
OAI22X1 OAI22X1_44 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n380_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n372_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n381_));
OAI22X1 OAI22X1_45 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n81_), .D(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n397_));
OAI22X1 OAI22X1_46 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n308_));
OAI22X1 OAI22X1_47 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n313_));
OAI22X1 OAI22X1_48 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n206_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n326_));
OAI22X1 OAI22X1_49 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n334_));
OAI22X1 OAI22X1_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n102_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n122_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_12_));
OAI22X1 OAI22X1_50 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n337_));
OAI22X1 OAI22X1_51 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n341_));
OAI22X1 OAI22X1_52 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n342_));
OAI22X1 OAI22X1_53 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n354_));
OAI22X1 OAI22X1_54 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n355_));
OAI22X1 OAI22X1_55 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n380_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n372_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n381_));
OAI22X1 OAI22X1_56 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n81_), .D(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n397_));
OAI22X1 OAI22X1_57 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n308_));
OAI22X1 OAI22X1_58 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n313_));
OAI22X1 OAI22X1_59 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n206_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n326_));
OAI22X1 OAI22X1_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n97_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n89_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n139_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_13_));
OAI22X1 OAI22X1_60 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n334_));
OAI22X1 OAI22X1_61 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n337_));
OAI22X1 OAI22X1_62 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n341_));
OAI22X1 OAI22X1_63 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n342_));
OAI22X1 OAI22X1_64 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n354_));
OAI22X1 OAI22X1_65 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n355_));
OAI22X1 OAI22X1_66 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n380_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n372_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n381_));
OAI22X1 OAI22X1_67 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n81_), .D(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n397_));
OAI22X1 OAI22X1_68 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n308_));
OAI22X1 OAI22X1_69 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n313_));
OAI22X1 OAI22X1_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n119_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_14_));
OAI22X1 OAI22X1_70 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n172_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n206_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n204_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n326_));
OAI22X1 OAI22X1_71 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n334_));
OAI22X1 OAI22X1_72 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n337_));
OAI22X1 OAI22X1_73 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n302_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n341_));
OAI22X1 OAI22X1_74 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n312_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n342_));
OAI22X1 OAI22X1_75 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n289_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n292_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n330_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n333_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n354_));
OAI22X1 OAI22X1_76 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n309_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n310_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n335_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n336_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n355_));
OAI22X1 OAI22X1_77 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n380_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n372_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n381_));
OAI22X1 OAI22X1_78 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n66_), .C(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n81_), .D(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n78_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n397_));
OAI22X1 OAI22X1_8 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n162_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n190_), .C(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_), .D(AES_CORE_CONTROL_UNIT__abc_15585_new_n183_), .Y(AES_CORE_CONTROL_UNIT_col_sel_1_));
OAI22X1 OAI22X1_9 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3115_), .B(AES_CORE_DATAPATH__abc_15863_new_n3089_), .C(AES_CORE_DATAPATH__abc_15863_new_n3116_), .D(AES_CORE_DATAPATH__abc_15863_new_n3117_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3118_));
OR2X2 OR2X2_1 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .B(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n91_));
OR2X2 OR2X2_10 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3207_), .B(AES_CORE_DATAPATH__abc_15863_new_n3211_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_));
OR2X2 OR2X2_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3229_), .B(AES_CORE_DATAPATH__abc_15863_new_n3233_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_));
OR2X2 OR2X2_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3251_), .B(AES_CORE_DATAPATH__abc_15863_new_n3255_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_));
OR2X2 OR2X2_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3273_), .B(AES_CORE_DATAPATH__abc_15863_new_n3277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_));
OR2X2 OR2X2_14 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3295_), .B(AES_CORE_DATAPATH__abc_15863_new_n3299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_));
OR2X2 OR2X2_15 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3317_), .B(AES_CORE_DATAPATH__abc_15863_new_n3321_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_));
OR2X2 OR2X2_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3339_), .B(AES_CORE_DATAPATH__abc_15863_new_n3343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_));
OR2X2 OR2X2_17 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3361_), .B(AES_CORE_DATAPATH__abc_15863_new_n3365_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_));
OR2X2 OR2X2_18 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3383_), .B(AES_CORE_DATAPATH__abc_15863_new_n3387_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_));
OR2X2 OR2X2_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3405_), .B(AES_CORE_DATAPATH__abc_15863_new_n3409_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_));
OR2X2 OR2X2_2 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n133_), .Y(AES_CORE_CONTROL_UNIT_bypass_key_en));
OR2X2 OR2X2_20 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3427_), .B(AES_CORE_DATAPATH__abc_15863_new_n3431_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_));
OR2X2 OR2X2_21 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3449_), .B(AES_CORE_DATAPATH__abc_15863_new_n3453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_));
OR2X2 OR2X2_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3471_), .B(AES_CORE_DATAPATH__abc_15863_new_n3475_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_));
OR2X2 OR2X2_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3493_), .B(AES_CORE_DATAPATH__abc_15863_new_n3497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_));
OR2X2 OR2X2_24 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3515_), .B(AES_CORE_DATAPATH__abc_15863_new_n3519_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_));
OR2X2 OR2X2_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3537_), .B(AES_CORE_DATAPATH__abc_15863_new_n3541_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_));
OR2X2 OR2X2_26 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3559_), .B(AES_CORE_DATAPATH__abc_15863_new_n3563_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_));
OR2X2 OR2X2_27 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3581_), .B(AES_CORE_DATAPATH__abc_15863_new_n3585_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_));
OR2X2 OR2X2_28 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3603_), .B(AES_CORE_DATAPATH__abc_15863_new_n3607_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_));
OR2X2 OR2X2_29 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3625_), .B(AES_CORE_DATAPATH__abc_15863_new_n3629_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_));
OR2X2 OR2X2_3 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT_key_en_0_));
OR2X2 OR2X2_30 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3647_), .B(AES_CORE_DATAPATH__abc_15863_new_n3651_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_));
OR2X2 OR2X2_31 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3669_), .B(AES_CORE_DATAPATH__abc_15863_new_n3673_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_));
OR2X2 OR2X2_32 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3691_), .B(AES_CORE_DATAPATH__abc_15863_new_n3695_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_));
OR2X2 OR2X2_33 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3713_), .B(AES_CORE_DATAPATH__abc_15863_new_n3717_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_));
OR2X2 OR2X2_34 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3735_), .B(AES_CORE_DATAPATH__abc_15863_new_n3739_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_));
OR2X2 OR2X2_35 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3757_), .B(AES_CORE_DATAPATH__abc_15863_new_n3761_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_));
OR2X2 OR2X2_36 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3779_), .B(AES_CORE_DATAPATH__abc_15863_new_n3783_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_));
OR2X2 OR2X2_37 ( .A(AES_CORE_DATAPATH__abc_15863_new_n4032_), .B(start), .Y(AES_CORE_DATAPATH__abc_15863_new_n4033_));
OR2X2 OR2X2_38 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7073_), .B(AES_CORE_DATAPATH__abc_15863_new_n7072_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7074_));
OR2X2 OR2X2_39 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7079_), .B(AES_CORE_DATAPATH__abc_15863_new_n7078_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7080_));
OR2X2 OR2X2_4 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_15863_new_n2710_));
OR2X2 OR2X2_40 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7085_), .B(AES_CORE_DATAPATH__abc_15863_new_n7086_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7087_));
OR2X2 OR2X2_41 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3090_), .B(AES_CORE_DATAPATH__abc_15863_new_n3096_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_));
OR2X2 OR2X2_42 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec));
OR2X2 OR2X2_43 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n101_));
OR2X2 OR2X2_44 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n135_));
OR2X2 OR2X2_45 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n238_));
OR2X2 OR2X2_46 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n51_));
OR2X2 OR2X2_47 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n103_));
OR2X2 OR2X2_48 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n195_));
OR2X2 OR2X2_49 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n232_));
OR2X2 OR2X2_5 ( .A(AES_CORE_DATAPATH_col_sel_host_0_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_0_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3082_));
OR2X2 OR2X2_50 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n300_));
OR2X2 OR2X2_51 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n476_));
OR2X2 OR2X2_52 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n51_));
OR2X2 OR2X2_53 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n103_));
OR2X2 OR2X2_54 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n195_));
OR2X2 OR2X2_55 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n232_));
OR2X2 OR2X2_56 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n300_));
OR2X2 OR2X2_57 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n476_));
OR2X2 OR2X2_58 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n51_));
OR2X2 OR2X2_59 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n103_));
OR2X2 OR2X2_6 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3118_), .B(AES_CORE_DATAPATH__abc_15863_new_n3122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_));
OR2X2 OR2X2_60 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n195_));
OR2X2 OR2X2_61 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n232_));
OR2X2 OR2X2_62 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n300_));
OR2X2 OR2X2_63 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n476_));
OR2X2 OR2X2_64 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n51_));
OR2X2 OR2X2_65 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n103_));
OR2X2 OR2X2_66 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n152_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n195_));
OR2X2 OR2X2_67 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n232_));
OR2X2 OR2X2_68 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n216_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n300_));
OR2X2 OR2X2_69 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n476_));
OR2X2 OR2X2_7 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3140_), .B(AES_CORE_DATAPATH__abc_15863_new_n3144_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_));
OR2X2 OR2X2_8 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3162_), .B(AES_CORE_DATAPATH__abc_15863_new_n3166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_));
OR2X2 OR2X2_9 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3185_), .B(AES_CORE_DATAPATH__abc_15863_new_n3189_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_));
XNOR2X1 XNOR2X1_1 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n157_), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n158_));
XNOR2X1 XNOR2X1_10 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n348_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n349_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_));
XNOR2X1 XNOR2X1_100 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n409_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n407_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_));
XNOR2X1 XNOR2X1_101 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n420_));
XNOR2X1 XNOR2X1_102 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n420_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n419_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n421_));
XNOR2X1 XNOR2X1_103 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n431_));
XNOR2X1 XNOR2X1_104 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_));
XNOR2X1 XNOR2X1_105 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n433_));
XNOR2X1 XNOR2X1_106 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n433_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n431_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_));
XNOR2X1 XNOR2X1_107 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n350_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n110_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n435_));
XNOR2X1 XNOR2X1_108 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n435_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_));
XNOR2X1 XNOR2X1_109 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n437_));
XNOR2X1 XNOR2X1_11 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n351_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n352_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_));
XNOR2X1 XNOR2X1_110 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n97_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n438_));
XNOR2X1 XNOR2X1_111 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n438_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n437_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_));
XNOR2X1 XNOR2X1_112 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n120_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_));
XNOR2X1 XNOR2X1_113 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n371_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n441_));
XNOR2X1 XNOR2X1_114 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n442_));
XNOR2X1 XNOR2X1_115 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n437_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n442_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n443_));
XNOR2X1 XNOR2X1_116 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n443_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n441_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_));
XNOR2X1 XNOR2X1_117 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n449_));
XNOR2X1 XNOR2X1_118 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n449_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n124_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_));
XNOR2X1 XNOR2X1_119 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n194_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_));
XNOR2X1 XNOR2X1_12 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n354_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n355_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_));
XNOR2X1 XNOR2X1_120 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n452_));
XNOR2X1 XNOR2X1_121 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n437_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n452_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n453_));
XNOR2X1 XNOR2X1_122 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n198_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n454_));
XNOR2X1 XNOR2X1_123 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n453_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n454_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_));
XNOR2X1 XNOR2X1_124 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n460_));
XNOR2X1 XNOR2X1_125 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n437_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n460_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n461_));
XNOR2X1 XNOR2X1_126 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n407_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n346_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n462_));
XNOR2X1 XNOR2X1_127 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n461_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n462_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_));
XNOR2X1 XNOR2X1_128 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n235_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n107_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n468_));
XNOR2X1 XNOR2X1_129 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n468_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n110_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n469_));
XNOR2X1 XNOR2X1_13 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n357_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n358_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_));
XNOR2X1 XNOR2X1_130 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n474_));
XNOR2X1 XNOR2X1_131 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n474_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n475_));
XNOR2X1 XNOR2X1_132 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n475_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n342_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n476_));
XNOR2X1 XNOR2X1_133 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n481_));
XNOR2X1 XNOR2X1_134 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n482_));
XNOR2X1 XNOR2X1_135 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n482_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n481_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_));
XNOR2X1 XNOR2X1_136 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n351_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_));
XNOR2X1 XNOR2X1_137 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n442_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n485_));
XNOR2X1 XNOR2X1_138 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n485_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_));
XNOR2X1 XNOR2X1_139 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n488_));
XNOR2X1 XNOR2X1_14 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n360_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n361_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_));
XNOR2X1 XNOR2X1_140 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n488_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n489_));
XNOR2X1 XNOR2X1_141 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n371_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n217_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n490_));
XNOR2X1 XNOR2X1_142 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n360_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n496_));
XNOR2X1 XNOR2X1_143 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n496_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n452_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_));
XNOR2X1 XNOR2X1_144 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n378_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_));
XNOR2X1 XNOR2X1_145 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n499_));
XNOR2X1 XNOR2X1_146 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n499_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n500_));
XNOR2X1 XNOR2X1_147 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n294_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n501_));
XNOR2X1 XNOR2X1_148 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n500_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n501_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n502_));
XNOR2X1 XNOR2X1_149 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n345_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n507_));
XNOR2X1 XNOR2X1_15 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n363_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n364_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_));
XNOR2X1 XNOR2X1_150 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n380_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n432_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n508_));
XNOR2X1 XNOR2X1_151 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n508_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n507_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n510_));
XNOR2X1 XNOR2X1_152 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n104_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n515_));
XNOR2X1 XNOR2X1_153 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n515_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n514_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n516_));
XNOR2X1 XNOR2X1_154 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n408_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n170_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n521_));
XNOR2X1 XNOR2X1_155 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n521_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n144_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_));
XNOR2X1 XNOR2X1_156 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n128_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n527_));
XNOR2X1 XNOR2X1_157 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n527_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n324_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_));
XNOR2X1 XNOR2X1_158 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n435_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_));
XNOR2X1 XNOR2X1_159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n54_));
XNOR2X1 XNOR2X1_16 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n366_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n367_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_));
XNOR2X1 XNOR2X1_160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n55_));
XNOR2X1 XNOR2X1_161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n79_));
XNOR2X1 XNOR2X1_162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n97_));
XNOR2X1 XNOR2X1_163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n100_));
XNOR2X1 XNOR2X1_164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n121_));
XNOR2X1 XNOR2X1_165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n127_));
XNOR2X1 XNOR2X1_166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n129_));
XNOR2X1 XNOR2X1_167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n131_));
XNOR2X1 XNOR2X1_168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n196_));
XNOR2X1 XNOR2X1_169 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n224_));
XNOR2X1 XNOR2X1_17 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n369_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n370_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_));
XNOR2X1 XNOR2X1_170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n278_));
XNOR2X1 XNOR2X1_171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n282_));
XNOR2X1 XNOR2X1_172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n301_));
XNOR2X1 XNOR2X1_173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n306_));
XNOR2X1 XNOR2X1_174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n347_));
XNOR2X1 XNOR2X1_175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n364_));
XNOR2X1 XNOR2X1_176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n353_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_));
XNOR2X1 XNOR2X1_177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n369_));
XNOR2X1 XNOR2X1_178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n413_));
XNOR2X1 XNOR2X1_179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n425_));
XNOR2X1 XNOR2X1_18 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n372_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n373_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_));
XNOR2X1 XNOR2X1_180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n407_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n437_));
XNOR2X1 XNOR2X1_181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n54_));
XNOR2X1 XNOR2X1_182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n55_));
XNOR2X1 XNOR2X1_183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n79_));
XNOR2X1 XNOR2X1_184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n97_));
XNOR2X1 XNOR2X1_185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n100_));
XNOR2X1 XNOR2X1_186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n121_));
XNOR2X1 XNOR2X1_187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n127_));
XNOR2X1 XNOR2X1_188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n129_));
XNOR2X1 XNOR2X1_189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n131_));
XNOR2X1 XNOR2X1_19 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n376_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_));
XNOR2X1 XNOR2X1_190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n196_));
XNOR2X1 XNOR2X1_191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n224_));
XNOR2X1 XNOR2X1_192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n278_));
XNOR2X1 XNOR2X1_193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n282_));
XNOR2X1 XNOR2X1_194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n301_));
XNOR2X1 XNOR2X1_195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n306_));
XNOR2X1 XNOR2X1_196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n347_));
XNOR2X1 XNOR2X1_197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n364_));
XNOR2X1 XNOR2X1_198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n353_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_));
XNOR2X1 XNOR2X1_199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n369_));
XNOR2X1 XNOR2X1_2 ( .A(AES_CORE_DATAPATH__abc_15863_new_n7015_), .B(AES_CORE_DATAPATH__abc_15863_new_n2520_), .Y(AES_CORE_DATAPATH__abc_15863_new_n7023_));
XNOR2X1 XNOR2X1_20 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n378_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n379_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_));
XNOR2X1 XNOR2X1_200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n413_));
XNOR2X1 XNOR2X1_201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n425_));
XNOR2X1 XNOR2X1_202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n407_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n437_));
XNOR2X1 XNOR2X1_203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n54_));
XNOR2X1 XNOR2X1_204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n55_));
XNOR2X1 XNOR2X1_205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n79_));
XNOR2X1 XNOR2X1_206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n97_));
XNOR2X1 XNOR2X1_207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n100_));
XNOR2X1 XNOR2X1_208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n121_));
XNOR2X1 XNOR2X1_209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n127_));
XNOR2X1 XNOR2X1_21 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n381_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n382_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_));
XNOR2X1 XNOR2X1_210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n129_));
XNOR2X1 XNOR2X1_211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n131_));
XNOR2X1 XNOR2X1_212 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n196_));
XNOR2X1 XNOR2X1_213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n224_));
XNOR2X1 XNOR2X1_214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n278_));
XNOR2X1 XNOR2X1_215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n282_));
XNOR2X1 XNOR2X1_216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n301_));
XNOR2X1 XNOR2X1_217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n306_));
XNOR2X1 XNOR2X1_218 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n347_));
XNOR2X1 XNOR2X1_219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n364_));
XNOR2X1 XNOR2X1_22 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n384_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n385_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_));
XNOR2X1 XNOR2X1_220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n353_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_));
XNOR2X1 XNOR2X1_221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n369_));
XNOR2X1 XNOR2X1_222 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n413_));
XNOR2X1 XNOR2X1_223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n425_));
XNOR2X1 XNOR2X1_224 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n407_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n437_));
XNOR2X1 XNOR2X1_225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n54_));
XNOR2X1 XNOR2X1_226 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n55_));
XNOR2X1 XNOR2X1_227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n79_));
XNOR2X1 XNOR2X1_228 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n97_));
XNOR2X1 XNOR2X1_229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n99_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n100_));
XNOR2X1 XNOR2X1_23 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n387_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n388_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_));
XNOR2X1 XNOR2X1_230 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n121_));
XNOR2X1 XNOR2X1_231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n127_));
XNOR2X1 XNOR2X1_232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n129_));
XNOR2X1 XNOR2X1_233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n131_));
XNOR2X1 XNOR2X1_234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n196_));
XNOR2X1 XNOR2X1_235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n224_));
XNOR2X1 XNOR2X1_236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n278_));
XNOR2X1 XNOR2X1_237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n282_));
XNOR2X1 XNOR2X1_238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n220_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n301_));
XNOR2X1 XNOR2X1_239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n219_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n306_));
XNOR2X1 XNOR2X1_24 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n390_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n391_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_));
XNOR2X1 XNOR2X1_240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n347_));
XNOR2X1 XNOR2X1_241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n364_));
XNOR2X1 XNOR2X1_242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n353_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_));
XNOR2X1 XNOR2X1_243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n223_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n369_));
XNOR2X1 XNOR2X1_244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n413_));
XNOR2X1 XNOR2X1_245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n425_));
XNOR2X1 XNOR2X1_246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n407_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n437_));
XNOR2X1 XNOR2X1_25 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n393_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n394_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_));
XNOR2X1 XNOR2X1_26 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n396_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n397_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_));
XNOR2X1 XNOR2X1_27 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n409_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n399_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_));
XNOR2X1 XNOR2X1_28 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n429_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n411_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_));
XNOR2X1 XNOR2X1_29 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n479_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n481_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n490_));
XNOR2X1 XNOR2X1_3 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n327_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n328_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_));
XNOR2X1 XNOR2X1_30 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n516_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n508_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_));
XNOR2X1 XNOR2X1_31 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n525_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n518_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_));
XNOR2X1 XNOR2X1_32 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n680_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_));
XNOR2X1 XNOR2X1_33 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n692_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_));
XNOR2X1 XNOR2X1_34 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n694_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_));
XNOR2X1 XNOR2X1_35 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n97_));
XNOR2X1 XNOR2X1_36 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_));
XNOR2X1 XNOR2X1_37 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n99_));
XNOR2X1 XNOR2X1_38 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n99_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n97_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_));
XNOR2X1 XNOR2X1_39 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n104_));
XNOR2X1 XNOR2X1_4 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n330_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n331_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_));
XNOR2X1 XNOR2X1_40 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n110_));
XNOR2X1 XNOR2X1_41 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n120_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_));
XNOR2X1 XNOR2X1_42 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n122_));
XNOR2X1 XNOR2X1_43 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n122_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n123_));
XNOR2X1 XNOR2X1_44 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n124_));
XNOR2X1 XNOR2X1_45 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n124_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n125_));
XNOR2X1 XNOR2X1_46 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n123_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n125_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_));
XNOR2X1 XNOR2X1_47 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n103_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n141_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n142_));
XNOR2X1 XNOR2X1_48 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n144_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n141_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n145_));
XNOR2X1 XNOR2X1_49 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n159_));
XNOR2X1 XNOR2X1_5 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n333_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n334_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_));
XNOR2X1 XNOR2X1_50 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n159_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n160_));
XNOR2X1 XNOR2X1_51 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_));
XNOR2X1 XNOR2X1_52 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n160_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n161_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_));
XNOR2X1 XNOR2X1_53 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n167_));
XNOR2X1 XNOR2X1_54 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n194_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_));
XNOR2X1 XNOR2X1_55 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n196_));
XNOR2X1 XNOR2X1_56 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n196_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n197_));
XNOR2X1 XNOR2X1_57 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n198_));
XNOR2X1 XNOR2X1_58 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n198_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n199_));
XNOR2X1 XNOR2X1_59 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n197_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_));
XNOR2X1 XNOR2X1_6 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n336_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n337_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_));
XNOR2X1 XNOR2X1_60 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n233_));
XNOR2X1 XNOR2X1_61 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n98_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n233_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n234_));
XNOR2X1 XNOR2X1_62 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n235_));
XNOR2X1 XNOR2X1_63 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n235_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n236_));
XNOR2X1 XNOR2X1_64 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n234_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n236_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_));
XNOR2X1 XNOR2X1_65 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n110_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n290_));
XNOR2X1 XNOR2X1_66 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n290_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n291_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n292_));
XNOR2X1 XNOR2X1_67 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n322_));
XNOR2X1 XNOR2X1_68 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n322_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n323_));
XNOR2X1 XNOR2X1_69 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_));
XNOR2X1 XNOR2X1_7 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n339_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n340_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_));
XNOR2X1 XNOR2X1_70 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n198_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n328_));
XNOR2X1 XNOR2X1_71 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n198_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n330_));
XNOR2X1 XNOR2X1_72 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n342_));
XNOR2X1 XNOR2X1_73 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n342_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n343_));
XNOR2X1 XNOR2X1_74 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n343_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n181_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_));
XNOR2X1 XNOR2X1_75 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n349_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n350_));
XNOR2X1 XNOR2X1_76 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n350_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n104_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n351_));
XNOR2X1 XNOR2X1_77 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n351_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_));
XNOR2X1 XNOR2X1_78 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_));
XNOR2X1 XNOR2X1_79 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n167_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n354_));
XNOR2X1 XNOR2X1_8 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n342_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n343_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_));
XNOR2X1 XNOR2X1_80 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n354_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_));
XNOR2X1 XNOR2X1_81 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n118_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n174_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n356_));
XNOR2X1 XNOR2X1_82 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n358_));
XNOR2X1 XNOR2X1_83 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n358_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n359_));
XNOR2X1 XNOR2X1_84 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n360_));
XNOR2X1 XNOR2X1_85 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n360_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n219_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n361_));
XNOR2X1 XNOR2X1_86 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n371_));
XNOR2X1 XNOR2X1_87 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n240_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n372_));
XNOR2X1 XNOR2X1_88 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n372_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n371_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_));
XNOR2X1 XNOR2X1_89 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n378_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_));
XNOR2X1 XNOR2X1_9 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n345_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n346_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_));
XNOR2X1 XNOR2X1_90 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n380_));
XNOR2X1 XNOR2X1_91 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n380_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n381_));
XNOR2X1 XNOR2X1_92 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n382_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n383_));
XNOR2X1 XNOR2X1_93 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n383_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n381_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n384_));
XNOR2X1 XNOR2X1_94 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n346_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n393_));
XNOR2X1 XNOR2X1_95 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n394_));
XNOR2X1 XNOR2X1_96 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n353_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n394_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n395_));
XNOR2X1 XNOR2X1_97 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n395_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n393_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n397_));
XNOR2X1 XNOR2X1_98 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n408_));
XNOR2X1 XNOR2X1_99 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n408_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n107_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n409_));
XOR2X1 XOR2X1_1 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2740_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2741_));
XOR2X1 XOR2X1_10 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2870_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2871_));
XOR2X1 XOR2X1_100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_));
XOR2X1 XOR2X1_101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_));
XOR2X1 XOR2X1_102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_));
XOR2X1 XOR2X1_103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_));
XOR2X1 XOR2X1_104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_));
XOR2X1 XOR2X1_105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_));
XOR2X1 XOR2X1_106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_));
XOR2X1 XOR2X1_107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_));
XOR2X1 XOR2X1_108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_));
XOR2X1 XOR2X1_109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_));
XOR2X1 XOR2X1_11 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2880_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2881_));
XOR2X1 XOR2X1_110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_));
XOR2X1 XOR2X1_111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_));
XOR2X1 XOR2X1_112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_));
XOR2X1 XOR2X1_113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_));
XOR2X1 XOR2X1_114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_));
XOR2X1 XOR2X1_115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_));
XOR2X1 XOR2X1_116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n408_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_));
XOR2X1 XOR2X1_117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n468_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_));
XOR2X1 XOR2X1_118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n490_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_));
XOR2X1 XOR2X1_119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_));
XOR2X1 XOR2X1_12 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2890_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2891_));
XOR2X1 XOR2X1_120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_));
XOR2X1 XOR2X1_121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_));
XOR2X1 XOR2X1_122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_));
XOR2X1 XOR2X1_123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_));
XOR2X1 XOR2X1_124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_));
XOR2X1 XOR2X1_125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_));
XOR2X1 XOR2X1_126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_));
XOR2X1 XOR2X1_127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_));
XOR2X1 XOR2X1_128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_));
XOR2X1 XOR2X1_129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_));
XOR2X1 XOR2X1_13 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2900_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2901_));
XOR2X1 XOR2X1_130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_));
XOR2X1 XOR2X1_131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_));
XOR2X1 XOR2X1_132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_));
XOR2X1 XOR2X1_133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_));
XOR2X1 XOR2X1_134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_));
XOR2X1 XOR2X1_135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_));
XOR2X1 XOR2X1_136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_));
XOR2X1 XOR2X1_137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_));
XOR2X1 XOR2X1_138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_));
XOR2X1 XOR2X1_139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_));
XOR2X1 XOR2X1_14 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2911_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2912_));
XOR2X1 XOR2X1_140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_));
XOR2X1 XOR2X1_141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_));
XOR2X1 XOR2X1_142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_));
XOR2X1 XOR2X1_143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_));
XOR2X1 XOR2X1_144 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_));
XOR2X1 XOR2X1_145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_));
XOR2X1 XOR2X1_146 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_));
XOR2X1 XOR2X1_147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_));
XOR2X1 XOR2X1_148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_));
XOR2X1 XOR2X1_149 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_));
XOR2X1 XOR2X1_15 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2920_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2921_));
XOR2X1 XOR2X1_150 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_));
XOR2X1 XOR2X1_151 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n105_));
XOR2X1 XOR2X1_152 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n123_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n125_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n127_));
XOR2X1 XOR2X1_153 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n164_));
XOR2X1 XOR2X1_154 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n175_));
XOR2X1 XOR2X1_155 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n197_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n201_));
XOR2X1 XOR2X1_156 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n203_));
XOR2X1 XOR2X1_157 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n234_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n236_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n285_));
XOR2X1 XOR2X1_158 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n291_));
XOR2X1 XOR2X1_159 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n294_));
XOR2X1 XOR2X1_16 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2930_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2931_));
XOR2X1 XOR2X1_160 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n324_));
XOR2X1 XOR2X1_161 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n323_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n324_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_));
XOR2X1 XOR2X1_162 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n356_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_));
XOR2X1 XOR2X1_163 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n359_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n361_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_));
XOR2X1 XOR2X1_164 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n382_));
XOR2X1 XOR2X1_165 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n395_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n393_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_));
XOR2X1 XOR2X1_166 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n407_));
XOR2X1 XOR2X1_167 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n419_));
XOR2X1 XOR2X1_168 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n443_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n441_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n445_));
XOR2X1 XOR2X1_169 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n453_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n454_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n456_));
XOR2X1 XOR2X1_17 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2940_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2941_));
XOR2X1 XOR2X1_170 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n461_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n462_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n465_));
XOR2X1 XOR2X1_171 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n356_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_));
XOR2X1 XOR2X1_172 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n489_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n490_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_));
XOR2X1 XOR2X1_173 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n508_), .B(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n507_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_));
XOR2X1 XOR2X1_174 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_22016_new_n514_));
XOR2X1 XOR2X1_175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n205_));
XOR2X1 XOR2X1_176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_));
XOR2X1 XOR2X1_177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n282_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_));
XOR2X1 XOR2X1_178 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_));
XOR2X1 XOR2X1_179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n412_));
XOR2X1 XOR2X1_18 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2963_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2964_));
XOR2X1 XOR2X1_180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_22451_new_n500_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_));
XOR2X1 XOR2X1_181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n205_));
XOR2X1 XOR2X1_182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_));
XOR2X1 XOR2X1_183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n282_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_));
XOR2X1 XOR2X1_184 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_));
XOR2X1 XOR2X1_185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n412_));
XOR2X1 XOR2X1_186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_22451_new_n500_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_));
XOR2X1 XOR2X1_187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n205_));
XOR2X1 XOR2X1_188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_));
XOR2X1 XOR2X1_189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n282_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_));
XOR2X1 XOR2X1_19 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2973_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2974_));
XOR2X1 XOR2X1_190 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_));
XOR2X1 XOR2X1_191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n412_));
XOR2X1 XOR2X1_192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_22451_new_n500_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_));
XOR2X1 XOR2X1_193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n205_));
XOR2X1 XOR2X1_194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_));
XOR2X1 XOR2X1_195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n282_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_));
XOR2X1 XOR2X1_196 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n224_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_));
XOR2X1 XOR2X1_197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n412_));
XOR2X1 XOR2X1_198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_22451_new_n500_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_));
XOR2X1 XOR2X1_2 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2764_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2765_));
XOR2X1 XOR2X1_20 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3009_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3010_));
XOR2X1 XOR2X1_21 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3019_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3020_));
XOR2X1 XOR2X1_22 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3029_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3030_));
XOR2X1 XOR2X1_23 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3040_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3041_));
XOR2X1 XOR2X1_24 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3050_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3051_));
XOR2X1 XOR2X1_25 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3060_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3061_));
XOR2X1 XOR2X1_26 ( .A(AES_CORE_DATAPATH__abc_15863_new_n3069_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_15863_new_n3070_));
XOR2X1 XOR2X1_27 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n327_));
XOR2X1 XOR2X1_28 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n330_));
XOR2X1 XOR2X1_29 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n333_));
XOR2X1 XOR2X1_3 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2774_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2775_));
XOR2X1 XOR2X1_30 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n336_));
XOR2X1 XOR2X1_31 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n339_));
XOR2X1 XOR2X1_32 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n342_));
XOR2X1 XOR2X1_33 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n345_));
XOR2X1 XOR2X1_34 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n348_));
XOR2X1 XOR2X1_35 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n351_));
XOR2X1 XOR2X1_36 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n354_));
XOR2X1 XOR2X1_37 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n357_));
XOR2X1 XOR2X1_38 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n360_));
XOR2X1 XOR2X1_39 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n363_));
XOR2X1 XOR2X1_4 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2784_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2785_));
XOR2X1 XOR2X1_40 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n366_));
XOR2X1 XOR2X1_41 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n369_));
XOR2X1 XOR2X1_42 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n372_));
XOR2X1 XOR2X1_43 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n375_));
XOR2X1 XOR2X1_44 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n378_));
XOR2X1 XOR2X1_45 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n381_));
XOR2X1 XOR2X1_46 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n384_));
XOR2X1 XOR2X1_47 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n387_));
XOR2X1 XOR2X1_48 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n390_));
XOR2X1 XOR2X1_49 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n393_));
XOR2X1 XOR2X1_5 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2794_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2795_));
XOR2X1 XOR2X1_50 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n396_));
XOR2X1 XOR2X1_51 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n399_));
XOR2X1 XOR2X1_52 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n407_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n408_));
XOR2X1 XOR2X1_53 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n411_));
XOR2X1 XOR2X1_54 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n431_));
XOR2X1 XOR2X1_55 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n456_));
XOR2X1 XOR2X1_56 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n475_));
XOR2X1 XOR2X1_57 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n493_));
XOR2X1 XOR2X1_58 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n508_));
XOR2X1 XOR2X1_59 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_21614_new_n518_));
XOR2X1 XOR2X1_6 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2804_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2805_));
XOR2X1 XOR2X1_60 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_));
XOR2X1 XOR2X1_61 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_));
XOR2X1 XOR2X1_62 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_));
XOR2X1 XOR2X1_63 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_));
XOR2X1 XOR2X1_64 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_));
XOR2X1 XOR2X1_65 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_));
XOR2X1 XOR2X1_66 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_));
XOR2X1 XOR2X1_67 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_));
XOR2X1 XOR2X1_68 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_));
XOR2X1 XOR2X1_69 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_));
XOR2X1 XOR2X1_7 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2840_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2841_));
XOR2X1 XOR2X1_70 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_));
XOR2X1 XOR2X1_71 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_));
XOR2X1 XOR2X1_72 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_));
XOR2X1 XOR2X1_73 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_));
XOR2X1 XOR2X1_74 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_));
XOR2X1 XOR2X1_75 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_));
XOR2X1 XOR2X1_76 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_));
XOR2X1 XOR2X1_77 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_));
XOR2X1 XOR2X1_78 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_));
XOR2X1 XOR2X1_79 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_));
XOR2X1 XOR2X1_8 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2851_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2852_));
XOR2X1 XOR2X1_80 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_));
XOR2X1 XOR2X1_81 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_));
XOR2X1 XOR2X1_82 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_));
XOR2X1 XOR2X1_83 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_));
XOR2X1 XOR2X1_84 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_));
XOR2X1 XOR2X1_85 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_));
XOR2X1 XOR2X1_86 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_));
XOR2X1 XOR2X1_87 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_));
XOR2X1 XOR2X1_88 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_));
XOR2X1 XOR2X1_89 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_));
XOR2X1 XOR2X1_9 ( .A(AES_CORE_DATAPATH__abc_15863_new_n2860_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_15863_new_n2861_));
XOR2X1 XOR2X1_90 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_));
XOR2X1 XOR2X1_91 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_));
XOR2X1 XOR2X1_92 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_));
XOR2X1 XOR2X1_93 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_));
XOR2X1 XOR2X1_94 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_));
XOR2X1 XOR2X1_95 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_));
XOR2X1 XOR2X1_96 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_));
XOR2X1 XOR2X1_97 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_));
XOR2X1 XOR2X1_98 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_));
XOR2X1 XOR2X1_99 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_));


endmodule