module aes_core(\bus_in[0] , \bus_in[1] , \bus_in[2] , \bus_in[3] , \bus_in[4] , \bus_in[5] , \bus_in[6] , \bus_in[7] , \bus_in[8] , \bus_in[9] , \bus_in[10] , \bus_in[11] , \bus_in[12] , \bus_in[13] , \bus_in[14] , \bus_in[15] , \bus_in[16] , \bus_in[17] , \bus_in[18] , \bus_in[19] , \bus_in[20] , \bus_in[21] , \bus_in[22] , \bus_in[23] , \bus_in[24] , \bus_in[25] , \bus_in[26] , \bus_in[27] , \bus_in[28] , \bus_in[29] , \bus_in[30] , \bus_in[31] , \iv_en[0] , \iv_en[1] , \iv_en[2] , \iv_en[3] , \iv_sel_rd[0] , \iv_sel_rd[1] , \iv_sel_rd[2] , \iv_sel_rd[3] , \key_en[0] , \key_en[1] , \key_en[2] , \key_en[3] , \key_sel_rd[0] , \key_sel_rd[1] , \data_type[0] , \data_type[1] , \addr[0] , \addr[1] , \op_mode[0] , \op_mode[1] , \aes_mode[0] , \aes_mode[1] , start, disable_core, write_en, read_en, first_block, rst_n, clk, \col_out[0] , \col_out[1] , \col_out[2] , \col_out[3] , \col_out[4] , \col_out[5] , \col_out[6] , \col_out[7] , \col_out[8] , \col_out[9] , \col_out[10] , \col_out[11] , \col_out[12] , \col_out[13] , \col_out[14] , \col_out[15] , \col_out[16] , \col_out[17] , \col_out[18] , \col_out[19] , \col_out[20] , \col_out[21] , \col_out[22] , \col_out[23] , \col_out[24] , \col_out[25] , \col_out[26] , \col_out[27] , \col_out[28] , \col_out[29] , \col_out[30] , \col_out[31] , \key_out[0] , \key_out[1] , \key_out[2] , \key_out[3] , \key_out[4] , \key_out[5] , \key_out[6] , \key_out[7] , \key_out[8] , \key_out[9] , \key_out[10] , \key_out[11] , \key_out[12] , \key_out[13] , \key_out[14] , \key_out[15] , \key_out[16] , \key_out[17] , \key_out[18] , \key_out[19] , \key_out[20] , \key_out[21] , \key_out[22] , \key_out[23] , \key_out[24] , \key_out[25] , \key_out[26] , \key_out[27] , \key_out[28] , \key_out[29] , \key_out[30] , \key_out[31] , \iv_out[0] , \iv_out[1] , \iv_out[2] , \iv_out[3] , \iv_out[4] , \iv_out[5] , \iv_out[6] , \iv_out[7] , \iv_out[8] , \iv_out[9] , \iv_out[10] , \iv_out[11] , \iv_out[12] , \iv_out[13] , \iv_out[14] , \iv_out[15] , \iv_out[16] , \iv_out[17] , \iv_out[18] , \iv_out[19] , \iv_out[20] , \iv_out[21] , \iv_out[22] , \iv_out[23] , \iv_out[24] , \iv_out[25] , \iv_out[26] , \iv_out[27] , \iv_out[28] , \iv_out[29] , \iv_out[30] , \iv_out[31] , end_aes);

wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__0_; 
wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__1_; 
wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__2_; 
wire AES_CORE_CONTROL_UNIT__0rd_count_3_0__3_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1817; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1856; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1897; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1928; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_0_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_10_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_12_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_13_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_14_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_1_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_2_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_4_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_5_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_6_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_8_; 
wire AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_9_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n100_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n101_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n102_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n103_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n104_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n105_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n106_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n107_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n108_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n109_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n111_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n112_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n113_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n114_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n115_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n117_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n118_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n119_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n121_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n122_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n123_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n125_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n126_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n127_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n128_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n129_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n130_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n131_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n132_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n133_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n135_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n136_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n138_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n139_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n141_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n142_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n143_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n144_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n145_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n146_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n147_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n149_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n150_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n152_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n153_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n154_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n156_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n157_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n159_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n160_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n161_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n163_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n164_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n167_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n168_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n169_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n170_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n172_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n173_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n174_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n175_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n177_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n178_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n179_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n180_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n182_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n183_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n184_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n185_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n187_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n188_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n189_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n191_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n192_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n193_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n197_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n198_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n199_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n200_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n201_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n202_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n203_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n205_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n206_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n208_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n209_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n211_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n212_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n213_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n214_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n215_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n216_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n217_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n218_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n219_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n220_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n221_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n222_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n223_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n224_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n225_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n227_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n228_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n229_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n230_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n231_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n232_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n233_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n234_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n238_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n239_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n240_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n243_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n244_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n245_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n247_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n248_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n249_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n251_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n252_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n253_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n257_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n258_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n73_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n74_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n76_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n77_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n78_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n79_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n80_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n81_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n82_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n83_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n84_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n86_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n87_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n88_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n90_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n91_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n92_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n93_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n94_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n95_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n96_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n97_; 
wire AES_CORE_CONTROL_UNIT__abc_15585_new_n99_; 
wire AES_CORE_CONTROL_UNIT_bypass_key_en; 
wire AES_CORE_CONTROL_UNIT_bypass_rk; 
wire AES_CORE_CONTROL_UNIT_col_en_0_; 
wire AES_CORE_CONTROL_UNIT_col_en_1_; 
wire AES_CORE_CONTROL_UNIT_col_en_2_; 
wire AES_CORE_CONTROL_UNIT_col_en_3_; 
wire AES_CORE_CONTROL_UNIT_col_sel_0_; 
wire AES_CORE_CONTROL_UNIT_col_sel_1_; 
wire AES_CORE_CONTROL_UNIT_encrypt_decrypt; 
wire AES_CORE_CONTROL_UNIT_iv_cnt_en; 
wire AES_CORE_CONTROL_UNIT_key_derivation_en; 
wire AES_CORE_CONTROL_UNIT_key_en_0_; 
wire AES_CORE_CONTROL_UNIT_key_en_1_; 
wire AES_CORE_CONTROL_UNIT_key_en_2_; 
wire AES_CORE_CONTROL_UNIT_key_en_3_; 
wire AES_CORE_CONTROL_UNIT_key_gen; 
wire AES_CORE_CONTROL_UNIT_key_out_sel_0_; 
wire AES_CORE_CONTROL_UNIT_key_out_sel_1_; 
wire AES_CORE_CONTROL_UNIT_key_sel; 
wire AES_CORE_CONTROL_UNIT_last_round; 
wire AES_CORE_CONTROL_UNIT_mode_cbc; 
wire AES_CORE_CONTROL_UNIT_mode_ctr; 
wire AES_CORE_CONTROL_UNIT_rd_count_0_; 
wire AES_CORE_CONTROL_UNIT_rd_count_1_; 
wire AES_CORE_CONTROL_UNIT_rd_count_2_; 
wire AES_CORE_CONTROL_UNIT_rd_count_3_; 
wire AES_CORE_CONTROL_UNIT_rk_sel_0_; 
wire AES_CORE_CONTROL_UNIT_rk_sel_1_; 
wire AES_CORE_CONTROL_UNIT_sbox_sel_0_; 
wire AES_CORE_CONTROL_UNIT_sbox_sel_1_; 
wire AES_CORE_CONTROL_UNIT_sbox_sel_2_; 
wire AES_CORE_CONTROL_UNIT_state_0_; 
wire AES_CORE_CONTROL_UNIT_state_11_; 
wire AES_CORE_CONTROL_UNIT_state_12_; 
wire AES_CORE_CONTROL_UNIT_state_13_; 
wire AES_CORE_CONTROL_UNIT_state_14_; 
wire AES_CORE_CONTROL_UNIT_state_15_; 
wire AES_CORE_CONTROL_UNIT_state_1_; 
wire AES_CORE_CONTROL_UNIT_state_2_; 
wire AES_CORE_CONTROL_UNIT_state_3_; 
wire AES_CORE_CONTROL_UNIT_state_4_; 
wire AES_CORE_CONTROL_UNIT_state_6_; 
wire AES_CORE_CONTROL_UNIT_state_7_; 
wire AES_CORE_CONTROL_UNIT_state_8_; 
wire AES_CORE_CONTROL_UNIT_state_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1000_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1001_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1003_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1004_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1006_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1007_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1008_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1010_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1011_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1013_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1014_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1015_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1017_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1018_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1020_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1021_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1022_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1024_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1025_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1026_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1028_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1029_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1030_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1032_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1033_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1034_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1036_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1037_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1038_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1040_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1041_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1042_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1044_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1045_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1046_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1048_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1049_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1050_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1052_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1053_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1054_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1056_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1057_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1058_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1060_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1061_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1062_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1064_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1065_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1066_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1068_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1069_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1070_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1072_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1073_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1074_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1076_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1077_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1078_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1080_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1081_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1082_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1084_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1085_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1086_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1088_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1089_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1090_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1092_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1093_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1094_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1096_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1097_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1098_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1100_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1101_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1102_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1104_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1105_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1106_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1108_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1109_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1110_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1112_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1113_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1114_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1116_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1117_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1118_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1120_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1121_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1122_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1124_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1125_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1126_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1128_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1129_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1130_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1132_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1133_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1134_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1135_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1137_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1138_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1139_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1141_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1142_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1143_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1144_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1146_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1147_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1148_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1150_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1151_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1152_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1154_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1155_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1156_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1158_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1159_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1160_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1162_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1163_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1164_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1166_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1167_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1168_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1170_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1171_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1172_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1174_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1175_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1176_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1178_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1179_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1180_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1182_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1183_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1184_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1186_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1187_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1188_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1190_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1191_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1192_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1194_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1195_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1196_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1198_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1199_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1200_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1202_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1203_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1204_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1206_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1207_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1208_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1210_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1211_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1212_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1214_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1215_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1216_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1218_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1219_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1220_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1222_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1223_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1224_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1226_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1227_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1228_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1230_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1231_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1232_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1234_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1235_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1236_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1238_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1239_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1240_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1242_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1243_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1244_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1246_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1247_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1248_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1250_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1251_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1252_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1254_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1255_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1256_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1258_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1259_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1260_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1262_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1263_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1264_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1266_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1267_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1268_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1270_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1271_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1272_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1274_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1275_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1276_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n327_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n328_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n329_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n330_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n331_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n332_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n333_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n334_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n335_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n336_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n338_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n339_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n340_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n341_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n342_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n343_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n344_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n345_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n346_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n347_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n349_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n350_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n351_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n352_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n353_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n354_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n355_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n356_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n357_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n358_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n360_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n361_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n362_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n363_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n364_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n365_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n366_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n367_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n368_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n369_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n371_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n372_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n373_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n374_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n375_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n376_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n377_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n378_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n379_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n380_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n382_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n383_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n384_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n385_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n386_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n387_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n388_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n389_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n390_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n391_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n393_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n394_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n395_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n396_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n397_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n398_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n399_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n400_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n401_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n402_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n404_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n405_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n406_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n407_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n408_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n409_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n410_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n411_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n412_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n413_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n415_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n416_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n417_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n418_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n419_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n420_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n421_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n422_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n423_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n424_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n426_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n427_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n428_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n429_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n430_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n431_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n432_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n433_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n434_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n435_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n437_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n438_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n439_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n440_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n441_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n442_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n443_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n444_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n445_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n446_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n448_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n449_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n450_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n451_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n452_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n453_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n454_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n455_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n456_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n457_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n459_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n460_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n461_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n462_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n463_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n464_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n465_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n466_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n467_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n468_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n470_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n471_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n472_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n473_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n474_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n475_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n476_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n477_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n478_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n479_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n481_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n482_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n483_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n484_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n485_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n486_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n487_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n488_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n489_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n490_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n492_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n493_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n494_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n495_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n496_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n497_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n498_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n499_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n500_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n501_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n503_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n504_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n505_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n506_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n507_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n508_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n509_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n510_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n511_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n512_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n514_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n515_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n516_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n517_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n518_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n519_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n520_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n521_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n522_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n523_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n525_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n526_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n527_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n528_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n529_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n530_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n531_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n532_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n533_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n534_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n536_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n537_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n538_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n539_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n540_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n541_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n542_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n543_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n544_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n545_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n547_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n548_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n549_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n550_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n551_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n552_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n553_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n554_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n555_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n556_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n558_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n559_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n560_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n561_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n562_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n563_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n564_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n565_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n566_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n567_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n569_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n570_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n571_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n572_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n573_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n574_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n575_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n576_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n577_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n578_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n580_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n581_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n582_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n583_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n584_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n585_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n586_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n587_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n588_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n589_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n591_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n592_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n593_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n594_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n595_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n596_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n597_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n599_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n600_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n601_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n602_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n603_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n604_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n605_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n606_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n607_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n608_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n609_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n610_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n611_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n612_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n613_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n614_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n616_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n617_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n618_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n619_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n620_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n621_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n622_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n623_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n624_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n625_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n626_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n627_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n628_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n629_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n630_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n631_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n632_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n633_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n634_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n635_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n636_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n637_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n638_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n639_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n640_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n641_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n643_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n644_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n645_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n646_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n648_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n649_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n650_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n651_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n652_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n653_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n654_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n655_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n656_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n657_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n658_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n659_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n660_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n661_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n662_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n663_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n664_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n665_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n666_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n667_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n668_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n669_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n670_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n671_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n672_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n673_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n674_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n675_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n676_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n677_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n678_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n679_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n680_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n681_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n682_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n683_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n684_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n685_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n686_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n687_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n688_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n689_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n690_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n692_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n693_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n694_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n695_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n696_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n697_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n698_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n699_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n700_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n701_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n702_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n703_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n704_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n705_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n706_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n707_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n708_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n709_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n710_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n711_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n713_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n714_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n715_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n716_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n717_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n718_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n719_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n720_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n721_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n722_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n723_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n724_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n725_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n726_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n727_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n728_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n729_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n730_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n731_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n732_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n733_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n735_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n736_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n737_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n738_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n739_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n740_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n741_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n742_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n743_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n744_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n745_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n746_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n747_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n748_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n749_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n750_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n751_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n752_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n753_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n754_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n755_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n756_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n757_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n759_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n760_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n761_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n762_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n763_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n764_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n765_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n766_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n767_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n768_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n769_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n770_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n771_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n772_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n773_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n774_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n776_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n777_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n778_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n779_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n780_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n781_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n782_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n783_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n784_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n785_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n786_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n787_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n788_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n789_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n790_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n791_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n792_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n793_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n794_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n796_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n797_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n798_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n800_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n801_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n803_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n804_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n805_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n807_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n808_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n810_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n811_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n812_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n814_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n815_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n817_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n818_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n819_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n821_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n822_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n824_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n825_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n826_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n828_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n829_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n831_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n832_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n833_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n835_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n836_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n838_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n839_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n840_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n842_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n843_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n845_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n846_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n847_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n849_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n850_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n852_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n853_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n854_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n856_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n857_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n859_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n860_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n861_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n863_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n864_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n866_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n867_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n868_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n870_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n871_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n873_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n874_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n875_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n877_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n878_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n880_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n881_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n882_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n884_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n885_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n887_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n888_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n889_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n891_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n892_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n894_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n895_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n896_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n898_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n899_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n901_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n902_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n903_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n905_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n906_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n908_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n909_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n910_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n912_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n913_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n915_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n916_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n917_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n919_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n920_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n922_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n923_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n924_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n926_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n927_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n929_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n930_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n931_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n933_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n934_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n936_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n937_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n938_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n940_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n941_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n943_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n944_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n945_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n947_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n948_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n950_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n951_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n952_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n954_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n955_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n957_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n958_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n959_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n961_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n962_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n964_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n965_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n966_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n968_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n969_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n971_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n972_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n973_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n975_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n976_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n978_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n979_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n980_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n982_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n983_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n985_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n986_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n987_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n989_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n990_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n992_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n993_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n994_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n996_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n997_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n999_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_0_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_1_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_2_; 
wire AES_CORE_DATAPATH_KEY_EXPANDER_round_3_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n100_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n101_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n102_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n103_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n104_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n105_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n106_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n108_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n109_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n110_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n111_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n112_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n113_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n114_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n115_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n116_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n117_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n119_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n120_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n121_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n122_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n123_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n125_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n126_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n127_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n128_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n129_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n130_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n131_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n133_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n134_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n136_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n137_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n138_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n139_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n140_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n142_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n144_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n145_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n146_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n148_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n149_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n151_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n153_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n154_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n155_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n157_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n159_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n161_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n162_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n163_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n164_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n165_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n166_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n167_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n168_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n169_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n170_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n171_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n172_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n173_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n174_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n176_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n177_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n178_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n179_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n180_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n181_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n182_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n183_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n185_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n186_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n187_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n189_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n191_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n193_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n196_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n197_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n198_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n200_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n201_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n202_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n204_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n205_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n206_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n207_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n208_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n210_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n211_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n212_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n213_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n214_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n215_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n216_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n217_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n218_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n219_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n221_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n222_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n223_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n224_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n225_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n226_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n227_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n228_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n229_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n231_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n232_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n233_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n234_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n235_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n236_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n237_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n239_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n240_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n241_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n242_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n243_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n244_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n245_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n246_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n247_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n248_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n249_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n250_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n252_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n253_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n254_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n256_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n257_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n258_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n259_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n260_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n261_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n262_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n263_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n264_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n265_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n266_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n267_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n268_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n269_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n270_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n271_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n272_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n273_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n274_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n276_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n277_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n278_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n279_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n280_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n281_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n282_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n283_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n284_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n286_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n287_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n288_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n289_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n290_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n291_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n292_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n293_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n294_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n295_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n296_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n297_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n298_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n300_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n301_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n302_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n303_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n304_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n305_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n306_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n307_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n308_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n309_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n310_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n311_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n312_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n313_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n314_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n315_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n316_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n317_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n318_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n319_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n320_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n321_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n322_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n323_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n324_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n325_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n326_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n327_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n328_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n329_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n330_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n331_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n332_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n333_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n334_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n335_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n336_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n337_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n339_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n340_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n341_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n342_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n343_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n344_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n345_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n346_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n347_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n348_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n349_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n350_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n351_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n353_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n354_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n355_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n356_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n357_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n358_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n359_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n360_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n361_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n363_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n364_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n365_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n366_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n367_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n368_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n369_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n370_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n371_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n372_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n373_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n374_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n375_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n376_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n377_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n378_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n379_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n380_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n381_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n382_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n383_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n384_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n385_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n386_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n387_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n388_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n389_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n390_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n391_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n392_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n393_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n394_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n395_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n396_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n397_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n398_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n399_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n401_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n402_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n403_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n404_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n405_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n406_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n407_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n408_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n409_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n410_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n411_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n412_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n414_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n415_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n416_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n417_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n418_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n419_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n420_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n421_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n422_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n423_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n424_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n425_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n426_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n427_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n428_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n429_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n430_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n431_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n432_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n433_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n434_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n435_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n436_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n437_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n438_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n439_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n440_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n441_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n442_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n444_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n445_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n446_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n447_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n448_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n449_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n450_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n451_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n452_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n453_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n454_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n455_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n456_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n457_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n459_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n460_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n461_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n463_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n464_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n465_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n466_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n467_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n468_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n469_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n470_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n471_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n472_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n473_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n474_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n475_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n476_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n477_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n479_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n480_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n481_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n482_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n483_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n484_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n485_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n486_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n487_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n488_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n490_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n491_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n492_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n493_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n494_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n495_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n496_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n497_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n498_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n499_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n500_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n502_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n503_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n505_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n506_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n507_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n508_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n509_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n511_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n513_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n514_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n515_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n516_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n517_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n518_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n519_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n521_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n522_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n523_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n524_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n525_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n526_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n527_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n528_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n529_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n530_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n531_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n532_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n533_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n534_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n535_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n537_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n538_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n539_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n540_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n541_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n542_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n544_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n545_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n546_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n547_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n548_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n549_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n550_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n551_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n552_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n553_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n555_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n556_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n557_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n558_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n559_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n560_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n561_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n563_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n564_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n565_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n566_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n567_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n568_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n569_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n570_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n571_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n572_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n573_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n574_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n575_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n576_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n578_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n579_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n580_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n581_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n582_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n583_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n584_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n585_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n586_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n588_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n589_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n590_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n591_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n592_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n593_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n594_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n595_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n596_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n597_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n598_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n599_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n600_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n601_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n603_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n604_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n605_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n606_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n607_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n608_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n609_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n610_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n611_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n613_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n614_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n615_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n616_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n617_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n618_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n619_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n620_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n621_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n622_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n624_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n625_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n626_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n627_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n628_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n629_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n630_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n631_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n632_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n634_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n635_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n636_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n637_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n638_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n639_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n640_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n641_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n642_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n643_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n644_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n646_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n647_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n648_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n649_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n650_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n651_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n653_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n654_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n655_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n656_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n657_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n658_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n660_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n661_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n662_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n663_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n664_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n665_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n666_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n667_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n669_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n670_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n671_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n672_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n673_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n674_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n676_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n677_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n678_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n679_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n680_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n681_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n682_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n683_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n685_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n687_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n688_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n689_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n691_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n692_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n693_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n694_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n695_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n696_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n697_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n698_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n699_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n700_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n701_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n702_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n703_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n704_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n705_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n707_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n708_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n710_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n711_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n712_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n713_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n714_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n715_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n716_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n717_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n718_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n719_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n721_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n722_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n723_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n725_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n726_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n727_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n728_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n729_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n730_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n731_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n732_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n733_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n734_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n735_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n736_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n737_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n739_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n740_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n741_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n743_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n744_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n745_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n746_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n747_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n748_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n749_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n750_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n751_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n752_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n753_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n754_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n755_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n756_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n757_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n759_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n760_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n762_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n763_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n764_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n765_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n766_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n767_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n768_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n769_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n770_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n771_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n772_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n774_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n775_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n777_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n778_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n779_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n780_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n781_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n782_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n783_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n784_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n785_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n786_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n788_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n789_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n790_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n792_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n793_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n794_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n795_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n796_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n797_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n798_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n799_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n800_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n801_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n802_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n804_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n805_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n807_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n808_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n809_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n810_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n811_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n812_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n814_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n815_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n816_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n818_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n819_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n820_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n821_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n822_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n823_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n824_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n825_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n826_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n827_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n828_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n829_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n830_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n831_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n832_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n834_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n835_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n837_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n838_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n839_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n840_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n841_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n842_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n843_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n844_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n845_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n846_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n847_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n849_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n850_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n852_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n853_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n854_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n855_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n856_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n857_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n858_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n859_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n860_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n861_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n862_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n863_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n864_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n865_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n867_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n868_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n869_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n871_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n872_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n873_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n874_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n875_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n876_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n877_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n878_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n879_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n880_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n881_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n882_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n883_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n884_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n885_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n887_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n888_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n890_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n891_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n892_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n893_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n894_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n895_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n896_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n897_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n898_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n899_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n900_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n902_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n903_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n905_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n906_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n907_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n908_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n909_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n910_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n911_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n912_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n913_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n914_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n916_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n917_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n918_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n920_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n921_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n922_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n923_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n924_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n925_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n926_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n928_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n929_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n97_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n98_; 
wire AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n99_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_0__7_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_1__7_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_2__7_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__0_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__1_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__2_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__3_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__4_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__5_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__6_; 
wire AES_CORE_DATAPATH_MIX_COL_col_3__7_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_; 
wire AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n108_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n120_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n124_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n126_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n134_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n225_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n276_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n283_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n314_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n325_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n338_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n345_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n346_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n350_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n363_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n367_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n384_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n422_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n455_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n475_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n490_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n499_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n501_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n502_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n503_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n504_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n505_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n506_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n507_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n508_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n509_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n510_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n511_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n512_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n513_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n514_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n515_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n516_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n518_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n519_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n520_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n521_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n522_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n523_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n524_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n525_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n526_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n527_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n528_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n529_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n530_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n531_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n532_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n533_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n535_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n536_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n537_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n538_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n539_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n540_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n541_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n542_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n543_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n544_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n545_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n546_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n547_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n548_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n550_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n551_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n552_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n554_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n555_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n68_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n83_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n96_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n108_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n120_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n124_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n126_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n134_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n225_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n276_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n283_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n314_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n325_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n338_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n345_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n346_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n350_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n363_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n367_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n384_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n422_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n455_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n475_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n490_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n499_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n501_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n502_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n503_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n504_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n505_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n506_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n507_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n508_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n509_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n510_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n511_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n512_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n513_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n514_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n515_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n516_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n518_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n519_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n520_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n521_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n522_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n523_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n524_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n525_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n526_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n527_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n528_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n529_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n530_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n531_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n532_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n533_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n535_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n536_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n537_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n538_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n539_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n540_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n541_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n542_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n543_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n544_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n545_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n546_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n547_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n548_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n550_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n551_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n552_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n554_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n555_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n68_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n83_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n96_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n108_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n120_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n124_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n126_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n134_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n225_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n276_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n283_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n314_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n325_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n338_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n345_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n346_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n350_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n363_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n367_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n384_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n422_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n455_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n475_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n490_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n499_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n501_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n502_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n503_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n504_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n505_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n506_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n507_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n508_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n509_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n510_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n511_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n512_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n513_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n514_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n515_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n516_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n518_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n519_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n520_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n521_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n522_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n523_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n524_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n525_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n526_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n527_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n528_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n529_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n530_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n531_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n532_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n533_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n535_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n536_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n537_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n538_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n539_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n540_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n541_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n542_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n543_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n544_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n545_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n546_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n547_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n548_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n550_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n551_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n552_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n554_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n555_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n68_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n83_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n96_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n100_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n102_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n103_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n104_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n105_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n106_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n107_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n108_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n109_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n110_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n111_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n112_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n113_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n114_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n115_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n117_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n118_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n119_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n120_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n121_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n122_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n123_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n124_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n125_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n126_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n128_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n129_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n130_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n131_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n132_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n133_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n134_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n135_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n136_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n138_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n139_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n140_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n142_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n143_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n144_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n145_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n146_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n147_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n148_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n149_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n150_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n151_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n152_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n153_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n154_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n156_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n157_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n158_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n159_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n160_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n161_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n162_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n163_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n164_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n166_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n167_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n168_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n169_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n170_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n171_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n172_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n173_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n174_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n175_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n177_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n178_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n179_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n180_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n181_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n182_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n183_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n184_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n185_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n186_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n187_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n188_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n189_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n190_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n191_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n192_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n193_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n194_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n195_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n196_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n197_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n198_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n199_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n200_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n201_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n202_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n204_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n205_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n206_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n207_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n208_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n209_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n210_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n211_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n212_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n213_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n214_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n215_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n216_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n217_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n218_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n219_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n220_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n221_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n222_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n223_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n224_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n225_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n226_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n227_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n228_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n229_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n230_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n231_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n232_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n233_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n234_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n235_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n236_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n237_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n238_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n239_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n240_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n241_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n242_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n243_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n246_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n247_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n248_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n249_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n250_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n251_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n252_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n253_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n254_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n255_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n256_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n257_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n258_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n259_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n260_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n261_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n262_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n263_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n264_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n265_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n266_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n267_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n268_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n269_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n270_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n271_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n272_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n273_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n274_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n275_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n276_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n277_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n279_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n280_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n281_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n282_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n283_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n284_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n285_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n286_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n287_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n288_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n289_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n290_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n291_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n292_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n293_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n294_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n295_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n296_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n297_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n298_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n299_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n300_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n302_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n303_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n304_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n305_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n306_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n307_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n308_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n309_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n310_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n311_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n312_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n313_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n314_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n315_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n316_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n317_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n318_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n319_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n320_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n321_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n323_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n324_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n325_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n326_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n327_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n328_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n329_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n330_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n331_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n332_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n333_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n334_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n335_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n337_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n338_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n339_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n340_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n341_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n342_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n343_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n344_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n345_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n346_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n347_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n348_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n349_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n350_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n351_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n352_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n353_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n354_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n355_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n356_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n357_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n358_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n359_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n360_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n361_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n362_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n363_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n364_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n365_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n366_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n367_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n369_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n370_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n371_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n372_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n373_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n374_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n376_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n378_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n379_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n380_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n381_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n382_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n383_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n384_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n385_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n386_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n387_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n389_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n390_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n391_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n392_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n393_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n394_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n395_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n396_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n397_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n398_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n399_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n400_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n401_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n402_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n404_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n405_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n406_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n407_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n408_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n409_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n410_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n411_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n412_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n414_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n416_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n417_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n418_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n420_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n421_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n422_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n423_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n424_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n425_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n426_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n427_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n429_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n430_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n432_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n433_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n435_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n436_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n438_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n439_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n440_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n442_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n443_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n444_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n445_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n446_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n447_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n448_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n449_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n450_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n451_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n452_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n453_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n454_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n455_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n456_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n457_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n458_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n459_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n460_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n461_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n462_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n463_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n464_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n465_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n466_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n468_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n469_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n470_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n471_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n472_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n473_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n474_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n475_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n476_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n477_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n478_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n479_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n480_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n481_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n482_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n483_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n485_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n486_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n487_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n488_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n489_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n490_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n491_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n492_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n493_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n494_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n495_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n496_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n497_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n498_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n499_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n500_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n501_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n502_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n503_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n504_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n505_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n506_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n507_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n508_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n509_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n50_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n510_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n511_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n512_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n513_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n514_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n515_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n516_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n518_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n519_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n51_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n520_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n521_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n522_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n523_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n524_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n525_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n526_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n527_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n528_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n529_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n52_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n530_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n531_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n532_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n533_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n535_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n536_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n537_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n538_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n539_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n53_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n540_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n541_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n542_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n543_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n544_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n545_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n546_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n547_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n548_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n54_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n550_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n551_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n552_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n554_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n555_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n55_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n56_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n57_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n58_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n59_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n60_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n61_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n62_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n63_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n64_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n65_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n67_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n68_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n69_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n70_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n71_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n72_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n73_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n74_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n75_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n76_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n78_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n80_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n81_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n82_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n83_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n84_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n85_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n86_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n87_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n88_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n90_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n91_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n92_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n93_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n94_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n95_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n96_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n97_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n98_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n99_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_; 
wire AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_; 
wire AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n101_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n102_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n103_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n104_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n105_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n106_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n108_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n109_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n110_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n111_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n112_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n113_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n115_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n116_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n117_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n118_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n119_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n120_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n122_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n123_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n124_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n125_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n126_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n127_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n129_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n130_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n131_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n132_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n133_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n134_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n136_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n137_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n138_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n139_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n140_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n141_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n143_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n144_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n145_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n146_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n147_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n148_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n150_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n151_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n152_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n153_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n154_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n155_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n157_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n158_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n159_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n160_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n161_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n162_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n164_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n165_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n166_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n167_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n168_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n169_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n171_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n172_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n173_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n174_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n175_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n176_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n178_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n179_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n180_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n181_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n182_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n183_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n185_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n186_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n187_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n188_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n189_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n190_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n192_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n193_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n194_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n195_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n196_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n197_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n199_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n200_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n201_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n202_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n203_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n204_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n206_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n207_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n208_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n209_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n210_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n211_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n213_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n214_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n215_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n216_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n217_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n218_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n220_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n221_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n222_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n223_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n224_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n225_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n227_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n228_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n229_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n230_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n231_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n232_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n234_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n235_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n236_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n237_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n238_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n239_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n241_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n242_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n243_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n244_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n245_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n246_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n248_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n249_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n250_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n251_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n252_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n253_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n255_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n256_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n257_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n258_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n259_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n260_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n262_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n263_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n264_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n265_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n266_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n267_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n269_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n270_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n271_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n272_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n273_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n274_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n276_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n277_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n278_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n279_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n280_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n281_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n283_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n284_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n285_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n286_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n287_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n288_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n290_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n291_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n292_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n293_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n294_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n295_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n67_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n69_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n70_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n72_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n73_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n75_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n77_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n78_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n80_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n81_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n82_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n83_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n84_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n85_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n87_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n88_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n89_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n90_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n91_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n92_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n94_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n95_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n96_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n97_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n98_; 
wire AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n99_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_0_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_10_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_11_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_12_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_13_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_14_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_15_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_16_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_17_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_18_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_19_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_1_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_20_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_21_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_22_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_23_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_24_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_25_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_26_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_27_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_28_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_29_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_2_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_30_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_31_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_3_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_4_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_5_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_6_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_7_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_8_; 
wire AES_CORE_DATAPATH_SWAP_IN_data_swap_9_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n101_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n102_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n103_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n104_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n105_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n106_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n108_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n109_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n110_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n111_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n112_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n113_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n115_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n116_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n117_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n118_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n119_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n120_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n122_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n123_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n124_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n125_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n126_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n127_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n129_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n130_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n131_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n132_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n133_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n134_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n136_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n137_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n138_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n139_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n140_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n141_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n143_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n144_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n145_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n146_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n147_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n148_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n150_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n151_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n152_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n153_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n154_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n155_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n157_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n158_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n159_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n160_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n161_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n162_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n164_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n165_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n166_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n167_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n168_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n169_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n171_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n172_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n173_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n174_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n175_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n176_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n178_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n179_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n180_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n181_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n182_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n183_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n185_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n186_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n187_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n188_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n189_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n190_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n192_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n193_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n194_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n195_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n196_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n197_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n199_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n200_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n201_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n202_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n203_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n204_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n206_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n207_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n208_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n209_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n210_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n211_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n213_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n214_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n215_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n216_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n217_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n218_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n220_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n221_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n222_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n223_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n224_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n225_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n227_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n228_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n229_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n230_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n231_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n232_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n234_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n235_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n236_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n237_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n238_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n239_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n241_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n242_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n243_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n244_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n245_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n246_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n248_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n249_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n250_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n251_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n252_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n253_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n255_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n256_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n257_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n258_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n259_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n260_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n262_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n263_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n264_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n265_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n266_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n267_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n269_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n270_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n271_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n272_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n273_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n274_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n276_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n277_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n278_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n279_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n280_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n281_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n283_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n284_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n285_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n286_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n287_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n288_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n290_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n291_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n292_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n293_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n294_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n295_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n67_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n69_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n70_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n72_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n73_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n75_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n77_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n78_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n80_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n81_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n82_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n83_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n84_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n85_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n87_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n88_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n89_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n90_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n91_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n92_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n94_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n95_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n96_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n97_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n98_; 
wire AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n99_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_0__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_0__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_1__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_2__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1_3__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_1__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_2__31_0__9_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__0_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__10_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__11_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__12_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__13_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__14_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__15_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__16_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__17_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__18_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__19_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__1_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__20_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__21_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__22_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__23_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__24_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__25_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__26_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__27_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__28_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__29_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__2_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__30_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__31_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__3_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__4_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__5_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__6_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__7_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__8_; 
wire AES_CORE_DATAPATH__0bkp_3__31_0__9_; 
wire AES_CORE_DATAPATH__0col_0__31_0__0_; 
wire AES_CORE_DATAPATH__0col_0__31_0__10_; 
wire AES_CORE_DATAPATH__0col_0__31_0__11_; 
wire AES_CORE_DATAPATH__0col_0__31_0__12_; 
wire AES_CORE_DATAPATH__0col_0__31_0__13_; 
wire AES_CORE_DATAPATH__0col_0__31_0__14_; 
wire AES_CORE_DATAPATH__0col_0__31_0__15_; 
wire AES_CORE_DATAPATH__0col_0__31_0__16_; 
wire AES_CORE_DATAPATH__0col_0__31_0__17_; 
wire AES_CORE_DATAPATH__0col_0__31_0__18_; 
wire AES_CORE_DATAPATH__0col_0__31_0__19_; 
wire AES_CORE_DATAPATH__0col_0__31_0__1_; 
wire AES_CORE_DATAPATH__0col_0__31_0__20_; 
wire AES_CORE_DATAPATH__0col_0__31_0__21_; 
wire AES_CORE_DATAPATH__0col_0__31_0__22_; 
wire AES_CORE_DATAPATH__0col_0__31_0__23_; 
wire AES_CORE_DATAPATH__0col_0__31_0__24_; 
wire AES_CORE_DATAPATH__0col_0__31_0__25_; 
wire AES_CORE_DATAPATH__0col_0__31_0__26_; 
wire AES_CORE_DATAPATH__0col_0__31_0__27_; 
wire AES_CORE_DATAPATH__0col_0__31_0__28_; 
wire AES_CORE_DATAPATH__0col_0__31_0__29_; 
wire AES_CORE_DATAPATH__0col_0__31_0__2_; 
wire AES_CORE_DATAPATH__0col_0__31_0__30_; 
wire AES_CORE_DATAPATH__0col_0__31_0__31_; 
wire AES_CORE_DATAPATH__0col_0__31_0__3_; 
wire AES_CORE_DATAPATH__0col_0__31_0__4_; 
wire AES_CORE_DATAPATH__0col_0__31_0__5_; 
wire AES_CORE_DATAPATH__0col_0__31_0__6_; 
wire AES_CORE_DATAPATH__0col_0__31_0__7_; 
wire AES_CORE_DATAPATH__0col_0__31_0__8_; 
wire AES_CORE_DATAPATH__0col_0__31_0__9_; 
wire AES_CORE_DATAPATH__0col_1__31_0__0_; 
wire AES_CORE_DATAPATH__0col_1__31_0__10_; 
wire AES_CORE_DATAPATH__0col_1__31_0__11_; 
wire AES_CORE_DATAPATH__0col_1__31_0__12_; 
wire AES_CORE_DATAPATH__0col_1__31_0__13_; 
wire AES_CORE_DATAPATH__0col_1__31_0__14_; 
wire AES_CORE_DATAPATH__0col_1__31_0__15_; 
wire AES_CORE_DATAPATH__0col_1__31_0__16_; 
wire AES_CORE_DATAPATH__0col_1__31_0__17_; 
wire AES_CORE_DATAPATH__0col_1__31_0__18_; 
wire AES_CORE_DATAPATH__0col_1__31_0__19_; 
wire AES_CORE_DATAPATH__0col_1__31_0__1_; 
wire AES_CORE_DATAPATH__0col_1__31_0__20_; 
wire AES_CORE_DATAPATH__0col_1__31_0__21_; 
wire AES_CORE_DATAPATH__0col_1__31_0__22_; 
wire AES_CORE_DATAPATH__0col_1__31_0__23_; 
wire AES_CORE_DATAPATH__0col_1__31_0__24_; 
wire AES_CORE_DATAPATH__0col_1__31_0__25_; 
wire AES_CORE_DATAPATH__0col_1__31_0__26_; 
wire AES_CORE_DATAPATH__0col_1__31_0__27_; 
wire AES_CORE_DATAPATH__0col_1__31_0__28_; 
wire AES_CORE_DATAPATH__0col_1__31_0__29_; 
wire AES_CORE_DATAPATH__0col_1__31_0__2_; 
wire AES_CORE_DATAPATH__0col_1__31_0__30_; 
wire AES_CORE_DATAPATH__0col_1__31_0__31_; 
wire AES_CORE_DATAPATH__0col_1__31_0__3_; 
wire AES_CORE_DATAPATH__0col_1__31_0__4_; 
wire AES_CORE_DATAPATH__0col_1__31_0__5_; 
wire AES_CORE_DATAPATH__0col_1__31_0__6_; 
wire AES_CORE_DATAPATH__0col_1__31_0__7_; 
wire AES_CORE_DATAPATH__0col_1__31_0__8_; 
wire AES_CORE_DATAPATH__0col_1__31_0__9_; 
wire AES_CORE_DATAPATH__0col_2__31_0__0_; 
wire AES_CORE_DATAPATH__0col_2__31_0__10_; 
wire AES_CORE_DATAPATH__0col_2__31_0__11_; 
wire AES_CORE_DATAPATH__0col_2__31_0__12_; 
wire AES_CORE_DATAPATH__0col_2__31_0__13_; 
wire AES_CORE_DATAPATH__0col_2__31_0__14_; 
wire AES_CORE_DATAPATH__0col_2__31_0__15_; 
wire AES_CORE_DATAPATH__0col_2__31_0__16_; 
wire AES_CORE_DATAPATH__0col_2__31_0__17_; 
wire AES_CORE_DATAPATH__0col_2__31_0__18_; 
wire AES_CORE_DATAPATH__0col_2__31_0__19_; 
wire AES_CORE_DATAPATH__0col_2__31_0__1_; 
wire AES_CORE_DATAPATH__0col_2__31_0__20_; 
wire AES_CORE_DATAPATH__0col_2__31_0__21_; 
wire AES_CORE_DATAPATH__0col_2__31_0__22_; 
wire AES_CORE_DATAPATH__0col_2__31_0__23_; 
wire AES_CORE_DATAPATH__0col_2__31_0__24_; 
wire AES_CORE_DATAPATH__0col_2__31_0__25_; 
wire AES_CORE_DATAPATH__0col_2__31_0__26_; 
wire AES_CORE_DATAPATH__0col_2__31_0__27_; 
wire AES_CORE_DATAPATH__0col_2__31_0__28_; 
wire AES_CORE_DATAPATH__0col_2__31_0__29_; 
wire AES_CORE_DATAPATH__0col_2__31_0__2_; 
wire AES_CORE_DATAPATH__0col_2__31_0__30_; 
wire AES_CORE_DATAPATH__0col_2__31_0__31_; 
wire AES_CORE_DATAPATH__0col_2__31_0__3_; 
wire AES_CORE_DATAPATH__0col_2__31_0__4_; 
wire AES_CORE_DATAPATH__0col_2__31_0__5_; 
wire AES_CORE_DATAPATH__0col_2__31_0__6_; 
wire AES_CORE_DATAPATH__0col_2__31_0__7_; 
wire AES_CORE_DATAPATH__0col_2__31_0__8_; 
wire AES_CORE_DATAPATH__0col_2__31_0__9_; 
wire AES_CORE_DATAPATH__0col_3__31_0__0_; 
wire AES_CORE_DATAPATH__0col_3__31_0__10_; 
wire AES_CORE_DATAPATH__0col_3__31_0__11_; 
wire AES_CORE_DATAPATH__0col_3__31_0__12_; 
wire AES_CORE_DATAPATH__0col_3__31_0__13_; 
wire AES_CORE_DATAPATH__0col_3__31_0__14_; 
wire AES_CORE_DATAPATH__0col_3__31_0__15_; 
wire AES_CORE_DATAPATH__0col_3__31_0__16_; 
wire AES_CORE_DATAPATH__0col_3__31_0__17_; 
wire AES_CORE_DATAPATH__0col_3__31_0__18_; 
wire AES_CORE_DATAPATH__0col_3__31_0__19_; 
wire AES_CORE_DATAPATH__0col_3__31_0__1_; 
wire AES_CORE_DATAPATH__0col_3__31_0__20_; 
wire AES_CORE_DATAPATH__0col_3__31_0__21_; 
wire AES_CORE_DATAPATH__0col_3__31_0__22_; 
wire AES_CORE_DATAPATH__0col_3__31_0__23_; 
wire AES_CORE_DATAPATH__0col_3__31_0__24_; 
wire AES_CORE_DATAPATH__0col_3__31_0__25_; 
wire AES_CORE_DATAPATH__0col_3__31_0__26_; 
wire AES_CORE_DATAPATH__0col_3__31_0__27_; 
wire AES_CORE_DATAPATH__0col_3__31_0__28_; 
wire AES_CORE_DATAPATH__0col_3__31_0__29_; 
wire AES_CORE_DATAPATH__0col_3__31_0__2_; 
wire AES_CORE_DATAPATH__0col_3__31_0__30_; 
wire AES_CORE_DATAPATH__0col_3__31_0__31_; 
wire AES_CORE_DATAPATH__0col_3__31_0__3_; 
wire AES_CORE_DATAPATH__0col_3__31_0__4_; 
wire AES_CORE_DATAPATH__0col_3__31_0__5_; 
wire AES_CORE_DATAPATH__0col_3__31_0__6_; 
wire AES_CORE_DATAPATH__0col_3__31_0__7_; 
wire AES_CORE_DATAPATH__0col_3__31_0__8_; 
wire AES_CORE_DATAPATH__0col_3__31_0__9_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__0_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__1_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__2_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__3_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__0_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__1_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__2_; 
wire AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__3_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_0__31_0__9_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_1__31_0__9_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_2__31_0__9_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__0_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__10_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__11_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__12_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__13_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__14_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__15_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__16_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__17_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__18_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__19_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__1_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__20_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__21_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__22_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__23_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__24_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__25_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__26_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__27_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__28_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__29_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__2_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__30_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__31_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__3_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__4_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__5_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__6_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__7_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__8_; 
wire AES_CORE_DATAPATH__0iv_3__31_0__9_; 
wire AES_CORE_DATAPATH__0key_0__31_0__0_; 
wire AES_CORE_DATAPATH__0key_0__31_0__10_; 
wire AES_CORE_DATAPATH__0key_0__31_0__11_; 
wire AES_CORE_DATAPATH__0key_0__31_0__12_; 
wire AES_CORE_DATAPATH__0key_0__31_0__13_; 
wire AES_CORE_DATAPATH__0key_0__31_0__14_; 
wire AES_CORE_DATAPATH__0key_0__31_0__15_; 
wire AES_CORE_DATAPATH__0key_0__31_0__16_; 
wire AES_CORE_DATAPATH__0key_0__31_0__17_; 
wire AES_CORE_DATAPATH__0key_0__31_0__18_; 
wire AES_CORE_DATAPATH__0key_0__31_0__19_; 
wire AES_CORE_DATAPATH__0key_0__31_0__1_; 
wire AES_CORE_DATAPATH__0key_0__31_0__20_; 
wire AES_CORE_DATAPATH__0key_0__31_0__21_; 
wire AES_CORE_DATAPATH__0key_0__31_0__22_; 
wire AES_CORE_DATAPATH__0key_0__31_0__23_; 
wire AES_CORE_DATAPATH__0key_0__31_0__24_; 
wire AES_CORE_DATAPATH__0key_0__31_0__25_; 
wire AES_CORE_DATAPATH__0key_0__31_0__26_; 
wire AES_CORE_DATAPATH__0key_0__31_0__27_; 
wire AES_CORE_DATAPATH__0key_0__31_0__28_; 
wire AES_CORE_DATAPATH__0key_0__31_0__29_; 
wire AES_CORE_DATAPATH__0key_0__31_0__2_; 
wire AES_CORE_DATAPATH__0key_0__31_0__30_; 
wire AES_CORE_DATAPATH__0key_0__31_0__31_; 
wire AES_CORE_DATAPATH__0key_0__31_0__3_; 
wire AES_CORE_DATAPATH__0key_0__31_0__4_; 
wire AES_CORE_DATAPATH__0key_0__31_0__5_; 
wire AES_CORE_DATAPATH__0key_0__31_0__6_; 
wire AES_CORE_DATAPATH__0key_0__31_0__7_; 
wire AES_CORE_DATAPATH__0key_0__31_0__8_; 
wire AES_CORE_DATAPATH__0key_0__31_0__9_; 
wire AES_CORE_DATAPATH__0key_1__31_0__0_; 
wire AES_CORE_DATAPATH__0key_1__31_0__10_; 
wire AES_CORE_DATAPATH__0key_1__31_0__11_; 
wire AES_CORE_DATAPATH__0key_1__31_0__12_; 
wire AES_CORE_DATAPATH__0key_1__31_0__13_; 
wire AES_CORE_DATAPATH__0key_1__31_0__14_; 
wire AES_CORE_DATAPATH__0key_1__31_0__15_; 
wire AES_CORE_DATAPATH__0key_1__31_0__16_; 
wire AES_CORE_DATAPATH__0key_1__31_0__17_; 
wire AES_CORE_DATAPATH__0key_1__31_0__18_; 
wire AES_CORE_DATAPATH__0key_1__31_0__19_; 
wire AES_CORE_DATAPATH__0key_1__31_0__1_; 
wire AES_CORE_DATAPATH__0key_1__31_0__20_; 
wire AES_CORE_DATAPATH__0key_1__31_0__21_; 
wire AES_CORE_DATAPATH__0key_1__31_0__22_; 
wire AES_CORE_DATAPATH__0key_1__31_0__23_; 
wire AES_CORE_DATAPATH__0key_1__31_0__24_; 
wire AES_CORE_DATAPATH__0key_1__31_0__25_; 
wire AES_CORE_DATAPATH__0key_1__31_0__26_; 
wire AES_CORE_DATAPATH__0key_1__31_0__27_; 
wire AES_CORE_DATAPATH__0key_1__31_0__28_; 
wire AES_CORE_DATAPATH__0key_1__31_0__29_; 
wire AES_CORE_DATAPATH__0key_1__31_0__2_; 
wire AES_CORE_DATAPATH__0key_1__31_0__30_; 
wire AES_CORE_DATAPATH__0key_1__31_0__31_; 
wire AES_CORE_DATAPATH__0key_1__31_0__3_; 
wire AES_CORE_DATAPATH__0key_1__31_0__4_; 
wire AES_CORE_DATAPATH__0key_1__31_0__5_; 
wire AES_CORE_DATAPATH__0key_1__31_0__6_; 
wire AES_CORE_DATAPATH__0key_1__31_0__7_; 
wire AES_CORE_DATAPATH__0key_1__31_0__8_; 
wire AES_CORE_DATAPATH__0key_1__31_0__9_; 
wire AES_CORE_DATAPATH__0key_2__31_0__0_; 
wire AES_CORE_DATAPATH__0key_2__31_0__10_; 
wire AES_CORE_DATAPATH__0key_2__31_0__11_; 
wire AES_CORE_DATAPATH__0key_2__31_0__12_; 
wire AES_CORE_DATAPATH__0key_2__31_0__13_; 
wire AES_CORE_DATAPATH__0key_2__31_0__14_; 
wire AES_CORE_DATAPATH__0key_2__31_0__15_; 
wire AES_CORE_DATAPATH__0key_2__31_0__16_; 
wire AES_CORE_DATAPATH__0key_2__31_0__17_; 
wire AES_CORE_DATAPATH__0key_2__31_0__18_; 
wire AES_CORE_DATAPATH__0key_2__31_0__19_; 
wire AES_CORE_DATAPATH__0key_2__31_0__1_; 
wire AES_CORE_DATAPATH__0key_2__31_0__20_; 
wire AES_CORE_DATAPATH__0key_2__31_0__21_; 
wire AES_CORE_DATAPATH__0key_2__31_0__22_; 
wire AES_CORE_DATAPATH__0key_2__31_0__23_; 
wire AES_CORE_DATAPATH__0key_2__31_0__24_; 
wire AES_CORE_DATAPATH__0key_2__31_0__25_; 
wire AES_CORE_DATAPATH__0key_2__31_0__26_; 
wire AES_CORE_DATAPATH__0key_2__31_0__27_; 
wire AES_CORE_DATAPATH__0key_2__31_0__28_; 
wire AES_CORE_DATAPATH__0key_2__31_0__29_; 
wire AES_CORE_DATAPATH__0key_2__31_0__2_; 
wire AES_CORE_DATAPATH__0key_2__31_0__30_; 
wire AES_CORE_DATAPATH__0key_2__31_0__31_; 
wire AES_CORE_DATAPATH__0key_2__31_0__3_; 
wire AES_CORE_DATAPATH__0key_2__31_0__4_; 
wire AES_CORE_DATAPATH__0key_2__31_0__5_; 
wire AES_CORE_DATAPATH__0key_2__31_0__6_; 
wire AES_CORE_DATAPATH__0key_2__31_0__7_; 
wire AES_CORE_DATAPATH__0key_2__31_0__8_; 
wire AES_CORE_DATAPATH__0key_2__31_0__9_; 
wire AES_CORE_DATAPATH__0key_3__31_0__0_; 
wire AES_CORE_DATAPATH__0key_3__31_0__10_; 
wire AES_CORE_DATAPATH__0key_3__31_0__11_; 
wire AES_CORE_DATAPATH__0key_3__31_0__12_; 
wire AES_CORE_DATAPATH__0key_3__31_0__13_; 
wire AES_CORE_DATAPATH__0key_3__31_0__14_; 
wire AES_CORE_DATAPATH__0key_3__31_0__15_; 
wire AES_CORE_DATAPATH__0key_3__31_0__16_; 
wire AES_CORE_DATAPATH__0key_3__31_0__17_; 
wire AES_CORE_DATAPATH__0key_3__31_0__18_; 
wire AES_CORE_DATAPATH__0key_3__31_0__19_; 
wire AES_CORE_DATAPATH__0key_3__31_0__1_; 
wire AES_CORE_DATAPATH__0key_3__31_0__20_; 
wire AES_CORE_DATAPATH__0key_3__31_0__21_; 
wire AES_CORE_DATAPATH__0key_3__31_0__22_; 
wire AES_CORE_DATAPATH__0key_3__31_0__23_; 
wire AES_CORE_DATAPATH__0key_3__31_0__24_; 
wire AES_CORE_DATAPATH__0key_3__31_0__25_; 
wire AES_CORE_DATAPATH__0key_3__31_0__26_; 
wire AES_CORE_DATAPATH__0key_3__31_0__27_; 
wire AES_CORE_DATAPATH__0key_3__31_0__28_; 
wire AES_CORE_DATAPATH__0key_3__31_0__29_; 
wire AES_CORE_DATAPATH__0key_3__31_0__2_; 
wire AES_CORE_DATAPATH__0key_3__31_0__30_; 
wire AES_CORE_DATAPATH__0key_3__31_0__31_; 
wire AES_CORE_DATAPATH__0key_3__31_0__3_; 
wire AES_CORE_DATAPATH__0key_3__31_0__4_; 
wire AES_CORE_DATAPATH__0key_3__31_0__5_; 
wire AES_CORE_DATAPATH__0key_3__31_0__6_; 
wire AES_CORE_DATAPATH__0key_3__31_0__7_; 
wire AES_CORE_DATAPATH__0key_3__31_0__8_; 
wire AES_CORE_DATAPATH__0key_3__31_0__9_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__0_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__1_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__2_; 
wire AES_CORE_DATAPATH__0key_en_pp1_3_0__3_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_0__31_0__9_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_1__31_0__9_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_2__31_0__9_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__0_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__10_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__11_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__12_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__13_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__14_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__15_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__16_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__17_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__18_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__19_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__1_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__20_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__21_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__22_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__23_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__24_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__25_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__26_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__27_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__28_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__29_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__2_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__30_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__31_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__3_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__4_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__5_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__6_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__7_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__8_; 
wire AES_CORE_DATAPATH__0key_host_3__31_0__9_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__0_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__10_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__11_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__12_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__13_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__14_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__15_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__16_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__17_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__18_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__19_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__1_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__20_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__21_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__22_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__23_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__24_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__25_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__26_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__27_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__28_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__29_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__2_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__30_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__31_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__3_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__4_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__5_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__6_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__7_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__8_; 
wire AES_CORE_DATAPATH__0sbox_pp2_31_0__9_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10010_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10018_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10042_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10054_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10058_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10060_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10066_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10082_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10090_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10110_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10114_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10126_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10130_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10139_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10154_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10160_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10166_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10172_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10178_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10184_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10190_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10202_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10208_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10210_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10218_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10220_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10226_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10235_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10238_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10244_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10250_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10260_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10275_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10280_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10299_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10307_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10310_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10323_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10347_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10360_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10363_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10371_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10377_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10395_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10407_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10410_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10413_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10419_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10425_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10427_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10431_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10437_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10440_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10443_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10449_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10452_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10455_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10458_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10467_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10476_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10485_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10491_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10500_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10512_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10530_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10540_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10552_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10564_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10570_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10576_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10588_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10600_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10612_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10620_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10659_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10660_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n10697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2458_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2467_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2470_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2476_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2485_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2491_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2494_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2512_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2534_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2552_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2558_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2564_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2576_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2582_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2588_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2606_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2612_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2659_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2668_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2677_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2686_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2692_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2695_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2704_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2708_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2713_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2716_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2722_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2731_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2732_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2736_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2749_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2763_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2769_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2772_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2781_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2785_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2787_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2793_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2799_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2808_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2810_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2817_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2826_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2832_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2835_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2841_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2844_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2853_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2857_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2881_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2883_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2889_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2905_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2910_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2928_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2929_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2937_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2947_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2953_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2960_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2961_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2964_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2969_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2977_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2985_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2993_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n2999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3001_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3009_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3017_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3018_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3042_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3054_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3060_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3066_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3081_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3090_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3110_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3114_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3126_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3139_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3153_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3160_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3169_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3177_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3178_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3193_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3210_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3216_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3218_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3234_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3235_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3243_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3250_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3255_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3258_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3260_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3267_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3275_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3279_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3291_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3299_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3303_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3307_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3313_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3319_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3322_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3323_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3325_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3331_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3337_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3340_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3343_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3347_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3349_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3355_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3358_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3360_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3361_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3363_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3367_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3371_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3373_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3376_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3377_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3379_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3385_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3391_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3394_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3395_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3397_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3403_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3407_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3410_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3413_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3419_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3422_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3425_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3427_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3431_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3437_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3440_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3443_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3446_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3449_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3452_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3455_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3458_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3470_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3476_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3485_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3491_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3494_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3500_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3510_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3530_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3534_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3540_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3552_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3558_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3564_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3570_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3582_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3588_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3600_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3606_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3612_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3620_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3630_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3660_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3668_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3677_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3680_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3686_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3692_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3695_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3700_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3708_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3710_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3713_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3716_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3720_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3722_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3731_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3732_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3740_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3749_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3760_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3763_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3769_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3772_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3781_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3785_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3790_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3793_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3799_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3808_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3810_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3817_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3826_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3835_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3841_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3844_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3848_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3853_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3857_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3860_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3866_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3878_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3881_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3884_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3889_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3902_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3905_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3910_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3914_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3920_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3929_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3932_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3937_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3938_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3950_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3953_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3961_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3964_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3969_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3974_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3977_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3985_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3993_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n3999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4001_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4009_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4010_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4017_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4018_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4042_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4054_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4058_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4060_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4066_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4081_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4082_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4090_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4110_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4114_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4126_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4130_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4153_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4154_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4160_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4166_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4169_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4172_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4177_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4178_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4190_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4193_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4202_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4208_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4210_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4218_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4220_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4226_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4234_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4238_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4243_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4244_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4250_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4255_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4258_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4260_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4275_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4279_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4291_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4303_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4307_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4310_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4313_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4316_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4319_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4322_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4323_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4325_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4328_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4334_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4337_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4340_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4343_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4346_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4347_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4349_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4352_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4355_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4358_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4360_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4361_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4364_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4367_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4370_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4371_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4373_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4377_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4379_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4382_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4385_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4388_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4391_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4394_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4397_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4400_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4403_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4406_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4407_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4410_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4413_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4419_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4422_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4425_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4431_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4437_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4443_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4446_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4449_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4452_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4455_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4458_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4467_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4470_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4476_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4485_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4491_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4494_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4500_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4512_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4530_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4558_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4564_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4570_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4576_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4582_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4588_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4600_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4606_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4612_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4620_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4630_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4660_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4680_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4692_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4700_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4708_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4710_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4716_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4720_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4732_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4736_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4760_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4763_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4769_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4772_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4781_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4787_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4790_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4793_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4799_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4800_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4808_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4810_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4817_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4826_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4832_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4835_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4841_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4844_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4853_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4860_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4866_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4878_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4881_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4884_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4889_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4896_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4902_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4905_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4914_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4920_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4929_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4932_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4938_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4947_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4950_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4953_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4960_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4961_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4969_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4974_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4977_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4985_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4992_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4993_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n4999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5001_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5010_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5017_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5042_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5058_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5060_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5066_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5082_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5110_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5114_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5130_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5139_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5154_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5177_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5210_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5216_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5218_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5234_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5243_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5255_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5258_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5260_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5267_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5279_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5280_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5291_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5303_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5307_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5310_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5313_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5316_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5319_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5322_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5325_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5328_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5331_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5334_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5337_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5340_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5343_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5346_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5349_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5352_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5355_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5358_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5360_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5361_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5363_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5364_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5367_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5370_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5373_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5376_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5379_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5382_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5385_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5388_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5391_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5394_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5397_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5400_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5403_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5406_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5410_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5422_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5427_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5440_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5510_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5534_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5540_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5620_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5659_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5668_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5677_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5680_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5686_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5692_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5695_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5700_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5704_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5710_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5713_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5716_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5722_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5731_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5736_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5740_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5749_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5760_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5763_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5769_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5772_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5781_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5785_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5787_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5790_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5793_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5799_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5800_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5808_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5817_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5826_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5832_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5835_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5841_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5844_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5848_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5853_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5857_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5866_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5878_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5881_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5883_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5884_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5889_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5896_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5902_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5905_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5914_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5920_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5928_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5929_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5932_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5937_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5938_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5947_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5950_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5953_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5961_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5964_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5969_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5974_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5977_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5985_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5992_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5993_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n5999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6001_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6009_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6017_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6018_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6042_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6054_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6058_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6066_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6081_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6082_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6090_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6114_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6126_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6130_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6139_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6153_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6154_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6166_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6169_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6172_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6177_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6178_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6184_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6190_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6193_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6202_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6208_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6216_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6218_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6220_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6226_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6234_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6235_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6238_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6243_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6244_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6250_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6255_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6258_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6267_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6275_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6279_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6280_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6291_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6299_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6303_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6307_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6313_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6316_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6319_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6322_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6323_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6325_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6328_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6331_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6334_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6337_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6340_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6343_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6346_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6347_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6349_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6352_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6355_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6358_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6361_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6363_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6364_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6367_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6370_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6371_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6373_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6376_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6377_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6379_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6382_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6385_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6388_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6391_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6394_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6395_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6397_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6400_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6403_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6406_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6407_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6413_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6419_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6422_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6425_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6427_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6431_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6437_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6440_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6443_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6446_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6449_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6452_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6455_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6458_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6467_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6470_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6476_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6485_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6491_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6494_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6500_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6512_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6530_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6534_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6540_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6552_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6558_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6564_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6570_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6576_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6582_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6588_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6600_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6606_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6612_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6620_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6630_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6659_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6668_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6677_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6680_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6686_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6692_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6695_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6700_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6704_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6708_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6713_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6716_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6720_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6722_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6731_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6732_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6736_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6740_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6749_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6763_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6769_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6772_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6781_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6785_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6787_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6790_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6793_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6799_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6800_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6808_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6817_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6826_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6832_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6835_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6841_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6844_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6848_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6853_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6857_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6866_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6878_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6881_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6883_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6884_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6889_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6896_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6902_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6905_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6914_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6920_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6928_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6929_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6932_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6937_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6938_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6947_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6950_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6953_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6961_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6964_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6969_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6974_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6977_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6985_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6992_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6993_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n6999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7001_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7009_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7017_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7018_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7042_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7054_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7058_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7066_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7081_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7082_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7090_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7114_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7126_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7130_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7139_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7153_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7154_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7166_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7169_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7172_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7177_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7178_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7184_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7190_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7193_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7202_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7208_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7216_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7218_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7220_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7226_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7234_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7235_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7238_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7243_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7244_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7250_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7255_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7258_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7267_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7275_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7279_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7280_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7291_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7299_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7303_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7307_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7313_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7316_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7319_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7322_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7323_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7325_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7328_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7331_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7334_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7337_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7340_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7343_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7346_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7347_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7349_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7352_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7355_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7358_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7361_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7363_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7364_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7367_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7370_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7371_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7373_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7376_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7379_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7382_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7385_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7388_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7391_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7394_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7397_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7400_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7403_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7406_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7407_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7410_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7419_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7425_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7427_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7437_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7443_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7446_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7452_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7455_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7470_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7491_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7500_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7510_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7534_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7540_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7552_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7558_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7564_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7570_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7576_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7582_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7588_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7600_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7606_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7612_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7630_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7660_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7700_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7708_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7720_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7732_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7736_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7760_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7763_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7772_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7781_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7787_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7790_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7799_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7800_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7808_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7810_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7826_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7832_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7835_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7844_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7848_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7853_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7860_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7866_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7878_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7883_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7884_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7896_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7902_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7910_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7914_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7920_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7928_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7932_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7938_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7947_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7950_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7960_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7964_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7974_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7992_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n7999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8007_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8010_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8017_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8030_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8054_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8060_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8078_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8081_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8102_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8110_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8126_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8139_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8151_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8153_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8160_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8165_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8166_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8169_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8172_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8177_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8184_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8190_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8192_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8193_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8204_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8208_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8216_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8220_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8230_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8235_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8238_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8243_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8244_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8255_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8260_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8267_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8279_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8280_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8303_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8310_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8313_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8316_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8319_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8322_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8325_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8328_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8334_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8337_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8340_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8343_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8346_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8349_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8352_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8358_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8360_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8361_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8364_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8367_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8370_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8373_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8376_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8377_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8382_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8385_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8388_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8391_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8394_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8397_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8400_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8406_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8407_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8410_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8413_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8416_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8422_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8425_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8428_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8431_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8434_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8437_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8440_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8446_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8449_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8452_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8455_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8458_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8461_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8464_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8470_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8473_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8476_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8479_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8482_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8485_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8488_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8494_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8497_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8500_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8508_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8510_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8512_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8516_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8524_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8530_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8532_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8548_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8556_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8572_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8580_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8596_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8604_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8620_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8628_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8630_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8636_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8644_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8652_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8659_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8660_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8668_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8676_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8677_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8680_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8684_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8686_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8692_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8695_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8704_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8708_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8710_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8713_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8716_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8720_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8722_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8724_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8731_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8732_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8740_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8748_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8749_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8756_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8760_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8766_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8769_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8775_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8778_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8784_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8785_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8787_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8793_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8796_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8800_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8802_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8805_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8810_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8811_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8814_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8820_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8823_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8829_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8832_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8838_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8841_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8847_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8848_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8850_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8857_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8860_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8863_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8866_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8869_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8872_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8875_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8878_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8881_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8883_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8884_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8887_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8890_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8893_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8896_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8899_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8902_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8905_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8908_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8910_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8911_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8914_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8917_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8920_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8923_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8926_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8928_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8932_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8935_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8937_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8938_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8941_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8944_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8947_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8950_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8953_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8960_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8961_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8969_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8977_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8992_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8993_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n8999_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9000_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9001_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9002_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9003_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9004_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9005_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9006_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9008_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9009_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9010_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9011_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9012_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9013_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9014_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9015_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9016_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9018_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9019_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9020_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9021_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9022_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9023_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9024_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9025_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9026_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9027_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9028_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9029_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9031_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9032_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9033_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9034_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9035_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9036_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9037_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9038_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9039_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9040_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9041_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9043_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9044_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9045_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9046_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9047_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9048_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9049_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9050_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9051_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9052_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9053_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9055_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9056_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9057_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9058_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9059_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9060_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9061_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9062_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9063_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9064_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9065_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9067_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9068_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9069_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9070_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9071_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9072_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9073_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9074_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9075_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9076_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9077_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9079_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9080_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9081_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9082_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9083_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9084_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9085_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9086_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9087_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9088_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9089_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9091_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9092_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9093_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9094_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9095_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9096_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9097_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9098_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9099_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9100_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9101_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9103_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9104_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9105_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9106_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9107_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9108_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9109_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9110_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9111_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9112_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9113_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9115_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9116_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9117_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9118_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9119_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9120_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9121_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9122_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9123_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9124_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9125_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9127_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9128_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9129_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9130_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9131_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9132_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9133_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9134_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9135_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9136_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9137_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9138_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9140_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9141_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9142_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9143_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9144_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9145_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9146_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9147_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9148_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9149_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9150_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9152_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9153_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9154_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9155_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9156_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9157_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9158_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9159_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9160_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9161_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9162_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9163_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9164_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9166_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9167_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9168_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9169_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9170_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9171_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9172_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9173_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9174_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9175_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9176_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9178_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9179_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9180_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9181_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9182_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9183_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9184_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9185_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9186_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9187_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9188_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9189_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9190_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9191_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9193_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9194_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9195_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9196_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9197_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9198_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9199_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9200_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9201_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9202_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9203_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9205_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9206_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9207_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9208_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9209_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9210_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9211_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9212_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9213_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9214_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9215_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9216_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9217_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9219_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9220_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9221_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9222_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9223_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9224_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9225_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9226_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9227_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9228_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9229_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9231_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9232_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9233_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9234_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9235_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9236_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9237_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9238_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9239_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9240_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9241_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9242_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9244_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9245_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9246_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9247_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9248_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9249_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9250_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9251_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9252_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9253_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9254_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9256_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9257_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9258_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9259_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9260_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9261_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9262_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9263_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9264_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9265_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9266_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9268_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9269_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9270_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9271_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9272_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9273_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9274_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9275_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9276_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9277_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9278_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9280_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9281_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9282_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9283_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9284_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9285_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9286_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9287_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9288_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9289_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9290_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9292_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9293_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9294_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9295_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9296_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9297_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9298_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9299_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9300_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9301_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9302_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9304_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9305_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9306_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9308_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9309_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9311_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9312_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9314_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9315_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9317_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9318_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9320_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9321_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9323_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9324_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9326_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9327_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9329_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9330_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9332_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9333_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9335_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9336_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9338_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9339_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9341_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9342_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9344_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9345_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9347_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9348_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9350_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9351_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9353_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9354_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9356_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9357_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9359_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9360_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9362_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9363_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9365_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9366_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9368_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9369_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9371_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9372_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9374_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9375_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9377_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9378_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9380_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9381_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9383_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9384_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9386_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9387_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9389_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9390_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9392_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9393_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9395_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9396_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9398_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9399_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9401_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9402_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9403_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9404_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9405_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9406_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9408_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9409_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9411_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9412_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9414_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9415_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9417_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9418_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9420_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9421_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9423_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9424_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9426_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9427_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9429_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9430_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9432_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9433_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9435_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9436_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9438_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9439_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9441_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9442_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9444_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9445_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9447_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9448_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9450_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9451_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9453_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9454_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9456_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9457_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9459_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9460_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9462_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9463_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9465_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9466_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9468_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9469_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9471_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9472_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9474_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9475_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9477_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9478_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9480_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9481_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9483_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9484_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9486_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9487_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9489_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9490_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9492_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9493_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9495_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9496_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9498_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9499_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9501_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9502_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9503_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9504_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9505_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9506_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9507_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9509_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9510_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9511_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9512_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9513_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9514_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9515_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9517_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9518_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9519_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9520_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9521_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9522_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9523_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9525_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9526_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9527_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9528_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9529_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9530_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9531_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9533_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9534_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9535_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9536_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9537_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9538_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9539_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9541_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9542_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9543_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9544_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9545_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9546_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9547_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9549_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9550_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9551_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9552_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9553_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9554_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9555_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9557_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9558_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9559_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9560_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9561_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9562_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9563_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9565_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9566_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9567_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9568_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9569_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9570_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9571_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9573_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9574_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9575_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9576_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9577_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9578_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9579_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9581_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9582_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9583_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9584_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9585_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9586_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9587_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9589_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9590_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9591_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9592_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9593_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9594_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9595_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9597_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9598_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9599_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9600_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9601_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9602_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9603_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9605_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9606_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9607_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9608_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9609_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9610_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9611_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9613_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9614_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9615_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9616_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9617_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9618_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9619_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9621_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9622_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9623_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9624_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9625_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9626_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9627_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9629_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9630_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9631_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9632_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9633_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9634_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9635_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9637_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9638_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9639_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9640_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9641_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9642_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9643_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9645_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9646_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9647_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9648_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9649_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9650_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9651_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9653_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9654_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9655_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9656_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9657_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9658_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9659_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9661_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9662_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9663_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9664_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9665_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9666_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9667_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9669_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9670_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9671_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9672_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9673_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9674_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9675_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9677_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9678_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9679_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9680_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9681_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9682_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9683_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9685_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9686_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9687_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9688_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9689_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9690_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9691_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9693_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9694_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9695_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9696_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9697_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9698_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9699_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9701_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9702_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9703_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9704_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9705_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9706_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9707_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9709_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9710_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9711_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9712_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9713_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9714_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9715_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9717_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9718_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9719_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9720_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9721_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9722_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9723_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9725_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9726_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9727_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9728_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9729_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9730_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9731_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9733_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9734_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9735_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9736_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9737_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9738_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9739_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9741_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9742_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9743_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9744_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9745_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9746_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9747_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9749_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9750_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9751_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9752_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9753_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9754_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9755_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9757_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9758_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9759_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9761_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9762_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9764_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9765_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9767_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9768_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9770_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9771_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9773_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9774_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9776_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9777_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9779_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9780_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9782_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9783_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9785_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9786_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9788_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9789_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9791_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9792_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9794_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9795_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9797_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9798_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9800_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9801_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9803_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9804_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9806_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9807_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9809_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9810_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9812_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9813_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9815_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9816_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9818_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9819_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9821_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9822_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9824_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9825_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9827_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9828_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9830_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9831_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9833_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9834_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9836_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9837_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9839_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9840_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9842_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9843_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9845_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9846_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9848_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9849_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9851_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9852_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9854_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9855_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9856_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9857_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9858_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9859_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9861_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9862_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9864_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9865_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9867_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9868_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9870_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9871_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9873_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9874_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9876_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9877_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9879_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9880_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9882_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9883_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9885_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9886_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9888_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9889_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9891_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9892_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9894_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9895_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9897_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9898_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9900_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9901_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9903_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9904_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9906_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9907_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9909_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9910_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9912_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9913_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9915_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9916_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9918_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9919_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9921_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9922_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9924_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9925_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9927_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9928_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9930_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9931_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9933_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9934_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9936_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9937_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9939_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9940_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9942_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9943_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9945_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9946_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9948_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9949_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9951_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9952_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9954_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9955_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9956_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9957_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9958_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9959_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9960_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9962_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9963_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9964_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9965_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9966_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9967_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9968_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9970_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9971_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9972_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9973_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9974_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9975_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9976_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9978_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9979_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9980_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9981_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9982_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9983_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9984_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9986_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9987_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9988_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9989_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9990_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9991_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9992_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9994_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9995_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9996_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9997_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9998_; 
wire AES_CORE_DATAPATH__abc_16009_new_n9999_; 
wire AES_CORE_DATAPATH_bkp_0__0_; 
wire AES_CORE_DATAPATH_bkp_0__10_; 
wire AES_CORE_DATAPATH_bkp_0__11_; 
wire AES_CORE_DATAPATH_bkp_0__12_; 
wire AES_CORE_DATAPATH_bkp_0__13_; 
wire AES_CORE_DATAPATH_bkp_0__14_; 
wire AES_CORE_DATAPATH_bkp_0__15_; 
wire AES_CORE_DATAPATH_bkp_0__16_; 
wire AES_CORE_DATAPATH_bkp_0__17_; 
wire AES_CORE_DATAPATH_bkp_0__18_; 
wire AES_CORE_DATAPATH_bkp_0__19_; 
wire AES_CORE_DATAPATH_bkp_0__1_; 
wire AES_CORE_DATAPATH_bkp_0__20_; 
wire AES_CORE_DATAPATH_bkp_0__21_; 
wire AES_CORE_DATAPATH_bkp_0__22_; 
wire AES_CORE_DATAPATH_bkp_0__23_; 
wire AES_CORE_DATAPATH_bkp_0__24_; 
wire AES_CORE_DATAPATH_bkp_0__25_; 
wire AES_CORE_DATAPATH_bkp_0__26_; 
wire AES_CORE_DATAPATH_bkp_0__27_; 
wire AES_CORE_DATAPATH_bkp_0__28_; 
wire AES_CORE_DATAPATH_bkp_0__29_; 
wire AES_CORE_DATAPATH_bkp_0__2_; 
wire AES_CORE_DATAPATH_bkp_0__30_; 
wire AES_CORE_DATAPATH_bkp_0__31_; 
wire AES_CORE_DATAPATH_bkp_0__3_; 
wire AES_CORE_DATAPATH_bkp_0__4_; 
wire AES_CORE_DATAPATH_bkp_0__5_; 
wire AES_CORE_DATAPATH_bkp_0__6_; 
wire AES_CORE_DATAPATH_bkp_0__7_; 
wire AES_CORE_DATAPATH_bkp_0__8_; 
wire AES_CORE_DATAPATH_bkp_0__9_; 
wire AES_CORE_DATAPATH_bkp_1_0__0_; 
wire AES_CORE_DATAPATH_bkp_1_0__10_; 
wire AES_CORE_DATAPATH_bkp_1_0__11_; 
wire AES_CORE_DATAPATH_bkp_1_0__12_; 
wire AES_CORE_DATAPATH_bkp_1_0__13_; 
wire AES_CORE_DATAPATH_bkp_1_0__14_; 
wire AES_CORE_DATAPATH_bkp_1_0__15_; 
wire AES_CORE_DATAPATH_bkp_1_0__16_; 
wire AES_CORE_DATAPATH_bkp_1_0__17_; 
wire AES_CORE_DATAPATH_bkp_1_0__18_; 
wire AES_CORE_DATAPATH_bkp_1_0__19_; 
wire AES_CORE_DATAPATH_bkp_1_0__1_; 
wire AES_CORE_DATAPATH_bkp_1_0__20_; 
wire AES_CORE_DATAPATH_bkp_1_0__21_; 
wire AES_CORE_DATAPATH_bkp_1_0__22_; 
wire AES_CORE_DATAPATH_bkp_1_0__23_; 
wire AES_CORE_DATAPATH_bkp_1_0__24_; 
wire AES_CORE_DATAPATH_bkp_1_0__25_; 
wire AES_CORE_DATAPATH_bkp_1_0__26_; 
wire AES_CORE_DATAPATH_bkp_1_0__27_; 
wire AES_CORE_DATAPATH_bkp_1_0__28_; 
wire AES_CORE_DATAPATH_bkp_1_0__29_; 
wire AES_CORE_DATAPATH_bkp_1_0__2_; 
wire AES_CORE_DATAPATH_bkp_1_0__30_; 
wire AES_CORE_DATAPATH_bkp_1_0__31_; 
wire AES_CORE_DATAPATH_bkp_1_0__3_; 
wire AES_CORE_DATAPATH_bkp_1_0__4_; 
wire AES_CORE_DATAPATH_bkp_1_0__5_; 
wire AES_CORE_DATAPATH_bkp_1_0__6_; 
wire AES_CORE_DATAPATH_bkp_1_0__7_; 
wire AES_CORE_DATAPATH_bkp_1_0__8_; 
wire AES_CORE_DATAPATH_bkp_1_0__9_; 
wire AES_CORE_DATAPATH_bkp_1_1__0_; 
wire AES_CORE_DATAPATH_bkp_1_1__10_; 
wire AES_CORE_DATAPATH_bkp_1_1__11_; 
wire AES_CORE_DATAPATH_bkp_1_1__12_; 
wire AES_CORE_DATAPATH_bkp_1_1__13_; 
wire AES_CORE_DATAPATH_bkp_1_1__14_; 
wire AES_CORE_DATAPATH_bkp_1_1__15_; 
wire AES_CORE_DATAPATH_bkp_1_1__16_; 
wire AES_CORE_DATAPATH_bkp_1_1__17_; 
wire AES_CORE_DATAPATH_bkp_1_1__18_; 
wire AES_CORE_DATAPATH_bkp_1_1__19_; 
wire AES_CORE_DATAPATH_bkp_1_1__1_; 
wire AES_CORE_DATAPATH_bkp_1_1__20_; 
wire AES_CORE_DATAPATH_bkp_1_1__21_; 
wire AES_CORE_DATAPATH_bkp_1_1__22_; 
wire AES_CORE_DATAPATH_bkp_1_1__23_; 
wire AES_CORE_DATAPATH_bkp_1_1__24_; 
wire AES_CORE_DATAPATH_bkp_1_1__25_; 
wire AES_CORE_DATAPATH_bkp_1_1__26_; 
wire AES_CORE_DATAPATH_bkp_1_1__27_; 
wire AES_CORE_DATAPATH_bkp_1_1__28_; 
wire AES_CORE_DATAPATH_bkp_1_1__29_; 
wire AES_CORE_DATAPATH_bkp_1_1__2_; 
wire AES_CORE_DATAPATH_bkp_1_1__30_; 
wire AES_CORE_DATAPATH_bkp_1_1__31_; 
wire AES_CORE_DATAPATH_bkp_1_1__3_; 
wire AES_CORE_DATAPATH_bkp_1_1__4_; 
wire AES_CORE_DATAPATH_bkp_1_1__5_; 
wire AES_CORE_DATAPATH_bkp_1_1__6_; 
wire AES_CORE_DATAPATH_bkp_1_1__7_; 
wire AES_CORE_DATAPATH_bkp_1_1__8_; 
wire AES_CORE_DATAPATH_bkp_1_1__9_; 
wire AES_CORE_DATAPATH_bkp_1_2__0_; 
wire AES_CORE_DATAPATH_bkp_1_2__10_; 
wire AES_CORE_DATAPATH_bkp_1_2__11_; 
wire AES_CORE_DATAPATH_bkp_1_2__12_; 
wire AES_CORE_DATAPATH_bkp_1_2__13_; 
wire AES_CORE_DATAPATH_bkp_1_2__14_; 
wire AES_CORE_DATAPATH_bkp_1_2__15_; 
wire AES_CORE_DATAPATH_bkp_1_2__16_; 
wire AES_CORE_DATAPATH_bkp_1_2__17_; 
wire AES_CORE_DATAPATH_bkp_1_2__18_; 
wire AES_CORE_DATAPATH_bkp_1_2__19_; 
wire AES_CORE_DATAPATH_bkp_1_2__1_; 
wire AES_CORE_DATAPATH_bkp_1_2__20_; 
wire AES_CORE_DATAPATH_bkp_1_2__21_; 
wire AES_CORE_DATAPATH_bkp_1_2__22_; 
wire AES_CORE_DATAPATH_bkp_1_2__23_; 
wire AES_CORE_DATAPATH_bkp_1_2__24_; 
wire AES_CORE_DATAPATH_bkp_1_2__25_; 
wire AES_CORE_DATAPATH_bkp_1_2__26_; 
wire AES_CORE_DATAPATH_bkp_1_2__27_; 
wire AES_CORE_DATAPATH_bkp_1_2__28_; 
wire AES_CORE_DATAPATH_bkp_1_2__29_; 
wire AES_CORE_DATAPATH_bkp_1_2__2_; 
wire AES_CORE_DATAPATH_bkp_1_2__30_; 
wire AES_CORE_DATAPATH_bkp_1_2__31_; 
wire AES_CORE_DATAPATH_bkp_1_2__3_; 
wire AES_CORE_DATAPATH_bkp_1_2__4_; 
wire AES_CORE_DATAPATH_bkp_1_2__5_; 
wire AES_CORE_DATAPATH_bkp_1_2__6_; 
wire AES_CORE_DATAPATH_bkp_1_2__7_; 
wire AES_CORE_DATAPATH_bkp_1_2__8_; 
wire AES_CORE_DATAPATH_bkp_1_2__9_; 
wire AES_CORE_DATAPATH_bkp_1_3__0_; 
wire AES_CORE_DATAPATH_bkp_1_3__10_; 
wire AES_CORE_DATAPATH_bkp_1_3__11_; 
wire AES_CORE_DATAPATH_bkp_1_3__12_; 
wire AES_CORE_DATAPATH_bkp_1_3__13_; 
wire AES_CORE_DATAPATH_bkp_1_3__14_; 
wire AES_CORE_DATAPATH_bkp_1_3__15_; 
wire AES_CORE_DATAPATH_bkp_1_3__16_; 
wire AES_CORE_DATAPATH_bkp_1_3__17_; 
wire AES_CORE_DATAPATH_bkp_1_3__18_; 
wire AES_CORE_DATAPATH_bkp_1_3__19_; 
wire AES_CORE_DATAPATH_bkp_1_3__1_; 
wire AES_CORE_DATAPATH_bkp_1_3__20_; 
wire AES_CORE_DATAPATH_bkp_1_3__21_; 
wire AES_CORE_DATAPATH_bkp_1_3__22_; 
wire AES_CORE_DATAPATH_bkp_1_3__23_; 
wire AES_CORE_DATAPATH_bkp_1_3__24_; 
wire AES_CORE_DATAPATH_bkp_1_3__25_; 
wire AES_CORE_DATAPATH_bkp_1_3__26_; 
wire AES_CORE_DATAPATH_bkp_1_3__27_; 
wire AES_CORE_DATAPATH_bkp_1_3__28_; 
wire AES_CORE_DATAPATH_bkp_1_3__29_; 
wire AES_CORE_DATAPATH_bkp_1_3__2_; 
wire AES_CORE_DATAPATH_bkp_1_3__30_; 
wire AES_CORE_DATAPATH_bkp_1_3__31_; 
wire AES_CORE_DATAPATH_bkp_1_3__3_; 
wire AES_CORE_DATAPATH_bkp_1_3__4_; 
wire AES_CORE_DATAPATH_bkp_1_3__5_; 
wire AES_CORE_DATAPATH_bkp_1_3__6_; 
wire AES_CORE_DATAPATH_bkp_1_3__7_; 
wire AES_CORE_DATAPATH_bkp_1_3__8_; 
wire AES_CORE_DATAPATH_bkp_1_3__9_; 
wire AES_CORE_DATAPATH_bkp_1__0_; 
wire AES_CORE_DATAPATH_bkp_1__10_; 
wire AES_CORE_DATAPATH_bkp_1__11_; 
wire AES_CORE_DATAPATH_bkp_1__12_; 
wire AES_CORE_DATAPATH_bkp_1__13_; 
wire AES_CORE_DATAPATH_bkp_1__14_; 
wire AES_CORE_DATAPATH_bkp_1__15_; 
wire AES_CORE_DATAPATH_bkp_1__16_; 
wire AES_CORE_DATAPATH_bkp_1__17_; 
wire AES_CORE_DATAPATH_bkp_1__18_; 
wire AES_CORE_DATAPATH_bkp_1__19_; 
wire AES_CORE_DATAPATH_bkp_1__1_; 
wire AES_CORE_DATAPATH_bkp_1__20_; 
wire AES_CORE_DATAPATH_bkp_1__21_; 
wire AES_CORE_DATAPATH_bkp_1__22_; 
wire AES_CORE_DATAPATH_bkp_1__23_; 
wire AES_CORE_DATAPATH_bkp_1__24_; 
wire AES_CORE_DATAPATH_bkp_1__25_; 
wire AES_CORE_DATAPATH_bkp_1__26_; 
wire AES_CORE_DATAPATH_bkp_1__27_; 
wire AES_CORE_DATAPATH_bkp_1__28_; 
wire AES_CORE_DATAPATH_bkp_1__29_; 
wire AES_CORE_DATAPATH_bkp_1__2_; 
wire AES_CORE_DATAPATH_bkp_1__30_; 
wire AES_CORE_DATAPATH_bkp_1__31_; 
wire AES_CORE_DATAPATH_bkp_1__3_; 
wire AES_CORE_DATAPATH_bkp_1__4_; 
wire AES_CORE_DATAPATH_bkp_1__5_; 
wire AES_CORE_DATAPATH_bkp_1__6_; 
wire AES_CORE_DATAPATH_bkp_1__7_; 
wire AES_CORE_DATAPATH_bkp_1__8_; 
wire AES_CORE_DATAPATH_bkp_1__9_; 
wire AES_CORE_DATAPATH_bkp_2__0_; 
wire AES_CORE_DATAPATH_bkp_2__10_; 
wire AES_CORE_DATAPATH_bkp_2__11_; 
wire AES_CORE_DATAPATH_bkp_2__12_; 
wire AES_CORE_DATAPATH_bkp_2__13_; 
wire AES_CORE_DATAPATH_bkp_2__14_; 
wire AES_CORE_DATAPATH_bkp_2__15_; 
wire AES_CORE_DATAPATH_bkp_2__16_; 
wire AES_CORE_DATAPATH_bkp_2__17_; 
wire AES_CORE_DATAPATH_bkp_2__18_; 
wire AES_CORE_DATAPATH_bkp_2__19_; 
wire AES_CORE_DATAPATH_bkp_2__1_; 
wire AES_CORE_DATAPATH_bkp_2__20_; 
wire AES_CORE_DATAPATH_bkp_2__21_; 
wire AES_CORE_DATAPATH_bkp_2__22_; 
wire AES_CORE_DATAPATH_bkp_2__23_; 
wire AES_CORE_DATAPATH_bkp_2__24_; 
wire AES_CORE_DATAPATH_bkp_2__25_; 
wire AES_CORE_DATAPATH_bkp_2__26_; 
wire AES_CORE_DATAPATH_bkp_2__27_; 
wire AES_CORE_DATAPATH_bkp_2__28_; 
wire AES_CORE_DATAPATH_bkp_2__29_; 
wire AES_CORE_DATAPATH_bkp_2__2_; 
wire AES_CORE_DATAPATH_bkp_2__30_; 
wire AES_CORE_DATAPATH_bkp_2__31_; 
wire AES_CORE_DATAPATH_bkp_2__3_; 
wire AES_CORE_DATAPATH_bkp_2__4_; 
wire AES_CORE_DATAPATH_bkp_2__5_; 
wire AES_CORE_DATAPATH_bkp_2__6_; 
wire AES_CORE_DATAPATH_bkp_2__7_; 
wire AES_CORE_DATAPATH_bkp_2__8_; 
wire AES_CORE_DATAPATH_bkp_2__9_; 
wire AES_CORE_DATAPATH_bkp_3__0_; 
wire AES_CORE_DATAPATH_bkp_3__10_; 
wire AES_CORE_DATAPATH_bkp_3__11_; 
wire AES_CORE_DATAPATH_bkp_3__12_; 
wire AES_CORE_DATAPATH_bkp_3__13_; 
wire AES_CORE_DATAPATH_bkp_3__14_; 
wire AES_CORE_DATAPATH_bkp_3__15_; 
wire AES_CORE_DATAPATH_bkp_3__16_; 
wire AES_CORE_DATAPATH_bkp_3__17_; 
wire AES_CORE_DATAPATH_bkp_3__18_; 
wire AES_CORE_DATAPATH_bkp_3__19_; 
wire AES_CORE_DATAPATH_bkp_3__1_; 
wire AES_CORE_DATAPATH_bkp_3__20_; 
wire AES_CORE_DATAPATH_bkp_3__21_; 
wire AES_CORE_DATAPATH_bkp_3__22_; 
wire AES_CORE_DATAPATH_bkp_3__23_; 
wire AES_CORE_DATAPATH_bkp_3__24_; 
wire AES_CORE_DATAPATH_bkp_3__25_; 
wire AES_CORE_DATAPATH_bkp_3__26_; 
wire AES_CORE_DATAPATH_bkp_3__27_; 
wire AES_CORE_DATAPATH_bkp_3__28_; 
wire AES_CORE_DATAPATH_bkp_3__29_; 
wire AES_CORE_DATAPATH_bkp_3__2_; 
wire AES_CORE_DATAPATH_bkp_3__30_; 
wire AES_CORE_DATAPATH_bkp_3__31_; 
wire AES_CORE_DATAPATH_bkp_3__3_; 
wire AES_CORE_DATAPATH_bkp_3__4_; 
wire AES_CORE_DATAPATH_bkp_3__5_; 
wire AES_CORE_DATAPATH_bkp_3__6_; 
wire AES_CORE_DATAPATH_bkp_3__7_; 
wire AES_CORE_DATAPATH_bkp_3__8_; 
wire AES_CORE_DATAPATH_bkp_3__9_; 
wire AES_CORE_DATAPATH_col_0__0_; 
wire AES_CORE_DATAPATH_col_0__10_; 
wire AES_CORE_DATAPATH_col_0__11_; 
wire AES_CORE_DATAPATH_col_0__12_; 
wire AES_CORE_DATAPATH_col_0__13_; 
wire AES_CORE_DATAPATH_col_0__14_; 
wire AES_CORE_DATAPATH_col_0__15_; 
wire AES_CORE_DATAPATH_col_0__16_; 
wire AES_CORE_DATAPATH_col_0__17_; 
wire AES_CORE_DATAPATH_col_0__18_; 
wire AES_CORE_DATAPATH_col_0__19_; 
wire AES_CORE_DATAPATH_col_0__1_; 
wire AES_CORE_DATAPATH_col_0__20_; 
wire AES_CORE_DATAPATH_col_0__21_; 
wire AES_CORE_DATAPATH_col_0__22_; 
wire AES_CORE_DATAPATH_col_0__23_; 
wire AES_CORE_DATAPATH_col_0__24_; 
wire AES_CORE_DATAPATH_col_0__25_; 
wire AES_CORE_DATAPATH_col_0__26_; 
wire AES_CORE_DATAPATH_col_0__27_; 
wire AES_CORE_DATAPATH_col_0__28_; 
wire AES_CORE_DATAPATH_col_0__29_; 
wire AES_CORE_DATAPATH_col_0__2_; 
wire AES_CORE_DATAPATH_col_0__30_; 
wire AES_CORE_DATAPATH_col_0__31_; 
wire AES_CORE_DATAPATH_col_0__3_; 
wire AES_CORE_DATAPATH_col_0__4_; 
wire AES_CORE_DATAPATH_col_0__5_; 
wire AES_CORE_DATAPATH_col_0__6_; 
wire AES_CORE_DATAPATH_col_0__7_; 
wire AES_CORE_DATAPATH_col_0__8_; 
wire AES_CORE_DATAPATH_col_0__9_; 
wire AES_CORE_DATAPATH_col_3__0_; 
wire AES_CORE_DATAPATH_col_3__10_; 
wire AES_CORE_DATAPATH_col_3__11_; 
wire AES_CORE_DATAPATH_col_3__12_; 
wire AES_CORE_DATAPATH_col_3__13_; 
wire AES_CORE_DATAPATH_col_3__14_; 
wire AES_CORE_DATAPATH_col_3__15_; 
wire AES_CORE_DATAPATH_col_3__16_; 
wire AES_CORE_DATAPATH_col_3__17_; 
wire AES_CORE_DATAPATH_col_3__18_; 
wire AES_CORE_DATAPATH_col_3__19_; 
wire AES_CORE_DATAPATH_col_3__1_; 
wire AES_CORE_DATAPATH_col_3__20_; 
wire AES_CORE_DATAPATH_col_3__21_; 
wire AES_CORE_DATAPATH_col_3__22_; 
wire AES_CORE_DATAPATH_col_3__23_; 
wire AES_CORE_DATAPATH_col_3__24_; 
wire AES_CORE_DATAPATH_col_3__25_; 
wire AES_CORE_DATAPATH_col_3__26_; 
wire AES_CORE_DATAPATH_col_3__27_; 
wire AES_CORE_DATAPATH_col_3__28_; 
wire AES_CORE_DATAPATH_col_3__29_; 
wire AES_CORE_DATAPATH_col_3__2_; 
wire AES_CORE_DATAPATH_col_3__30_; 
wire AES_CORE_DATAPATH_col_3__31_; 
wire AES_CORE_DATAPATH_col_3__3_; 
wire AES_CORE_DATAPATH_col_3__4_; 
wire AES_CORE_DATAPATH_col_3__5_; 
wire AES_CORE_DATAPATH_col_3__6_; 
wire AES_CORE_DATAPATH_col_3__7_; 
wire AES_CORE_DATAPATH_col_3__8_; 
wire AES_CORE_DATAPATH_col_3__9_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_; 
wire AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_; 
wire AES_CORE_DATAPATH_col_en_host_0_; 
wire AES_CORE_DATAPATH_col_en_host_1_; 
wire AES_CORE_DATAPATH_col_en_host_2_; 
wire AES_CORE_DATAPATH_col_en_host_3_; 
wire AES_CORE_DATAPATH_col_sel_host_0_; 
wire AES_CORE_DATAPATH_col_sel_host_1_; 
wire AES_CORE_DATAPATH_col_sel_pp1_0_; 
wire AES_CORE_DATAPATH_col_sel_pp1_1_; 
wire AES_CORE_DATAPATH_col_sel_pp2_0_; 
wire AES_CORE_DATAPATH_col_sel_pp2_1_; 
wire AES_CORE_DATAPATH_iv_0__0_; 
wire AES_CORE_DATAPATH_iv_0__10_; 
wire AES_CORE_DATAPATH_iv_0__11_; 
wire AES_CORE_DATAPATH_iv_0__12_; 
wire AES_CORE_DATAPATH_iv_0__13_; 
wire AES_CORE_DATAPATH_iv_0__14_; 
wire AES_CORE_DATAPATH_iv_0__15_; 
wire AES_CORE_DATAPATH_iv_0__16_; 
wire AES_CORE_DATAPATH_iv_0__17_; 
wire AES_CORE_DATAPATH_iv_0__18_; 
wire AES_CORE_DATAPATH_iv_0__19_; 
wire AES_CORE_DATAPATH_iv_0__1_; 
wire AES_CORE_DATAPATH_iv_0__20_; 
wire AES_CORE_DATAPATH_iv_0__21_; 
wire AES_CORE_DATAPATH_iv_0__22_; 
wire AES_CORE_DATAPATH_iv_0__23_; 
wire AES_CORE_DATAPATH_iv_0__24_; 
wire AES_CORE_DATAPATH_iv_0__25_; 
wire AES_CORE_DATAPATH_iv_0__26_; 
wire AES_CORE_DATAPATH_iv_0__27_; 
wire AES_CORE_DATAPATH_iv_0__28_; 
wire AES_CORE_DATAPATH_iv_0__29_; 
wire AES_CORE_DATAPATH_iv_0__2_; 
wire AES_CORE_DATAPATH_iv_0__30_; 
wire AES_CORE_DATAPATH_iv_0__31_; 
wire AES_CORE_DATAPATH_iv_0__3_; 
wire AES_CORE_DATAPATH_iv_0__4_; 
wire AES_CORE_DATAPATH_iv_0__5_; 
wire AES_CORE_DATAPATH_iv_0__6_; 
wire AES_CORE_DATAPATH_iv_0__7_; 
wire AES_CORE_DATAPATH_iv_0__8_; 
wire AES_CORE_DATAPATH_iv_0__9_; 
wire AES_CORE_DATAPATH_iv_1__0_; 
wire AES_CORE_DATAPATH_iv_1__10_; 
wire AES_CORE_DATAPATH_iv_1__11_; 
wire AES_CORE_DATAPATH_iv_1__12_; 
wire AES_CORE_DATAPATH_iv_1__13_; 
wire AES_CORE_DATAPATH_iv_1__14_; 
wire AES_CORE_DATAPATH_iv_1__15_; 
wire AES_CORE_DATAPATH_iv_1__16_; 
wire AES_CORE_DATAPATH_iv_1__17_; 
wire AES_CORE_DATAPATH_iv_1__18_; 
wire AES_CORE_DATAPATH_iv_1__19_; 
wire AES_CORE_DATAPATH_iv_1__1_; 
wire AES_CORE_DATAPATH_iv_1__20_; 
wire AES_CORE_DATAPATH_iv_1__21_; 
wire AES_CORE_DATAPATH_iv_1__22_; 
wire AES_CORE_DATAPATH_iv_1__23_; 
wire AES_CORE_DATAPATH_iv_1__24_; 
wire AES_CORE_DATAPATH_iv_1__25_; 
wire AES_CORE_DATAPATH_iv_1__26_; 
wire AES_CORE_DATAPATH_iv_1__27_; 
wire AES_CORE_DATAPATH_iv_1__28_; 
wire AES_CORE_DATAPATH_iv_1__29_; 
wire AES_CORE_DATAPATH_iv_1__2_; 
wire AES_CORE_DATAPATH_iv_1__30_; 
wire AES_CORE_DATAPATH_iv_1__31_; 
wire AES_CORE_DATAPATH_iv_1__3_; 
wire AES_CORE_DATAPATH_iv_1__4_; 
wire AES_CORE_DATAPATH_iv_1__5_; 
wire AES_CORE_DATAPATH_iv_1__6_; 
wire AES_CORE_DATAPATH_iv_1__7_; 
wire AES_CORE_DATAPATH_iv_1__8_; 
wire AES_CORE_DATAPATH_iv_1__9_; 
wire AES_CORE_DATAPATH_iv_2__0_; 
wire AES_CORE_DATAPATH_iv_2__10_; 
wire AES_CORE_DATAPATH_iv_2__11_; 
wire AES_CORE_DATAPATH_iv_2__12_; 
wire AES_CORE_DATAPATH_iv_2__13_; 
wire AES_CORE_DATAPATH_iv_2__14_; 
wire AES_CORE_DATAPATH_iv_2__15_; 
wire AES_CORE_DATAPATH_iv_2__16_; 
wire AES_CORE_DATAPATH_iv_2__17_; 
wire AES_CORE_DATAPATH_iv_2__18_; 
wire AES_CORE_DATAPATH_iv_2__19_; 
wire AES_CORE_DATAPATH_iv_2__1_; 
wire AES_CORE_DATAPATH_iv_2__20_; 
wire AES_CORE_DATAPATH_iv_2__21_; 
wire AES_CORE_DATAPATH_iv_2__22_; 
wire AES_CORE_DATAPATH_iv_2__23_; 
wire AES_CORE_DATAPATH_iv_2__24_; 
wire AES_CORE_DATAPATH_iv_2__25_; 
wire AES_CORE_DATAPATH_iv_2__26_; 
wire AES_CORE_DATAPATH_iv_2__27_; 
wire AES_CORE_DATAPATH_iv_2__28_; 
wire AES_CORE_DATAPATH_iv_2__29_; 
wire AES_CORE_DATAPATH_iv_2__2_; 
wire AES_CORE_DATAPATH_iv_2__30_; 
wire AES_CORE_DATAPATH_iv_2__31_; 
wire AES_CORE_DATAPATH_iv_2__3_; 
wire AES_CORE_DATAPATH_iv_2__4_; 
wire AES_CORE_DATAPATH_iv_2__5_; 
wire AES_CORE_DATAPATH_iv_2__6_; 
wire AES_CORE_DATAPATH_iv_2__7_; 
wire AES_CORE_DATAPATH_iv_2__8_; 
wire AES_CORE_DATAPATH_iv_2__9_; 
wire AES_CORE_DATAPATH_iv_3__0_; 
wire AES_CORE_DATAPATH_iv_3__10_; 
wire AES_CORE_DATAPATH_iv_3__11_; 
wire AES_CORE_DATAPATH_iv_3__12_; 
wire AES_CORE_DATAPATH_iv_3__13_; 
wire AES_CORE_DATAPATH_iv_3__14_; 
wire AES_CORE_DATAPATH_iv_3__15_; 
wire AES_CORE_DATAPATH_iv_3__16_; 
wire AES_CORE_DATAPATH_iv_3__17_; 
wire AES_CORE_DATAPATH_iv_3__18_; 
wire AES_CORE_DATAPATH_iv_3__19_; 
wire AES_CORE_DATAPATH_iv_3__1_; 
wire AES_CORE_DATAPATH_iv_3__20_; 
wire AES_CORE_DATAPATH_iv_3__21_; 
wire AES_CORE_DATAPATH_iv_3__22_; 
wire AES_CORE_DATAPATH_iv_3__23_; 
wire AES_CORE_DATAPATH_iv_3__24_; 
wire AES_CORE_DATAPATH_iv_3__25_; 
wire AES_CORE_DATAPATH_iv_3__26_; 
wire AES_CORE_DATAPATH_iv_3__27_; 
wire AES_CORE_DATAPATH_iv_3__28_; 
wire AES_CORE_DATAPATH_iv_3__29_; 
wire AES_CORE_DATAPATH_iv_3__2_; 
wire AES_CORE_DATAPATH_iv_3__30_; 
wire AES_CORE_DATAPATH_iv_3__31_; 
wire AES_CORE_DATAPATH_iv_3__3_; 
wire AES_CORE_DATAPATH_iv_3__4_; 
wire AES_CORE_DATAPATH_iv_3__5_; 
wire AES_CORE_DATAPATH_iv_3__6_; 
wire AES_CORE_DATAPATH_iv_3__7_; 
wire AES_CORE_DATAPATH_iv_3__8_; 
wire AES_CORE_DATAPATH_iv_3__9_; 
wire AES_CORE_DATAPATH_key_en_pp1_0_; 
wire AES_CORE_DATAPATH_key_en_pp1_1_; 
wire AES_CORE_DATAPATH_key_en_pp1_2_; 
wire AES_CORE_DATAPATH_key_en_pp1_3_; 
wire AES_CORE_DATAPATH_key_host_0__0_; 
wire AES_CORE_DATAPATH_key_host_0__10_; 
wire AES_CORE_DATAPATH_key_host_0__11_; 
wire AES_CORE_DATAPATH_key_host_0__12_; 
wire AES_CORE_DATAPATH_key_host_0__13_; 
wire AES_CORE_DATAPATH_key_host_0__14_; 
wire AES_CORE_DATAPATH_key_host_0__15_; 
wire AES_CORE_DATAPATH_key_host_0__16_; 
wire AES_CORE_DATAPATH_key_host_0__17_; 
wire AES_CORE_DATAPATH_key_host_0__18_; 
wire AES_CORE_DATAPATH_key_host_0__19_; 
wire AES_CORE_DATAPATH_key_host_0__1_; 
wire AES_CORE_DATAPATH_key_host_0__20_; 
wire AES_CORE_DATAPATH_key_host_0__21_; 
wire AES_CORE_DATAPATH_key_host_0__22_; 
wire AES_CORE_DATAPATH_key_host_0__23_; 
wire AES_CORE_DATAPATH_key_host_0__24_; 
wire AES_CORE_DATAPATH_key_host_0__25_; 
wire AES_CORE_DATAPATH_key_host_0__26_; 
wire AES_CORE_DATAPATH_key_host_0__27_; 
wire AES_CORE_DATAPATH_key_host_0__28_; 
wire AES_CORE_DATAPATH_key_host_0__29_; 
wire AES_CORE_DATAPATH_key_host_0__2_; 
wire AES_CORE_DATAPATH_key_host_0__30_; 
wire AES_CORE_DATAPATH_key_host_0__31_; 
wire AES_CORE_DATAPATH_key_host_0__3_; 
wire AES_CORE_DATAPATH_key_host_0__4_; 
wire AES_CORE_DATAPATH_key_host_0__5_; 
wire AES_CORE_DATAPATH_key_host_0__6_; 
wire AES_CORE_DATAPATH_key_host_0__7_; 
wire AES_CORE_DATAPATH_key_host_0__8_; 
wire AES_CORE_DATAPATH_key_host_0__9_; 
wire AES_CORE_DATAPATH_key_host_1__0_; 
wire AES_CORE_DATAPATH_key_host_1__10_; 
wire AES_CORE_DATAPATH_key_host_1__11_; 
wire AES_CORE_DATAPATH_key_host_1__12_; 
wire AES_CORE_DATAPATH_key_host_1__13_; 
wire AES_CORE_DATAPATH_key_host_1__14_; 
wire AES_CORE_DATAPATH_key_host_1__15_; 
wire AES_CORE_DATAPATH_key_host_1__16_; 
wire AES_CORE_DATAPATH_key_host_1__17_; 
wire AES_CORE_DATAPATH_key_host_1__18_; 
wire AES_CORE_DATAPATH_key_host_1__19_; 
wire AES_CORE_DATAPATH_key_host_1__1_; 
wire AES_CORE_DATAPATH_key_host_1__20_; 
wire AES_CORE_DATAPATH_key_host_1__21_; 
wire AES_CORE_DATAPATH_key_host_1__22_; 
wire AES_CORE_DATAPATH_key_host_1__23_; 
wire AES_CORE_DATAPATH_key_host_1__24_; 
wire AES_CORE_DATAPATH_key_host_1__25_; 
wire AES_CORE_DATAPATH_key_host_1__26_; 
wire AES_CORE_DATAPATH_key_host_1__27_; 
wire AES_CORE_DATAPATH_key_host_1__28_; 
wire AES_CORE_DATAPATH_key_host_1__29_; 
wire AES_CORE_DATAPATH_key_host_1__2_; 
wire AES_CORE_DATAPATH_key_host_1__30_; 
wire AES_CORE_DATAPATH_key_host_1__31_; 
wire AES_CORE_DATAPATH_key_host_1__3_; 
wire AES_CORE_DATAPATH_key_host_1__4_; 
wire AES_CORE_DATAPATH_key_host_1__5_; 
wire AES_CORE_DATAPATH_key_host_1__6_; 
wire AES_CORE_DATAPATH_key_host_1__7_; 
wire AES_CORE_DATAPATH_key_host_1__8_; 
wire AES_CORE_DATAPATH_key_host_1__9_; 
wire AES_CORE_DATAPATH_key_host_2__0_; 
wire AES_CORE_DATAPATH_key_host_2__10_; 
wire AES_CORE_DATAPATH_key_host_2__11_; 
wire AES_CORE_DATAPATH_key_host_2__12_; 
wire AES_CORE_DATAPATH_key_host_2__13_; 
wire AES_CORE_DATAPATH_key_host_2__14_; 
wire AES_CORE_DATAPATH_key_host_2__15_; 
wire AES_CORE_DATAPATH_key_host_2__16_; 
wire AES_CORE_DATAPATH_key_host_2__17_; 
wire AES_CORE_DATAPATH_key_host_2__18_; 
wire AES_CORE_DATAPATH_key_host_2__19_; 
wire AES_CORE_DATAPATH_key_host_2__1_; 
wire AES_CORE_DATAPATH_key_host_2__20_; 
wire AES_CORE_DATAPATH_key_host_2__21_; 
wire AES_CORE_DATAPATH_key_host_2__22_; 
wire AES_CORE_DATAPATH_key_host_2__23_; 
wire AES_CORE_DATAPATH_key_host_2__24_; 
wire AES_CORE_DATAPATH_key_host_2__25_; 
wire AES_CORE_DATAPATH_key_host_2__26_; 
wire AES_CORE_DATAPATH_key_host_2__27_; 
wire AES_CORE_DATAPATH_key_host_2__28_; 
wire AES_CORE_DATAPATH_key_host_2__29_; 
wire AES_CORE_DATAPATH_key_host_2__2_; 
wire AES_CORE_DATAPATH_key_host_2__30_; 
wire AES_CORE_DATAPATH_key_host_2__31_; 
wire AES_CORE_DATAPATH_key_host_2__3_; 
wire AES_CORE_DATAPATH_key_host_2__4_; 
wire AES_CORE_DATAPATH_key_host_2__5_; 
wire AES_CORE_DATAPATH_key_host_2__6_; 
wire AES_CORE_DATAPATH_key_host_2__7_; 
wire AES_CORE_DATAPATH_key_host_2__8_; 
wire AES_CORE_DATAPATH_key_host_2__9_; 
wire AES_CORE_DATAPATH_key_host_3__0_; 
wire AES_CORE_DATAPATH_key_host_3__10_; 
wire AES_CORE_DATAPATH_key_host_3__11_; 
wire AES_CORE_DATAPATH_key_host_3__12_; 
wire AES_CORE_DATAPATH_key_host_3__13_; 
wire AES_CORE_DATAPATH_key_host_3__14_; 
wire AES_CORE_DATAPATH_key_host_3__15_; 
wire AES_CORE_DATAPATH_key_host_3__16_; 
wire AES_CORE_DATAPATH_key_host_3__17_; 
wire AES_CORE_DATAPATH_key_host_3__18_; 
wire AES_CORE_DATAPATH_key_host_3__19_; 
wire AES_CORE_DATAPATH_key_host_3__1_; 
wire AES_CORE_DATAPATH_key_host_3__20_; 
wire AES_CORE_DATAPATH_key_host_3__21_; 
wire AES_CORE_DATAPATH_key_host_3__22_; 
wire AES_CORE_DATAPATH_key_host_3__23_; 
wire AES_CORE_DATAPATH_key_host_3__24_; 
wire AES_CORE_DATAPATH_key_host_3__25_; 
wire AES_CORE_DATAPATH_key_host_3__26_; 
wire AES_CORE_DATAPATH_key_host_3__27_; 
wire AES_CORE_DATAPATH_key_host_3__28_; 
wire AES_CORE_DATAPATH_key_host_3__29_; 
wire AES_CORE_DATAPATH_key_host_3__2_; 
wire AES_CORE_DATAPATH_key_host_3__30_; 
wire AES_CORE_DATAPATH_key_host_3__31_; 
wire AES_CORE_DATAPATH_key_host_3__3_; 
wire AES_CORE_DATAPATH_key_host_3__4_; 
wire AES_CORE_DATAPATH_key_host_3__5_; 
wire AES_CORE_DATAPATH_key_host_3__6_; 
wire AES_CORE_DATAPATH_key_host_3__7_; 
wire AES_CORE_DATAPATH_key_host_3__8_; 
wire AES_CORE_DATAPATH_key_host_3__9_; 
wire AES_CORE_DATAPATH_key_out_sel_pp1_0_; 
wire AES_CORE_DATAPATH_key_out_sel_pp1_1_; 
wire AES_CORE_DATAPATH_key_out_sel_pp2_0_; 
wire AES_CORE_DATAPATH_key_out_sel_pp2_1_; 
wire AES_CORE_DATAPATH_key_sel_pp1; 
wire AES_CORE_DATAPATH_last_round_pp1; 
wire AES_CORE_DATAPATH_last_round_pp2; 
wire AES_CORE_DATAPATH_rk_out_sel; 
wire AES_CORE_DATAPATH_rk_out_sel_pp1; 
wire AES_CORE_DATAPATH_rk_out_sel_pp2; 
wire AES_CORE_DATAPATH_rk_sel_pp1_0_; 
wire AES_CORE_DATAPATH_rk_sel_pp1_1_; 
wire AES_CORE_DATAPATH_rk_sel_pp2_0_; 
wire AES_CORE_DATAPATH_rk_sel_pp2_1_; 
wire _abc_15574_new_n11_; 
wire _abc_15574_new_n12_; 
wire _abc_15574_new_n13_; 
wire _abc_15574_new_n15_; 
input \addr[0] ;
input \addr[1] ;
input \aes_mode[0] ;
input \aes_mode[1] ;
input \bus_in[0] ;
input \bus_in[10] ;
input \bus_in[11] ;
input \bus_in[12] ;
input \bus_in[13] ;
input \bus_in[14] ;
input \bus_in[15] ;
input \bus_in[16] ;
input \bus_in[17] ;
input \bus_in[18] ;
input \bus_in[19] ;
input \bus_in[1] ;
input \bus_in[20] ;
input \bus_in[21] ;
input \bus_in[22] ;
input \bus_in[23] ;
input \bus_in[24] ;
input \bus_in[25] ;
input \bus_in[26] ;
input \bus_in[27] ;
input \bus_in[28] ;
input \bus_in[29] ;
input \bus_in[2] ;
input \bus_in[30] ;
input \bus_in[31] ;
input \bus_in[3] ;
input \bus_in[4] ;
input \bus_in[5] ;
input \bus_in[6] ;
input \bus_in[7] ;
input \bus_in[8] ;
input \bus_in[9] ;
input clk;
output \col_out[0] ;
output \col_out[10] ;
output \col_out[11] ;
output \col_out[12] ;
output \col_out[13] ;
output \col_out[14] ;
output \col_out[15] ;
output \col_out[16] ;
output \col_out[17] ;
output \col_out[18] ;
output \col_out[19] ;
output \col_out[1] ;
output \col_out[20] ;
output \col_out[21] ;
output \col_out[22] ;
output \col_out[23] ;
output \col_out[24] ;
output \col_out[25] ;
output \col_out[26] ;
output \col_out[27] ;
output \col_out[28] ;
output \col_out[29] ;
output \col_out[2] ;
output \col_out[30] ;
output \col_out[31] ;
output \col_out[3] ;
output \col_out[4] ;
output \col_out[5] ;
output \col_out[6] ;
output \col_out[7] ;
output \col_out[8] ;
output \col_out[9] ;
input \data_type[0] ;
input \data_type[1] ;
input disable_core;
output end_aes;
input first_block;
input \iv_en[0] ;
input \iv_en[1] ;
input \iv_en[2] ;
input \iv_en[3] ;
output \iv_out[0] ;
output \iv_out[10] ;
output \iv_out[11] ;
output \iv_out[12] ;
output \iv_out[13] ;
output \iv_out[14] ;
output \iv_out[15] ;
output \iv_out[16] ;
output \iv_out[17] ;
output \iv_out[18] ;
output \iv_out[19] ;
output \iv_out[1] ;
output \iv_out[20] ;
output \iv_out[21] ;
output \iv_out[22] ;
output \iv_out[23] ;
output \iv_out[24] ;
output \iv_out[25] ;
output \iv_out[26] ;
output \iv_out[27] ;
output \iv_out[28] ;
output \iv_out[29] ;
output \iv_out[2] ;
output \iv_out[30] ;
output \iv_out[31] ;
output \iv_out[3] ;
output \iv_out[4] ;
output \iv_out[5] ;
output \iv_out[6] ;
output \iv_out[7] ;
output \iv_out[8] ;
output \iv_out[9] ;
input \iv_sel_rd[0] ;
input \iv_sel_rd[1] ;
input \iv_sel_rd[2] ;
input \iv_sel_rd[3] ;
input \key_en[0] ;
input \key_en[1] ;
input \key_en[2] ;
input \key_en[3] ;
output \key_out[0] ;
output \key_out[10] ;
output \key_out[11] ;
output \key_out[12] ;
output \key_out[13] ;
output \key_out[14] ;
output \key_out[15] ;
output \key_out[16] ;
output \key_out[17] ;
output \key_out[18] ;
output \key_out[19] ;
output \key_out[1] ;
output \key_out[20] ;
output \key_out[21] ;
output \key_out[22] ;
output \key_out[23] ;
output \key_out[24] ;
output \key_out[25] ;
output \key_out[26] ;
output \key_out[27] ;
output \key_out[28] ;
output \key_out[29] ;
output \key_out[2] ;
output \key_out[30] ;
output \key_out[31] ;
output \key_out[3] ;
output \key_out[4] ;
output \key_out[5] ;
output \key_out[6] ;
output \key_out[7] ;
output \key_out[8] ;
output \key_out[9] ;
input \key_sel_rd[0] ;
input \key_sel_rd[1] ;
input \op_mode[0] ;
input \op_mode[1] ;
input read_en;
input rst_n;
input start;
input write_en;
AND2X2 AND2X2_1 ( .A(_abc_15574_new_n12_), .B(write_en), .Y(_abc_15574_new_n13_));
AND2X2 AND2X2_10 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n77_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n78_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n79_));
AND2X2 AND2X2_100 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n211_), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT_iv_cnt_en));
AND2X2 AND2X2_1000 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4463_));
AND2X2 AND2X2_1001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3496_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4464_));
AND2X2 AND2X2_1002 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4466_));
AND2X2 AND2X2_1003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3528_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4467_));
AND2X2 AND2X2_1004 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4469_));
AND2X2 AND2X2_1005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3560_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4470_));
AND2X2 AND2X2_1006 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4472_));
AND2X2 AND2X2_1007 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3592_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4473_));
AND2X2 AND2X2_1008 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4475_));
AND2X2 AND2X2_1009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3624_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4476_));
AND2X2 AND2X2_101 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1817));
AND2X2 AND2X2_1010 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4478_));
AND2X2 AND2X2_1011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3656_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4479_));
AND2X2 AND2X2_1012 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4481_));
AND2X2 AND2X2_1013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3688_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4482_));
AND2X2 AND2X2_1014 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4484_));
AND2X2 AND2X2_1015 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3720_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4485_));
AND2X2 AND2X2_1016 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4487_));
AND2X2 AND2X2_1017 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3752_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4488_));
AND2X2 AND2X2_1018 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4490_));
AND2X2 AND2X2_1019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3784_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4491_));
AND2X2 AND2X2_102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2458_));
AND2X2 AND2X2_1020 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4493_));
AND2X2 AND2X2_1021 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3816_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4494_));
AND2X2 AND2X2_1022 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4496_));
AND2X2 AND2X2_1023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3848_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4497_));
AND2X2 AND2X2_1024 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4499_));
AND2X2 AND2X2_1025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3880_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4500_));
AND2X2 AND2X2_1026 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4502_));
AND2X2 AND2X2_1027 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3912_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4503_));
AND2X2 AND2X2_1028 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4505_));
AND2X2 AND2X2_1029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3944_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4506_));
AND2X2 AND2X2_103 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2459_));
AND2X2 AND2X2_1030 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4508_));
AND2X2 AND2X2_1031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3976_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4509_));
AND2X2 AND2X2_1032 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4511_));
AND2X2 AND2X2_1033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4008_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4512_));
AND2X2 AND2X2_1034 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4514_));
AND2X2 AND2X2_1035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4040_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4515_));
AND2X2 AND2X2_1036 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4517_));
AND2X2 AND2X2_1037 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4072_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4518_));
AND2X2 AND2X2_1038 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4520_));
AND2X2 AND2X2_1039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4104_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4521_));
AND2X2 AND2X2_104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2463_));
AND2X2 AND2X2_1040 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4523_));
AND2X2 AND2X2_1041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4136_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4524_));
AND2X2 AND2X2_1042 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4526_));
AND2X2 AND2X2_1043 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4168_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4527_));
AND2X2 AND2X2_1044 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4529_));
AND2X2 AND2X2_1045 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4200_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4530_));
AND2X2 AND2X2_1046 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4532_));
AND2X2 AND2X2_1047 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4232_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4533_));
AND2X2 AND2X2_1048 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4535_));
AND2X2 AND2X2_1049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4264_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4536_));
AND2X2 AND2X2_105 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2464_));
AND2X2 AND2X2_1050 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4538_));
AND2X2 AND2X2_1051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4296_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4539_));
AND2X2 AND2X2_1052 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4541_));
AND2X2 AND2X2_1053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4328_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4542_));
AND2X2 AND2X2_1054 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4544_));
AND2X2 AND2X2_1055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4360_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4545_));
AND2X2 AND2X2_1056 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4547_));
AND2X2 AND2X2_1057 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4392_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4548_));
AND2X2 AND2X2_1058 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4550_));
AND2X2 AND2X2_1059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4424_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4551_));
AND2X2 AND2X2_106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2468_));
AND2X2 AND2X2_1060 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4553_));
AND2X2 AND2X2_1061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4456_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4554_));
AND2X2 AND2X2_1062 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4557_));
AND2X2 AND2X2_1063 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4558_));
AND2X2 AND2X2_1064 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4561_), .B(AES_CORE_DATAPATH__abc_16009_new_n4562_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4563_));
AND2X2 AND2X2_1065 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4560_), .B(AES_CORE_DATAPATH__abc_16009_new_n4563_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4564_));
AND2X2 AND2X2_1066 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_sel_pp1), .Y(AES_CORE_DATAPATH__abc_16009_new_n4565_));
AND2X2 AND2X2_1067 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_sel), .Y(AES_CORE_DATAPATH__abc_16009_new_n4566_));
AND2X2 AND2X2_1068 ( .A(\key_en[1] ), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4568_));
AND2X2 AND2X2_1069 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4569_));
AND2X2 AND2X2_107 ( .A(AES_CORE_CONTROL_UNIT_col_en_0_), .B(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_DATAPATH__abc_16009_new_n2469_));
AND2X2 AND2X2_1070 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4573_), .B(AES_CORE_DATAPATH__abc_16009_new_n4571_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4574_));
AND2X2 AND2X2_1071 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4575_), .B(AES_CORE_DATAPATH__abc_16009_new_n4577_), .Y(AES_CORE_DATAPATH__0key_1__31_0__0_));
AND2X2 AND2X2_1072 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4580_));
AND2X2 AND2X2_1073 ( .A(\key_en[1] ), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4581_));
AND2X2 AND2X2_1074 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4579_), .B(AES_CORE_DATAPATH__abc_16009_new_n4583_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4584_));
AND2X2 AND2X2_1075 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4584_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4585_));
AND2X2 AND2X2_1076 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4586_));
AND2X2 AND2X2_1077 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4589_));
AND2X2 AND2X2_1078 ( .A(\key_en[1] ), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4590_));
AND2X2 AND2X2_1079 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4588_), .B(AES_CORE_DATAPATH__abc_16009_new_n4592_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4593_));
AND2X2 AND2X2_108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2473_));
AND2X2 AND2X2_1080 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4593_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4594_));
AND2X2 AND2X2_1081 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4595_));
AND2X2 AND2X2_1082 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4598_));
AND2X2 AND2X2_1083 ( .A(\key_en[1] ), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4599_));
AND2X2 AND2X2_1084 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4597_), .B(AES_CORE_DATAPATH__abc_16009_new_n4601_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4602_));
AND2X2 AND2X2_1085 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4602_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4603_));
AND2X2 AND2X2_1086 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4604_));
AND2X2 AND2X2_1087 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4607_));
AND2X2 AND2X2_1088 ( .A(\key_en[1] ), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4608_));
AND2X2 AND2X2_1089 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4606_), .B(AES_CORE_DATAPATH__abc_16009_new_n4610_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4611_));
AND2X2 AND2X2_109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2474_), .B(AES_CORE_DATAPATH__abc_16009_new_n2476_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2477_));
AND2X2 AND2X2_1090 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4611_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4612_));
AND2X2 AND2X2_1091 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4613_));
AND2X2 AND2X2_1092 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4616_));
AND2X2 AND2X2_1093 ( .A(\key_en[1] ), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4617_));
AND2X2 AND2X2_1094 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4615_), .B(AES_CORE_DATAPATH__abc_16009_new_n4619_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4620_));
AND2X2 AND2X2_1095 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4620_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4621_));
AND2X2 AND2X2_1096 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4622_));
AND2X2 AND2X2_1097 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4625_));
AND2X2 AND2X2_1098 ( .A(\key_en[1] ), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4626_));
AND2X2 AND2X2_1099 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4624_), .B(AES_CORE_DATAPATH__abc_16009_new_n4628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4629_));
AND2X2 AND2X2_11 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n80_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n81_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_));
AND2X2 AND2X2_110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2479_));
AND2X2 AND2X2_1100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4629_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4630_));
AND2X2 AND2X2_1101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4631_));
AND2X2 AND2X2_1102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4634_));
AND2X2 AND2X2_1103 ( .A(\key_en[1] ), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4635_));
AND2X2 AND2X2_1104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4633_), .B(AES_CORE_DATAPATH__abc_16009_new_n4637_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4638_));
AND2X2 AND2X2_1105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4639_), .B(AES_CORE_DATAPATH__abc_16009_new_n4640_), .Y(AES_CORE_DATAPATH__0key_1__31_0__7_));
AND2X2 AND2X2_1106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4643_));
AND2X2 AND2X2_1107 ( .A(\key_en[1] ), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4644_));
AND2X2 AND2X2_1108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4642_), .B(AES_CORE_DATAPATH__abc_16009_new_n4646_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4647_));
AND2X2 AND2X2_1109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4647_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4648_));
AND2X2 AND2X2_111 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2480_));
AND2X2 AND2X2_1110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4649_));
AND2X2 AND2X2_1111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4652_));
AND2X2 AND2X2_1112 ( .A(\key_en[1] ), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4653_));
AND2X2 AND2X2_1113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4651_), .B(AES_CORE_DATAPATH__abc_16009_new_n4655_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4656_));
AND2X2 AND2X2_1114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4656_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4657_));
AND2X2 AND2X2_1115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4658_));
AND2X2 AND2X2_1116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4661_));
AND2X2 AND2X2_1117 ( .A(\key_en[1] ), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4662_));
AND2X2 AND2X2_1118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4660_), .B(AES_CORE_DATAPATH__abc_16009_new_n4664_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4665_));
AND2X2 AND2X2_1119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4666_), .B(AES_CORE_DATAPATH__abc_16009_new_n4667_), .Y(AES_CORE_DATAPATH__0key_1__31_0__10_));
AND2X2 AND2X2_112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2486_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2487_));
AND2X2 AND2X2_1120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4670_));
AND2X2 AND2X2_1121 ( .A(\key_en[1] ), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4671_));
AND2X2 AND2X2_1122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4669_), .B(AES_CORE_DATAPATH__abc_16009_new_n4673_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4674_));
AND2X2 AND2X2_1123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4675_), .B(AES_CORE_DATAPATH__abc_16009_new_n4676_), .Y(AES_CORE_DATAPATH__0key_1__31_0__11_));
AND2X2 AND2X2_1124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4679_));
AND2X2 AND2X2_1125 ( .A(\key_en[1] ), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4680_));
AND2X2 AND2X2_1126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4678_), .B(AES_CORE_DATAPATH__abc_16009_new_n4682_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4683_));
AND2X2 AND2X2_1127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4684_), .B(AES_CORE_DATAPATH__abc_16009_new_n4685_), .Y(AES_CORE_DATAPATH__0key_1__31_0__12_));
AND2X2 AND2X2_1128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4688_));
AND2X2 AND2X2_1129 ( .A(\key_en[1] ), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4689_));
AND2X2 AND2X2_113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2478_), .B(AES_CORE_DATAPATH__abc_16009_new_n2487_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2488_));
AND2X2 AND2X2_1130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4687_), .B(AES_CORE_DATAPATH__abc_16009_new_n4691_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4692_));
AND2X2 AND2X2_1131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4693_), .B(AES_CORE_DATAPATH__abc_16009_new_n4694_), .Y(AES_CORE_DATAPATH__0key_1__31_0__13_));
AND2X2 AND2X2_1132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4697_));
AND2X2 AND2X2_1133 ( .A(\key_en[1] ), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4698_));
AND2X2 AND2X2_1134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4696_), .B(AES_CORE_DATAPATH__abc_16009_new_n4700_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4701_));
AND2X2 AND2X2_1135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4701_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4702_));
AND2X2 AND2X2_1136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4703_));
AND2X2 AND2X2_1137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4706_));
AND2X2 AND2X2_1138 ( .A(\key_en[1] ), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4707_));
AND2X2 AND2X2_1139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4705_), .B(AES_CORE_DATAPATH__abc_16009_new_n4709_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4710_));
AND2X2 AND2X2_114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2489_));
AND2X2 AND2X2_1140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4710_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4711_));
AND2X2 AND2X2_1141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4712_));
AND2X2 AND2X2_1142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4715_));
AND2X2 AND2X2_1143 ( .A(\key_en[1] ), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4716_));
AND2X2 AND2X2_1144 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4714_), .B(AES_CORE_DATAPATH__abc_16009_new_n4718_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4719_));
AND2X2 AND2X2_1145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4720_), .B(AES_CORE_DATAPATH__abc_16009_new_n4721_), .Y(AES_CORE_DATAPATH__0key_1__31_0__16_));
AND2X2 AND2X2_1146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4724_));
AND2X2 AND2X2_1147 ( .A(\key_en[1] ), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4725_));
AND2X2 AND2X2_1148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4723_), .B(AES_CORE_DATAPATH__abc_16009_new_n4727_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4728_));
AND2X2 AND2X2_1149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4729_), .B(AES_CORE_DATAPATH__abc_16009_new_n4730_), .Y(AES_CORE_DATAPATH__0key_1__31_0__17_));
AND2X2 AND2X2_115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2491_));
AND2X2 AND2X2_1150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4733_));
AND2X2 AND2X2_1151 ( .A(\key_en[1] ), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4734_));
AND2X2 AND2X2_1152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4732_), .B(AES_CORE_DATAPATH__abc_16009_new_n4736_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4737_));
AND2X2 AND2X2_1153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4738_), .B(AES_CORE_DATAPATH__abc_16009_new_n4739_), .Y(AES_CORE_DATAPATH__0key_1__31_0__18_));
AND2X2 AND2X2_1154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4742_));
AND2X2 AND2X2_1155 ( .A(\key_en[1] ), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4743_));
AND2X2 AND2X2_1156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4741_), .B(AES_CORE_DATAPATH__abc_16009_new_n4745_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4746_));
AND2X2 AND2X2_1157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4746_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4747_));
AND2X2 AND2X2_1158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4748_));
AND2X2 AND2X2_1159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4751_));
AND2X2 AND2X2_116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2491_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2492_));
AND2X2 AND2X2_1160 ( .A(\key_en[1] ), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4752_));
AND2X2 AND2X2_1161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4750_), .B(AES_CORE_DATAPATH__abc_16009_new_n4754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4755_));
AND2X2 AND2X2_1162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4755_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4756_));
AND2X2 AND2X2_1163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4757_));
AND2X2 AND2X2_1164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4760_));
AND2X2 AND2X2_1165 ( .A(\key_en[1] ), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4761_));
AND2X2 AND2X2_1166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4759_), .B(AES_CORE_DATAPATH__abc_16009_new_n4763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4764_));
AND2X2 AND2X2_1167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4764_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4765_));
AND2X2 AND2X2_1168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4766_));
AND2X2 AND2X2_1169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4769_));
AND2X2 AND2X2_117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2493_));
AND2X2 AND2X2_1170 ( .A(\key_en[1] ), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4770_));
AND2X2 AND2X2_1171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4768_), .B(AES_CORE_DATAPATH__abc_16009_new_n4772_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4773_));
AND2X2 AND2X2_1172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4774_), .B(AES_CORE_DATAPATH__abc_16009_new_n4775_), .Y(AES_CORE_DATAPATH__0key_1__31_0__22_));
AND2X2 AND2X2_1173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4778_));
AND2X2 AND2X2_1174 ( .A(\key_en[1] ), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4779_));
AND2X2 AND2X2_1175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4777_), .B(AES_CORE_DATAPATH__abc_16009_new_n4781_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4782_));
AND2X2 AND2X2_1176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4782_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4783_));
AND2X2 AND2X2_1177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4784_));
AND2X2 AND2X2_1178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4787_));
AND2X2 AND2X2_1179 ( .A(\key_en[1] ), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4788_));
AND2X2 AND2X2_118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2496_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2497_));
AND2X2 AND2X2_1180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4786_), .B(AES_CORE_DATAPATH__abc_16009_new_n4790_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4791_));
AND2X2 AND2X2_1181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4792_), .B(AES_CORE_DATAPATH__abc_16009_new_n4793_), .Y(AES_CORE_DATAPATH__0key_1__31_0__24_));
AND2X2 AND2X2_1182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4796_));
AND2X2 AND2X2_1183 ( .A(\key_en[1] ), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4797_));
AND2X2 AND2X2_1184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4795_), .B(AES_CORE_DATAPATH__abc_16009_new_n4799_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4800_));
AND2X2 AND2X2_1185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4800_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4801_));
AND2X2 AND2X2_1186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4802_));
AND2X2 AND2X2_1187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4805_));
AND2X2 AND2X2_1188 ( .A(\key_en[1] ), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4806_));
AND2X2 AND2X2_1189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4804_), .B(AES_CORE_DATAPATH__abc_16009_new_n4808_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4809_));
AND2X2 AND2X2_119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2495_), .B(AES_CORE_DATAPATH__abc_16009_new_n2497_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2498_));
AND2X2 AND2X2_1190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4810_), .B(AES_CORE_DATAPATH__abc_16009_new_n4811_), .Y(AES_CORE_DATAPATH__0key_1__31_0__26_));
AND2X2 AND2X2_1191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4814_));
AND2X2 AND2X2_1192 ( .A(\key_en[1] ), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4815_));
AND2X2 AND2X2_1193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4813_), .B(AES_CORE_DATAPATH__abc_16009_new_n4817_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4818_));
AND2X2 AND2X2_1194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4818_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4819_));
AND2X2 AND2X2_1195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4820_));
AND2X2 AND2X2_1196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4823_));
AND2X2 AND2X2_1197 ( .A(\key_en[1] ), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4824_));
AND2X2 AND2X2_1198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4822_), .B(AES_CORE_DATAPATH__abc_16009_new_n4826_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4827_));
AND2X2 AND2X2_1199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4828_), .B(AES_CORE_DATAPATH__abc_16009_new_n4829_), .Y(AES_CORE_DATAPATH__0key_1__31_0__28_));
AND2X2 AND2X2_12 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n79_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n82_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n83_));
AND2X2 AND2X2_120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2499_));
AND2X2 AND2X2_1200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4832_));
AND2X2 AND2X2_1201 ( .A(\key_en[1] ), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4833_));
AND2X2 AND2X2_1202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4831_), .B(AES_CORE_DATAPATH__abc_16009_new_n4835_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4836_));
AND2X2 AND2X2_1203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4836_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4837_));
AND2X2 AND2X2_1204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4838_));
AND2X2 AND2X2_1205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4841_));
AND2X2 AND2X2_1206 ( .A(\key_en[1] ), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4842_));
AND2X2 AND2X2_1207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4840_), .B(AES_CORE_DATAPATH__abc_16009_new_n4844_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4845_));
AND2X2 AND2X2_1208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4846_), .B(AES_CORE_DATAPATH__abc_16009_new_n4847_), .Y(AES_CORE_DATAPATH__0key_1__31_0__30_));
AND2X2 AND2X2_1209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4562_), .B(AES_CORE_DATAPATH_key_host_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4849_));
AND2X2 AND2X2_121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2501_));
AND2X2 AND2X2_1210 ( .A(\key_en[1] ), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4850_));
AND2X2 AND2X2_1211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4853_), .B(AES_CORE_DATAPATH__abc_16009_new_n4852_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4854_));
AND2X2 AND2X2_1212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4854_), .B(AES_CORE_DATAPATH__abc_16009_new_n4576_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4855_));
AND2X2 AND2X2_1213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4856_));
AND2X2 AND2X2_1214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4858_));
AND2X2 AND2X2_1215 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4859_));
AND2X2 AND2X2_1216 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4561_), .B(AES_CORE_DATAPATH__abc_16009_new_n4862_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4863_));
AND2X2 AND2X2_1217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4861_), .B(AES_CORE_DATAPATH__abc_16009_new_n4863_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4864_));
AND2X2 AND2X2_1218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4866_));
AND2X2 AND2X2_1219 ( .A(\bus_in[0] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4867_));
AND2X2 AND2X2_122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2501_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2502_));
AND2X2 AND2X2_1220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4868_));
AND2X2 AND2X2_1221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH__abc_16009_new_n4869_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4870_));
AND2X2 AND2X2_1222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4871_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4872_));
AND2X2 AND2X2_1223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4873_));
AND2X2 AND2X2_1224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4876_));
AND2X2 AND2X2_1225 ( .A(\bus_in[1] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4877_));
AND2X2 AND2X2_1226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4875_), .B(AES_CORE_DATAPATH__abc_16009_new_n4879_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4880_));
AND2X2 AND2X2_1227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4880_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4881_));
AND2X2 AND2X2_1228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4882_));
AND2X2 AND2X2_1229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4885_));
AND2X2 AND2X2_123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2503_));
AND2X2 AND2X2_1230 ( .A(\bus_in[2] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4886_));
AND2X2 AND2X2_1231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4884_), .B(AES_CORE_DATAPATH__abc_16009_new_n4888_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4889_));
AND2X2 AND2X2_1232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4889_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4890_));
AND2X2 AND2X2_1233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4891_));
AND2X2 AND2X2_1234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4894_));
AND2X2 AND2X2_1235 ( .A(\bus_in[3] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4895_));
AND2X2 AND2X2_1236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4893_), .B(AES_CORE_DATAPATH__abc_16009_new_n4897_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4898_));
AND2X2 AND2X2_1237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4898_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4899_));
AND2X2 AND2X2_1238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4900_));
AND2X2 AND2X2_1239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4903_));
AND2X2 AND2X2_124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2506_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2507_));
AND2X2 AND2X2_1240 ( .A(\bus_in[4] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4904_));
AND2X2 AND2X2_1241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4902_), .B(AES_CORE_DATAPATH__abc_16009_new_n4906_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4907_));
AND2X2 AND2X2_1242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4908_), .B(AES_CORE_DATAPATH__abc_16009_new_n4909_), .Y(AES_CORE_DATAPATH__0key_0__31_0__4_));
AND2X2 AND2X2_1243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4912_));
AND2X2 AND2X2_1244 ( .A(\bus_in[5] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4913_));
AND2X2 AND2X2_1245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4911_), .B(AES_CORE_DATAPATH__abc_16009_new_n4915_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4916_));
AND2X2 AND2X2_1246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4916_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4917_));
AND2X2 AND2X2_1247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4918_));
AND2X2 AND2X2_1248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4921_));
AND2X2 AND2X2_1249 ( .A(\bus_in[6] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4922_));
AND2X2 AND2X2_125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2505_), .B(AES_CORE_DATAPATH__abc_16009_new_n2507_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2508_));
AND2X2 AND2X2_1250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4920_), .B(AES_CORE_DATAPATH__abc_16009_new_n4924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4925_));
AND2X2 AND2X2_1251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4926_), .B(AES_CORE_DATAPATH__abc_16009_new_n4927_), .Y(AES_CORE_DATAPATH__0key_0__31_0__6_));
AND2X2 AND2X2_1252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4930_));
AND2X2 AND2X2_1253 ( .A(\bus_in[7] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4931_));
AND2X2 AND2X2_1254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4929_), .B(AES_CORE_DATAPATH__abc_16009_new_n4933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4934_));
AND2X2 AND2X2_1255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4934_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4935_));
AND2X2 AND2X2_1256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4936_));
AND2X2 AND2X2_1257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4939_));
AND2X2 AND2X2_1258 ( .A(\bus_in[8] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4940_));
AND2X2 AND2X2_1259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4938_), .B(AES_CORE_DATAPATH__abc_16009_new_n4942_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4943_));
AND2X2 AND2X2_126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2509_));
AND2X2 AND2X2_1260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4943_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4944_));
AND2X2 AND2X2_1261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4945_));
AND2X2 AND2X2_1262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4948_));
AND2X2 AND2X2_1263 ( .A(\bus_in[9] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4949_));
AND2X2 AND2X2_1264 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4947_), .B(AES_CORE_DATAPATH__abc_16009_new_n4951_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4952_));
AND2X2 AND2X2_1265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4953_), .B(AES_CORE_DATAPATH__abc_16009_new_n4954_), .Y(AES_CORE_DATAPATH__0key_0__31_0__9_));
AND2X2 AND2X2_1266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4957_));
AND2X2 AND2X2_1267 ( .A(\bus_in[10] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4958_));
AND2X2 AND2X2_1268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4956_), .B(AES_CORE_DATAPATH__abc_16009_new_n4960_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4961_));
AND2X2 AND2X2_1269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4961_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4962_));
AND2X2 AND2X2_127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2511_));
AND2X2 AND2X2_1270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4963_));
AND2X2 AND2X2_1271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4966_));
AND2X2 AND2X2_1272 ( .A(\bus_in[11] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4967_));
AND2X2 AND2X2_1273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4965_), .B(AES_CORE_DATAPATH__abc_16009_new_n4969_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4970_));
AND2X2 AND2X2_1274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4970_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4971_));
AND2X2 AND2X2_1275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4972_));
AND2X2 AND2X2_1276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4975_));
AND2X2 AND2X2_1277 ( .A(\bus_in[12] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4976_));
AND2X2 AND2X2_1278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4974_), .B(AES_CORE_DATAPATH__abc_16009_new_n4978_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4979_));
AND2X2 AND2X2_1279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4979_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4980_));
AND2X2 AND2X2_128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2511_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2512_));
AND2X2 AND2X2_1280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4981_));
AND2X2 AND2X2_1281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4984_));
AND2X2 AND2X2_1282 ( .A(\bus_in[13] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4985_));
AND2X2 AND2X2_1283 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4983_), .B(AES_CORE_DATAPATH__abc_16009_new_n4987_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4988_));
AND2X2 AND2X2_1284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4989_), .B(AES_CORE_DATAPATH__abc_16009_new_n4990_), .Y(AES_CORE_DATAPATH__0key_0__31_0__13_));
AND2X2 AND2X2_1285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4993_));
AND2X2 AND2X2_1286 ( .A(\bus_in[14] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4994_));
AND2X2 AND2X2_1287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4992_), .B(AES_CORE_DATAPATH__abc_16009_new_n4996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4997_));
AND2X2 AND2X2_1288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4997_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4998_));
AND2X2 AND2X2_1289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4999_));
AND2X2 AND2X2_129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2513_));
AND2X2 AND2X2_1290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5002_));
AND2X2 AND2X2_1291 ( .A(\bus_in[15] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5003_));
AND2X2 AND2X2_1292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5001_), .B(AES_CORE_DATAPATH__abc_16009_new_n5005_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5006_));
AND2X2 AND2X2_1293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5006_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5007_));
AND2X2 AND2X2_1294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5008_));
AND2X2 AND2X2_1295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5011_));
AND2X2 AND2X2_1296 ( .A(\bus_in[16] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5012_));
AND2X2 AND2X2_1297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5010_), .B(AES_CORE_DATAPATH__abc_16009_new_n5014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5015_));
AND2X2 AND2X2_1298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5015_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5016_));
AND2X2 AND2X2_1299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5017_));
AND2X2 AND2X2_13 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n83_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_));
AND2X2 AND2X2_130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2516_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2517_));
AND2X2 AND2X2_1300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5020_));
AND2X2 AND2X2_1301 ( .A(\bus_in[17] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5021_));
AND2X2 AND2X2_1302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5019_), .B(AES_CORE_DATAPATH__abc_16009_new_n5023_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5024_));
AND2X2 AND2X2_1303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5024_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5025_));
AND2X2 AND2X2_1304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5026_));
AND2X2 AND2X2_1305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5029_));
AND2X2 AND2X2_1306 ( .A(\bus_in[18] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5030_));
AND2X2 AND2X2_1307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5028_), .B(AES_CORE_DATAPATH__abc_16009_new_n5032_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5033_));
AND2X2 AND2X2_1308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5033_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5034_));
AND2X2 AND2X2_1309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5035_));
AND2X2 AND2X2_131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2515_), .B(AES_CORE_DATAPATH__abc_16009_new_n2517_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2518_));
AND2X2 AND2X2_1310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5038_));
AND2X2 AND2X2_1311 ( .A(\bus_in[19] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5039_));
AND2X2 AND2X2_1312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5037_), .B(AES_CORE_DATAPATH__abc_16009_new_n5041_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5042_));
AND2X2 AND2X2_1313 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5042_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5043_));
AND2X2 AND2X2_1314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5044_));
AND2X2 AND2X2_1315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5047_));
AND2X2 AND2X2_1316 ( .A(\bus_in[20] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5048_));
AND2X2 AND2X2_1317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5046_), .B(AES_CORE_DATAPATH__abc_16009_new_n5050_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5051_));
AND2X2 AND2X2_1318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5052_), .B(AES_CORE_DATAPATH__abc_16009_new_n5053_), .Y(AES_CORE_DATAPATH__0key_0__31_0__20_));
AND2X2 AND2X2_1319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5056_));
AND2X2 AND2X2_132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2519_));
AND2X2 AND2X2_1320 ( .A(\bus_in[21] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5057_));
AND2X2 AND2X2_1321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5055_), .B(AES_CORE_DATAPATH__abc_16009_new_n5059_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5060_));
AND2X2 AND2X2_1322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5060_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5061_));
AND2X2 AND2X2_1323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5062_));
AND2X2 AND2X2_1324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5065_));
AND2X2 AND2X2_1325 ( .A(\bus_in[22] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5066_));
AND2X2 AND2X2_1326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5064_), .B(AES_CORE_DATAPATH__abc_16009_new_n5068_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5069_));
AND2X2 AND2X2_1327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5069_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5070_));
AND2X2 AND2X2_1328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5071_));
AND2X2 AND2X2_1329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5074_));
AND2X2 AND2X2_133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2521_));
AND2X2 AND2X2_1330 ( .A(\bus_in[23] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5075_));
AND2X2 AND2X2_1331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5073_), .B(AES_CORE_DATAPATH__abc_16009_new_n5077_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5078_));
AND2X2 AND2X2_1332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5079_), .B(AES_CORE_DATAPATH__abc_16009_new_n5080_), .Y(AES_CORE_DATAPATH__0key_0__31_0__23_));
AND2X2 AND2X2_1333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5083_));
AND2X2 AND2X2_1334 ( .A(\bus_in[24] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5084_));
AND2X2 AND2X2_1335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5082_), .B(AES_CORE_DATAPATH__abc_16009_new_n5086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5087_));
AND2X2 AND2X2_1336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5088_), .B(AES_CORE_DATAPATH__abc_16009_new_n5089_), .Y(AES_CORE_DATAPATH__0key_0__31_0__24_));
AND2X2 AND2X2_1337 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5092_));
AND2X2 AND2X2_1338 ( .A(\bus_in[25] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5093_));
AND2X2 AND2X2_1339 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5091_), .B(AES_CORE_DATAPATH__abc_16009_new_n5095_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5096_));
AND2X2 AND2X2_134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2521_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2522_));
AND2X2 AND2X2_1340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5096_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5097_));
AND2X2 AND2X2_1341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5098_));
AND2X2 AND2X2_1342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5101_));
AND2X2 AND2X2_1343 ( .A(\bus_in[26] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5102_));
AND2X2 AND2X2_1344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5100_), .B(AES_CORE_DATAPATH__abc_16009_new_n5104_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5105_));
AND2X2 AND2X2_1345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5106_), .B(AES_CORE_DATAPATH__abc_16009_new_n5107_), .Y(AES_CORE_DATAPATH__0key_0__31_0__26_));
AND2X2 AND2X2_1346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5110_));
AND2X2 AND2X2_1347 ( .A(\bus_in[27] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5111_));
AND2X2 AND2X2_1348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5109_), .B(AES_CORE_DATAPATH__abc_16009_new_n5113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5114_));
AND2X2 AND2X2_1349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5114_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5115_));
AND2X2 AND2X2_135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2523_));
AND2X2 AND2X2_1350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5116_));
AND2X2 AND2X2_1351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5119_));
AND2X2 AND2X2_1352 ( .A(\bus_in[28] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5120_));
AND2X2 AND2X2_1353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5118_), .B(AES_CORE_DATAPATH__abc_16009_new_n5122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5123_));
AND2X2 AND2X2_1354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5124_), .B(AES_CORE_DATAPATH__abc_16009_new_n5125_), .Y(AES_CORE_DATAPATH__0key_0__31_0__28_));
AND2X2 AND2X2_1355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5128_));
AND2X2 AND2X2_1356 ( .A(\bus_in[29] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5129_));
AND2X2 AND2X2_1357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5127_), .B(AES_CORE_DATAPATH__abc_16009_new_n5131_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5132_));
AND2X2 AND2X2_1358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5132_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5133_));
AND2X2 AND2X2_1359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5134_));
AND2X2 AND2X2_136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2526_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2527_));
AND2X2 AND2X2_1360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5137_));
AND2X2 AND2X2_1361 ( .A(\bus_in[30] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5138_));
AND2X2 AND2X2_1362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5136_), .B(AES_CORE_DATAPATH__abc_16009_new_n5140_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5141_));
AND2X2 AND2X2_1363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5142_), .B(AES_CORE_DATAPATH__abc_16009_new_n5143_), .Y(AES_CORE_DATAPATH__0key_0__31_0__30_));
AND2X2 AND2X2_1364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4862_), .B(AES_CORE_DATAPATH_key_host_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5145_));
AND2X2 AND2X2_1365 ( .A(\bus_in[31] ), .B(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5146_));
AND2X2 AND2X2_1366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5149_), .B(AES_CORE_DATAPATH__abc_16009_new_n5148_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5150_));
AND2X2 AND2X2_1367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5150_), .B(AES_CORE_DATAPATH__abc_16009_new_n4865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5151_));
AND2X2 AND2X2_1368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5152_));
AND2X2 AND2X2_1369 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5154_));
AND2X2 AND2X2_137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2525_), .B(AES_CORE_DATAPATH__abc_16009_new_n2527_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2528_));
AND2X2 AND2X2_1370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4869_), .B(AES_CORE_DATAPATH__abc_16009_new_n5155_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5156_));
AND2X2 AND2X2_1371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5159_), .B(AES_CORE_DATAPATH__abc_16009_new_n5158_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__1_));
AND2X2 AND2X2_1372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5162_), .B(AES_CORE_DATAPATH__abc_16009_new_n5161_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__2_));
AND2X2 AND2X2_1373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5165_), .B(AES_CORE_DATAPATH__abc_16009_new_n5164_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__3_));
AND2X2 AND2X2_1374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5168_), .B(AES_CORE_DATAPATH__abc_16009_new_n5167_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__4_));
AND2X2 AND2X2_1375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5171_), .B(AES_CORE_DATAPATH__abc_16009_new_n5170_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__5_));
AND2X2 AND2X2_1376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5174_), .B(AES_CORE_DATAPATH__abc_16009_new_n5173_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__6_));
AND2X2 AND2X2_1377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5177_), .B(AES_CORE_DATAPATH__abc_16009_new_n5176_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__7_));
AND2X2 AND2X2_1378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5180_), .B(AES_CORE_DATAPATH__abc_16009_new_n5179_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__8_));
AND2X2 AND2X2_1379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5183_), .B(AES_CORE_DATAPATH__abc_16009_new_n5182_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__9_));
AND2X2 AND2X2_138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2529_));
AND2X2 AND2X2_1380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5186_), .B(AES_CORE_DATAPATH__abc_16009_new_n5185_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__10_));
AND2X2 AND2X2_1381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5189_), .B(AES_CORE_DATAPATH__abc_16009_new_n5188_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__11_));
AND2X2 AND2X2_1382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5192_), .B(AES_CORE_DATAPATH__abc_16009_new_n5191_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__12_));
AND2X2 AND2X2_1383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5195_), .B(AES_CORE_DATAPATH__abc_16009_new_n5194_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__13_));
AND2X2 AND2X2_1384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5198_), .B(AES_CORE_DATAPATH__abc_16009_new_n5197_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__14_));
AND2X2 AND2X2_1385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5201_), .B(AES_CORE_DATAPATH__abc_16009_new_n5200_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__15_));
AND2X2 AND2X2_1386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5204_), .B(AES_CORE_DATAPATH__abc_16009_new_n5203_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__16_));
AND2X2 AND2X2_1387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5207_), .B(AES_CORE_DATAPATH__abc_16009_new_n5206_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__17_));
AND2X2 AND2X2_1388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5210_), .B(AES_CORE_DATAPATH__abc_16009_new_n5209_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__18_));
AND2X2 AND2X2_1389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5213_), .B(AES_CORE_DATAPATH__abc_16009_new_n5212_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__19_));
AND2X2 AND2X2_139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2531_));
AND2X2 AND2X2_1390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5216_), .B(AES_CORE_DATAPATH__abc_16009_new_n5215_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__20_));
AND2X2 AND2X2_1391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5219_), .B(AES_CORE_DATAPATH__abc_16009_new_n5218_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__21_));
AND2X2 AND2X2_1392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5222_), .B(AES_CORE_DATAPATH__abc_16009_new_n5221_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__22_));
AND2X2 AND2X2_1393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5225_), .B(AES_CORE_DATAPATH__abc_16009_new_n5224_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__23_));
AND2X2 AND2X2_1394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5228_), .B(AES_CORE_DATAPATH__abc_16009_new_n5227_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__24_));
AND2X2 AND2X2_1395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5231_), .B(AES_CORE_DATAPATH__abc_16009_new_n5230_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__25_));
AND2X2 AND2X2_1396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5234_), .B(AES_CORE_DATAPATH__abc_16009_new_n5233_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__26_));
AND2X2 AND2X2_1397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5237_), .B(AES_CORE_DATAPATH__abc_16009_new_n5236_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__27_));
AND2X2 AND2X2_1398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5240_), .B(AES_CORE_DATAPATH__abc_16009_new_n5239_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__28_));
AND2X2 AND2X2_1399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5243_), .B(AES_CORE_DATAPATH__abc_16009_new_n5242_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__29_));
AND2X2 AND2X2_14 ( .A(AES_CORE_CONTROL_UNIT_rd_count_1_), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n88_));
AND2X2 AND2X2_140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2531_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2532_));
AND2X2 AND2X2_1400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5246_), .B(AES_CORE_DATAPATH__abc_16009_new_n5245_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__30_));
AND2X2 AND2X2_1401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5248_), .B(AES_CORE_DATAPATH__abc_16009_new_n5249_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__31_));
AND2X2 AND2X2_1402 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5251_));
AND2X2 AND2X2_1403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5254_), .B(AES_CORE_DATAPATH__abc_16009_new_n5252_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5255_));
AND2X2 AND2X2_1404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5255_), .B(AES_CORE_DATAPATH__abc_16009_new_n5155_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5256_));
AND2X2 AND2X2_1405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5259_));
AND2X2 AND2X2_1406 ( .A(\bus_in[1] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5260_));
AND2X2 AND2X2_1407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5262_), .B(AES_CORE_DATAPATH__abc_16009_new_n5258_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__1_));
AND2X2 AND2X2_1408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5265_));
AND2X2 AND2X2_1409 ( .A(\bus_in[2] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5266_));
AND2X2 AND2X2_141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2533_));
AND2X2 AND2X2_1410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5268_), .B(AES_CORE_DATAPATH__abc_16009_new_n5264_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__2_));
AND2X2 AND2X2_1411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5271_));
AND2X2 AND2X2_1412 ( .A(\bus_in[3] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5272_));
AND2X2 AND2X2_1413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5274_), .B(AES_CORE_DATAPATH__abc_16009_new_n5270_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__3_));
AND2X2 AND2X2_1414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5277_));
AND2X2 AND2X2_1415 ( .A(\bus_in[4] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5278_));
AND2X2 AND2X2_1416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5280_), .B(AES_CORE_DATAPATH__abc_16009_new_n5276_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__4_));
AND2X2 AND2X2_1417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5283_));
AND2X2 AND2X2_1418 ( .A(\bus_in[5] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5284_));
AND2X2 AND2X2_1419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5286_), .B(AES_CORE_DATAPATH__abc_16009_new_n5282_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__5_));
AND2X2 AND2X2_142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2536_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2537_));
AND2X2 AND2X2_1420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5289_));
AND2X2 AND2X2_1421 ( .A(\bus_in[6] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5290_));
AND2X2 AND2X2_1422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5292_), .B(AES_CORE_DATAPATH__abc_16009_new_n5288_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__6_));
AND2X2 AND2X2_1423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5295_));
AND2X2 AND2X2_1424 ( .A(\bus_in[7] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5296_));
AND2X2 AND2X2_1425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5298_), .B(AES_CORE_DATAPATH__abc_16009_new_n5294_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__7_));
AND2X2 AND2X2_1426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5301_));
AND2X2 AND2X2_1427 ( .A(\bus_in[8] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5302_));
AND2X2 AND2X2_1428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5304_), .B(AES_CORE_DATAPATH__abc_16009_new_n5300_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__8_));
AND2X2 AND2X2_1429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5307_));
AND2X2 AND2X2_143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2535_), .B(AES_CORE_DATAPATH__abc_16009_new_n2537_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2538_));
AND2X2 AND2X2_1430 ( .A(\bus_in[9] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5308_));
AND2X2 AND2X2_1431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5310_), .B(AES_CORE_DATAPATH__abc_16009_new_n5306_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__9_));
AND2X2 AND2X2_1432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5313_));
AND2X2 AND2X2_1433 ( .A(\bus_in[10] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5314_));
AND2X2 AND2X2_1434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5316_), .B(AES_CORE_DATAPATH__abc_16009_new_n5312_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__10_));
AND2X2 AND2X2_1435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5319_));
AND2X2 AND2X2_1436 ( .A(\bus_in[11] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5320_));
AND2X2 AND2X2_1437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5322_), .B(AES_CORE_DATAPATH__abc_16009_new_n5318_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__11_));
AND2X2 AND2X2_1438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5325_));
AND2X2 AND2X2_1439 ( .A(\bus_in[12] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5326_));
AND2X2 AND2X2_144 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2539_));
AND2X2 AND2X2_1440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5328_), .B(AES_CORE_DATAPATH__abc_16009_new_n5324_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__12_));
AND2X2 AND2X2_1441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5331_));
AND2X2 AND2X2_1442 ( .A(\bus_in[13] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5332_));
AND2X2 AND2X2_1443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5334_), .B(AES_CORE_DATAPATH__abc_16009_new_n5330_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__13_));
AND2X2 AND2X2_1444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5337_));
AND2X2 AND2X2_1445 ( .A(\bus_in[14] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5338_));
AND2X2 AND2X2_1446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5340_), .B(AES_CORE_DATAPATH__abc_16009_new_n5336_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__14_));
AND2X2 AND2X2_1447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5343_));
AND2X2 AND2X2_1448 ( .A(\bus_in[15] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5344_));
AND2X2 AND2X2_1449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5346_), .B(AES_CORE_DATAPATH__abc_16009_new_n5342_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__15_));
AND2X2 AND2X2_145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2541_));
AND2X2 AND2X2_1450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5349_));
AND2X2 AND2X2_1451 ( .A(\bus_in[16] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5350_));
AND2X2 AND2X2_1452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5352_), .B(AES_CORE_DATAPATH__abc_16009_new_n5348_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__16_));
AND2X2 AND2X2_1453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5355_));
AND2X2 AND2X2_1454 ( .A(\bus_in[17] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5356_));
AND2X2 AND2X2_1455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5358_), .B(AES_CORE_DATAPATH__abc_16009_new_n5354_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__17_));
AND2X2 AND2X2_1456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5361_));
AND2X2 AND2X2_1457 ( .A(\bus_in[18] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5362_));
AND2X2 AND2X2_1458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5364_), .B(AES_CORE_DATAPATH__abc_16009_new_n5360_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__18_));
AND2X2 AND2X2_1459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5367_));
AND2X2 AND2X2_146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2541_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2542_));
AND2X2 AND2X2_1460 ( .A(\bus_in[19] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5368_));
AND2X2 AND2X2_1461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5370_), .B(AES_CORE_DATAPATH__abc_16009_new_n5366_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__19_));
AND2X2 AND2X2_1462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5373_));
AND2X2 AND2X2_1463 ( .A(\bus_in[20] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5374_));
AND2X2 AND2X2_1464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5376_), .B(AES_CORE_DATAPATH__abc_16009_new_n5372_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__20_));
AND2X2 AND2X2_1465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5379_));
AND2X2 AND2X2_1466 ( .A(\bus_in[21] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5380_));
AND2X2 AND2X2_1467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5382_), .B(AES_CORE_DATAPATH__abc_16009_new_n5378_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__21_));
AND2X2 AND2X2_1468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5385_));
AND2X2 AND2X2_1469 ( .A(\bus_in[22] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5386_));
AND2X2 AND2X2_147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2543_));
AND2X2 AND2X2_1470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5388_), .B(AES_CORE_DATAPATH__abc_16009_new_n5384_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__22_));
AND2X2 AND2X2_1471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5391_));
AND2X2 AND2X2_1472 ( .A(\bus_in[23] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5392_));
AND2X2 AND2X2_1473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5394_), .B(AES_CORE_DATAPATH__abc_16009_new_n5390_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__23_));
AND2X2 AND2X2_1474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5397_));
AND2X2 AND2X2_1475 ( .A(\bus_in[24] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5398_));
AND2X2 AND2X2_1476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5400_), .B(AES_CORE_DATAPATH__abc_16009_new_n5396_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__24_));
AND2X2 AND2X2_1477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5403_));
AND2X2 AND2X2_1478 ( .A(\bus_in[25] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5404_));
AND2X2 AND2X2_1479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5406_), .B(AES_CORE_DATAPATH__abc_16009_new_n5402_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__25_));
AND2X2 AND2X2_148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2546_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2547_));
AND2X2 AND2X2_1480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5409_));
AND2X2 AND2X2_1481 ( .A(\bus_in[26] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5410_));
AND2X2 AND2X2_1482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5412_), .B(AES_CORE_DATAPATH__abc_16009_new_n5408_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__26_));
AND2X2 AND2X2_1483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5415_));
AND2X2 AND2X2_1484 ( .A(\bus_in[27] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5416_));
AND2X2 AND2X2_1485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5418_), .B(AES_CORE_DATAPATH__abc_16009_new_n5414_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__27_));
AND2X2 AND2X2_1486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5421_));
AND2X2 AND2X2_1487 ( .A(\bus_in[28] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5422_));
AND2X2 AND2X2_1488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5424_), .B(AES_CORE_DATAPATH__abc_16009_new_n5420_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__28_));
AND2X2 AND2X2_1489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5427_));
AND2X2 AND2X2_149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2545_), .B(AES_CORE_DATAPATH__abc_16009_new_n2547_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2548_));
AND2X2 AND2X2_1490 ( .A(\bus_in[29] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5428_));
AND2X2 AND2X2_1491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5430_), .B(AES_CORE_DATAPATH__abc_16009_new_n5426_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__29_));
AND2X2 AND2X2_1492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5433_));
AND2X2 AND2X2_1493 ( .A(\bus_in[30] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5434_));
AND2X2 AND2X2_1494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5436_), .B(AES_CORE_DATAPATH__abc_16009_new_n5432_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__30_));
AND2X2 AND2X2_1495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(AES_CORE_DATAPATH_key_host_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5438_));
AND2X2 AND2X2_1496 ( .A(\bus_in[31] ), .B(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5439_));
AND2X2 AND2X2_1497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5441_), .B(AES_CORE_DATAPATH__abc_16009_new_n5442_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__31_));
AND2X2 AND2X2_1498 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5444_));
AND2X2 AND2X2_1499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4570_), .B(AES_CORE_DATAPATH__abc_16009_new_n5155_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5445_));
AND2X2 AND2X2_15 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n88_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .Y(AES_CORE_CONTROL_UNIT_last_round));
AND2X2 AND2X2_150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2549_));
AND2X2 AND2X2_1500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5447_), .B(AES_CORE_DATAPATH__abc_16009_new_n5448_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__1_));
AND2X2 AND2X2_1501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5450_), .B(AES_CORE_DATAPATH__abc_16009_new_n5451_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__2_));
AND2X2 AND2X2_1502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5453_), .B(AES_CORE_DATAPATH__abc_16009_new_n5454_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__3_));
AND2X2 AND2X2_1503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5456_), .B(AES_CORE_DATAPATH__abc_16009_new_n5457_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__4_));
AND2X2 AND2X2_1504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5459_), .B(AES_CORE_DATAPATH__abc_16009_new_n5460_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__5_));
AND2X2 AND2X2_1505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5462_), .B(AES_CORE_DATAPATH__abc_16009_new_n5463_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__6_));
AND2X2 AND2X2_1506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5465_), .B(AES_CORE_DATAPATH__abc_16009_new_n5466_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__7_));
AND2X2 AND2X2_1507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5468_), .B(AES_CORE_DATAPATH__abc_16009_new_n5469_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__8_));
AND2X2 AND2X2_1508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5471_), .B(AES_CORE_DATAPATH__abc_16009_new_n5472_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__9_));
AND2X2 AND2X2_1509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5474_), .B(AES_CORE_DATAPATH__abc_16009_new_n5475_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__10_));
AND2X2 AND2X2_151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2551_));
AND2X2 AND2X2_1510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5477_), .B(AES_CORE_DATAPATH__abc_16009_new_n5478_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__11_));
AND2X2 AND2X2_1511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5480_), .B(AES_CORE_DATAPATH__abc_16009_new_n5481_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__12_));
AND2X2 AND2X2_1512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5483_), .B(AES_CORE_DATAPATH__abc_16009_new_n5484_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__13_));
AND2X2 AND2X2_1513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5486_), .B(AES_CORE_DATAPATH__abc_16009_new_n5487_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__14_));
AND2X2 AND2X2_1514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5489_), .B(AES_CORE_DATAPATH__abc_16009_new_n5490_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__15_));
AND2X2 AND2X2_1515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5492_), .B(AES_CORE_DATAPATH__abc_16009_new_n5493_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__16_));
AND2X2 AND2X2_1516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5495_), .B(AES_CORE_DATAPATH__abc_16009_new_n5496_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__17_));
AND2X2 AND2X2_1517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5498_), .B(AES_CORE_DATAPATH__abc_16009_new_n5499_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__18_));
AND2X2 AND2X2_1518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5501_), .B(AES_CORE_DATAPATH__abc_16009_new_n5502_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__19_));
AND2X2 AND2X2_1519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5504_), .B(AES_CORE_DATAPATH__abc_16009_new_n5505_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__20_));
AND2X2 AND2X2_152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2551_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2552_));
AND2X2 AND2X2_1520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5507_), .B(AES_CORE_DATAPATH__abc_16009_new_n5508_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__21_));
AND2X2 AND2X2_1521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5510_), .B(AES_CORE_DATAPATH__abc_16009_new_n5511_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__22_));
AND2X2 AND2X2_1522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5513_), .B(AES_CORE_DATAPATH__abc_16009_new_n5514_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__23_));
AND2X2 AND2X2_1523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5516_), .B(AES_CORE_DATAPATH__abc_16009_new_n5517_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__24_));
AND2X2 AND2X2_1524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5519_), .B(AES_CORE_DATAPATH__abc_16009_new_n5520_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__25_));
AND2X2 AND2X2_1525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5522_), .B(AES_CORE_DATAPATH__abc_16009_new_n5523_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__26_));
AND2X2 AND2X2_1526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5525_), .B(AES_CORE_DATAPATH__abc_16009_new_n5526_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__27_));
AND2X2 AND2X2_1527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5528_), .B(AES_CORE_DATAPATH__abc_16009_new_n5529_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__28_));
AND2X2 AND2X2_1528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5531_), .B(AES_CORE_DATAPATH__abc_16009_new_n5532_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__29_));
AND2X2 AND2X2_1529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5534_), .B(AES_CORE_DATAPATH__abc_16009_new_n5535_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__30_));
AND2X2 AND2X2_153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2553_));
AND2X2 AND2X2_1530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5538_), .B(AES_CORE_DATAPATH__abc_16009_new_n5537_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__31_));
AND2X2 AND2X2_1531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5540_));
AND2X2 AND2X2_1532 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5541_));
AND2X2 AND2X2_1533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4561_), .B(AES_CORE_DATAPATH__abc_16009_new_n5253_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5544_));
AND2X2 AND2X2_1534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5543_), .B(AES_CORE_DATAPATH__abc_16009_new_n5544_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5545_));
AND2X2 AND2X2_1535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5547_), .B(AES_CORE_DATAPATH__abc_16009_new_n5546_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5548_));
AND2X2 AND2X2_1536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5549_), .B(AES_CORE_DATAPATH__abc_16009_new_n5551_), .Y(AES_CORE_DATAPATH__0key_2__31_0__0_));
AND2X2 AND2X2_1537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5554_), .B(AES_CORE_DATAPATH__abc_16009_new_n5553_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5555_));
AND2X2 AND2X2_1538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5556_), .B(AES_CORE_DATAPATH__abc_16009_new_n5557_), .Y(AES_CORE_DATAPATH__0key_2__31_0__1_));
AND2X2 AND2X2_1539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5560_), .B(AES_CORE_DATAPATH__abc_16009_new_n5559_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5561_));
AND2X2 AND2X2_154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2556_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2557_));
AND2X2 AND2X2_1540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5562_), .B(AES_CORE_DATAPATH__abc_16009_new_n5563_), .Y(AES_CORE_DATAPATH__0key_2__31_0__2_));
AND2X2 AND2X2_1541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5565_), .B(AES_CORE_DATAPATH__abc_16009_new_n5566_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5567_));
AND2X2 AND2X2_1542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5568_), .B(AES_CORE_DATAPATH__abc_16009_new_n5569_), .Y(AES_CORE_DATAPATH__0key_2__31_0__3_));
AND2X2 AND2X2_1543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5571_), .B(AES_CORE_DATAPATH__abc_16009_new_n5572_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5573_));
AND2X2 AND2X2_1544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5574_), .B(AES_CORE_DATAPATH__abc_16009_new_n5575_), .Y(AES_CORE_DATAPATH__0key_2__31_0__4_));
AND2X2 AND2X2_1545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5578_), .B(AES_CORE_DATAPATH__abc_16009_new_n5577_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5579_));
AND2X2 AND2X2_1546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5579_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5580_));
AND2X2 AND2X2_1547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5581_));
AND2X2 AND2X2_1548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5583_), .B(AES_CORE_DATAPATH__abc_16009_new_n5584_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5585_));
AND2X2 AND2X2_1549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5586_), .B(AES_CORE_DATAPATH__abc_16009_new_n5587_), .Y(AES_CORE_DATAPATH__0key_2__31_0__6_));
AND2X2 AND2X2_155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2555_), .B(AES_CORE_DATAPATH__abc_16009_new_n2557_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2558_));
AND2X2 AND2X2_1550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5590_), .B(AES_CORE_DATAPATH__abc_16009_new_n5589_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5591_));
AND2X2 AND2X2_1551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5592_), .B(AES_CORE_DATAPATH__abc_16009_new_n5593_), .Y(AES_CORE_DATAPATH__0key_2__31_0__7_));
AND2X2 AND2X2_1552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5596_), .B(AES_CORE_DATAPATH__abc_16009_new_n5595_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5597_));
AND2X2 AND2X2_1553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5598_), .B(AES_CORE_DATAPATH__abc_16009_new_n5599_), .Y(AES_CORE_DATAPATH__0key_2__31_0__8_));
AND2X2 AND2X2_1554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5602_), .B(AES_CORE_DATAPATH__abc_16009_new_n5601_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5603_));
AND2X2 AND2X2_1555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5603_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5604_));
AND2X2 AND2X2_1556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5605_));
AND2X2 AND2X2_1557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5608_), .B(AES_CORE_DATAPATH__abc_16009_new_n5607_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5609_));
AND2X2 AND2X2_1558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5609_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5610_));
AND2X2 AND2X2_1559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5611_));
AND2X2 AND2X2_156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2559_));
AND2X2 AND2X2_1560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5614_), .B(AES_CORE_DATAPATH__abc_16009_new_n5613_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5615_));
AND2X2 AND2X2_1561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5615_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5616_));
AND2X2 AND2X2_1562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5617_));
AND2X2 AND2X2_1563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5619_), .B(AES_CORE_DATAPATH__abc_16009_new_n5620_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5621_));
AND2X2 AND2X2_1564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5622_), .B(AES_CORE_DATAPATH__abc_16009_new_n5623_), .Y(AES_CORE_DATAPATH__0key_2__31_0__12_));
AND2X2 AND2X2_1565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5625_), .B(AES_CORE_DATAPATH__abc_16009_new_n5626_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5627_));
AND2X2 AND2X2_1566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5628_), .B(AES_CORE_DATAPATH__abc_16009_new_n5629_), .Y(AES_CORE_DATAPATH__0key_2__31_0__13_));
AND2X2 AND2X2_1567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5632_), .B(AES_CORE_DATAPATH__abc_16009_new_n5631_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5633_));
AND2X2 AND2X2_1568 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5633_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5634_));
AND2X2 AND2X2_1569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5635_));
AND2X2 AND2X2_157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2561_));
AND2X2 AND2X2_1570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5638_), .B(AES_CORE_DATAPATH__abc_16009_new_n5637_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5639_));
AND2X2 AND2X2_1571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5639_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5640_));
AND2X2 AND2X2_1572 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5641_));
AND2X2 AND2X2_1573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5643_), .B(AES_CORE_DATAPATH__abc_16009_new_n5644_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5645_));
AND2X2 AND2X2_1574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5646_), .B(AES_CORE_DATAPATH__abc_16009_new_n5647_), .Y(AES_CORE_DATAPATH__0key_2__31_0__16_));
AND2X2 AND2X2_1575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5650_), .B(AES_CORE_DATAPATH__abc_16009_new_n5649_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5651_));
AND2X2 AND2X2_1576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5651_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5652_));
AND2X2 AND2X2_1577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5653_));
AND2X2 AND2X2_1578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5656_), .B(AES_CORE_DATAPATH__abc_16009_new_n5655_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5657_));
AND2X2 AND2X2_1579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5657_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5658_));
AND2X2 AND2X2_158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2561_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2562_));
AND2X2 AND2X2_1580 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5659_));
AND2X2 AND2X2_1581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5661_), .B(AES_CORE_DATAPATH__abc_16009_new_n5662_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5663_));
AND2X2 AND2X2_1582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5664_), .B(AES_CORE_DATAPATH__abc_16009_new_n5665_), .Y(AES_CORE_DATAPATH__0key_2__31_0__19_));
AND2X2 AND2X2_1583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5668_), .B(AES_CORE_DATAPATH__abc_16009_new_n5667_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5669_));
AND2X2 AND2X2_1584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5669_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5670_));
AND2X2 AND2X2_1585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5671_));
AND2X2 AND2X2_1586 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5674_), .B(AES_CORE_DATAPATH__abc_16009_new_n5673_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5675_));
AND2X2 AND2X2_1587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5676_), .B(AES_CORE_DATAPATH__abc_16009_new_n5677_), .Y(AES_CORE_DATAPATH__0key_2__31_0__21_));
AND2X2 AND2X2_1588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5680_), .B(AES_CORE_DATAPATH__abc_16009_new_n5679_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5681_));
AND2X2 AND2X2_1589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5682_), .B(AES_CORE_DATAPATH__abc_16009_new_n5683_), .Y(AES_CORE_DATAPATH__0key_2__31_0__22_));
AND2X2 AND2X2_159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2563_));
AND2X2 AND2X2_1590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5686_), .B(AES_CORE_DATAPATH__abc_16009_new_n5685_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5687_));
AND2X2 AND2X2_1591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5688_), .B(AES_CORE_DATAPATH__abc_16009_new_n5689_), .Y(AES_CORE_DATAPATH__0key_2__31_0__23_));
AND2X2 AND2X2_1592 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5692_), .B(AES_CORE_DATAPATH__abc_16009_new_n5691_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5693_));
AND2X2 AND2X2_1593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5694_), .B(AES_CORE_DATAPATH__abc_16009_new_n5695_), .Y(AES_CORE_DATAPATH__0key_2__31_0__24_));
AND2X2 AND2X2_1594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5698_), .B(AES_CORE_DATAPATH__abc_16009_new_n5697_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5699_));
AND2X2 AND2X2_1595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5699_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5700_));
AND2X2 AND2X2_1596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5701_));
AND2X2 AND2X2_1597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5704_), .B(AES_CORE_DATAPATH__abc_16009_new_n5703_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5705_));
AND2X2 AND2X2_1598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5705_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5706_));
AND2X2 AND2X2_1599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5707_));
AND2X2 AND2X2_16 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_));
AND2X2 AND2X2_160 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2566_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2567_));
AND2X2 AND2X2_1600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5710_), .B(AES_CORE_DATAPATH__abc_16009_new_n5709_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5711_));
AND2X2 AND2X2_1601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5712_), .B(AES_CORE_DATAPATH__abc_16009_new_n5713_), .Y(AES_CORE_DATAPATH__0key_2__31_0__27_));
AND2X2 AND2X2_1602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5715_), .B(AES_CORE_DATAPATH__abc_16009_new_n5716_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5717_));
AND2X2 AND2X2_1603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5718_), .B(AES_CORE_DATAPATH__abc_16009_new_n5719_), .Y(AES_CORE_DATAPATH__0key_2__31_0__28_));
AND2X2 AND2X2_1604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5722_), .B(AES_CORE_DATAPATH__abc_16009_new_n5721_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5723_));
AND2X2 AND2X2_1605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5724_), .B(AES_CORE_DATAPATH__abc_16009_new_n5725_), .Y(AES_CORE_DATAPATH__0key_2__31_0__29_));
AND2X2 AND2X2_1606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5728_), .B(AES_CORE_DATAPATH__abc_16009_new_n5727_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5729_));
AND2X2 AND2X2_1607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5729_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5730_));
AND2X2 AND2X2_1608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5731_));
AND2X2 AND2X2_1609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5734_), .B(AES_CORE_DATAPATH__abc_16009_new_n5733_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5735_));
AND2X2 AND2X2_161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2565_), .B(AES_CORE_DATAPATH__abc_16009_new_n2567_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2568_));
AND2X2 AND2X2_1610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5735_), .B(AES_CORE_DATAPATH__abc_16009_new_n5550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5736_));
AND2X2 AND2X2_1611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5737_));
AND2X2 AND2X2_1612 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5740_));
AND2X2 AND2X2_1613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5741_));
AND2X2 AND2X2_1614 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_sel_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5742_));
AND2X2 AND2X2_1615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5745_));
AND2X2 AND2X2_1616 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_sel_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5746_));
AND2X2 AND2X2_1617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5744_), .B(AES_CORE_DATAPATH__abc_16009_new_n5748_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5749_));
AND2X2 AND2X2_1618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5750_));
AND2X2 AND2X2_1619 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5751_));
AND2X2 AND2X2_162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2569_));
AND2X2 AND2X2_1620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n5752_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5753_));
AND2X2 AND2X2_1621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5744_), .B(AES_CORE_DATAPATH__abc_16009_new_n5747_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5754_));
AND2X2 AND2X2_1622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3464_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5755_));
AND2X2 AND2X2_1623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5748_), .B(AES_CORE_DATAPATH__abc_16009_new_n5743_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5756_));
AND2X2 AND2X2_1624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2802_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n5758_));
AND2X2 AND2X2_1625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3464_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5760_));
AND2X2 AND2X2_1626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5761_));
AND2X2 AND2X2_1627 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2802_), .B(first_block), .Y(AES_CORE_DATAPATH__abc_16009_new_n5763_));
AND2X2 AND2X2_1628 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5765_));
AND2X2 AND2X2_1629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5765_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5766_));
AND2X2 AND2X2_163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2571_));
AND2X2 AND2X2_1630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5767_));
AND2X2 AND2X2_1631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5770_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5771_));
AND2X2 AND2X2_1632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5769_), .B(AES_CORE_DATAPATH__abc_16009_new_n5771_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5772_));
AND2X2 AND2X2_1633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5773_));
AND2X2 AND2X2_1634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5774_), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5775_));
AND2X2 AND2X2_1635 ( .A(\iv_out[0] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5776_));
AND2X2 AND2X2_1636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3452_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5780_));
AND2X2 AND2X2_1637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5780_), .B(AES_CORE_DATAPATH__abc_16009_new_n5779_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5781_));
AND2X2 AND2X2_1638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5784_), .B(AES_CORE_DATAPATH__abc_16009_new_n5785_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5786_));
AND2X2 AND2X2_1639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5778_), .B(AES_CORE_DATAPATH__abc_16009_new_n5788_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5789_));
AND2X2 AND2X2_164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2571_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2572_));
AND2X2 AND2X2_1640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5792_), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_16009_new_n5793_));
AND2X2 AND2X2_1641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5791_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5794_));
AND2X2 AND2X2_1642 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5790_), .B(AES_CORE_DATAPATH__abc_16009_new_n5794_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5795_));
AND2X2 AND2X2_1643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5796_));
AND2X2 AND2X2_1644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5799_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n5800_));
AND2X2 AND2X2_1645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5797_), .B(AES_CORE_DATAPATH__abc_16009_new_n5800_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5801_));
AND2X2 AND2X2_1646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2802_), .B(AES_CORE_DATAPATH__abc_16009_new_n5792_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5802_));
AND2X2 AND2X2_1647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5803_));
AND2X2 AND2X2_1648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5805_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5806_));
AND2X2 AND2X2_1649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5808_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5809_));
AND2X2 AND2X2_165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2573_));
AND2X2 AND2X2_1650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5811_));
AND2X2 AND2X2_1651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5812_));
AND2X2 AND2X2_1652 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5813_));
AND2X2 AND2X2_1653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n5814_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5815_));
AND2X2 AND2X2_1654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3487_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5817_));
AND2X2 AND2X2_1655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5817_), .B(AES_CORE_DATAPATH__abc_16009_new_n5816_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5818_));
AND2X2 AND2X2_1656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5820_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5821_));
AND2X2 AND2X2_1657 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5825_));
AND2X2 AND2X2_1658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5825_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5826_));
AND2X2 AND2X2_1659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5827_));
AND2X2 AND2X2_166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2576_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2577_));
AND2X2 AND2X2_1660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5830_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5831_));
AND2X2 AND2X2_1661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5829_), .B(AES_CORE_DATAPATH__abc_16009_new_n5831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5832_));
AND2X2 AND2X2_1662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5833_));
AND2X2 AND2X2_1663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5835_), .B(AES_CORE_DATAPATH__abc_16009_new_n5836_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5837_));
AND2X2 AND2X2_1664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5840_), .B(AES_CORE_DATAPATH__abc_16009_new_n5822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5841_));
AND2X2 AND2X2_1665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5839_), .B(AES_CORE_DATAPATH__abc_16009_new_n5842_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5843_));
AND2X2 AND2X2_1666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5845_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5846_));
AND2X2 AND2X2_1667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5844_), .B(AES_CORE_DATAPATH__abc_16009_new_n5846_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5847_));
AND2X2 AND2X2_1668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5849_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n5850_));
AND2X2 AND2X2_1669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5848_), .B(AES_CORE_DATAPATH__abc_16009_new_n5850_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5851_));
AND2X2 AND2X2_167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2575_), .B(AES_CORE_DATAPATH__abc_16009_new_n2577_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2578_));
AND2X2 AND2X2_1670 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5852_));
AND2X2 AND2X2_1671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5854_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5855_));
AND2X2 AND2X2_1672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3496_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5856_));
AND2X2 AND2X2_1673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5858_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5859_));
AND2X2 AND2X2_1674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5861_));
AND2X2 AND2X2_1675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5862_));
AND2X2 AND2X2_1676 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5863_));
AND2X2 AND2X2_1677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n5864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5865_));
AND2X2 AND2X2_1678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3528_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5866_));
AND2X2 AND2X2_1679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5867_));
AND2X2 AND2X2_168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2579_));
AND2X2 AND2X2_1680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5869_));
AND2X2 AND2X2_1681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5869_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5870_));
AND2X2 AND2X2_1682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5871_));
AND2X2 AND2X2_1683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5874_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5875_));
AND2X2 AND2X2_1684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5873_), .B(AES_CORE_DATAPATH__abc_16009_new_n5875_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5876_));
AND2X2 AND2X2_1685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5877_));
AND2X2 AND2X2_1686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5879_), .B(AES_CORE_DATAPATH__abc_16009_new_n5880_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5881_));
AND2X2 AND2X2_1687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3519_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5884_));
AND2X2 AND2X2_1688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5884_), .B(AES_CORE_DATAPATH__abc_16009_new_n5883_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5885_));
AND2X2 AND2X2_1689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5888_), .B(AES_CORE_DATAPATH__abc_16009_new_n5889_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5890_));
AND2X2 AND2X2_169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2581_));
AND2X2 AND2X2_1690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5882_), .B(AES_CORE_DATAPATH__abc_16009_new_n5892_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5893_));
AND2X2 AND2X2_1691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5895_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5896_));
AND2X2 AND2X2_1692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5894_), .B(AES_CORE_DATAPATH__abc_16009_new_n5896_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5897_));
AND2X2 AND2X2_1693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5899_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n5900_));
AND2X2 AND2X2_1694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5898_), .B(AES_CORE_DATAPATH__abc_16009_new_n5900_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5901_));
AND2X2 AND2X2_1695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5902_));
AND2X2 AND2X2_1696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5904_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5905_));
AND2X2 AND2X2_1697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3528_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5906_));
AND2X2 AND2X2_1698 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5908_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5909_));
AND2X2 AND2X2_1699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5911_));
AND2X2 AND2X2_17 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n91_));
AND2X2 AND2X2_170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2581_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2582_));
AND2X2 AND2X2_1700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5912_));
AND2X2 AND2X2_1701 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5913_));
AND2X2 AND2X2_1702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n5914_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5915_));
AND2X2 AND2X2_1703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3551_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5917_));
AND2X2 AND2X2_1704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5917_), .B(AES_CORE_DATAPATH__abc_16009_new_n5916_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5918_));
AND2X2 AND2X2_1705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5920_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5921_));
AND2X2 AND2X2_1706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5925_));
AND2X2 AND2X2_1707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5925_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5926_));
AND2X2 AND2X2_1708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5927_));
AND2X2 AND2X2_1709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5930_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5931_));
AND2X2 AND2X2_171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2583_));
AND2X2 AND2X2_1710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5929_), .B(AES_CORE_DATAPATH__abc_16009_new_n5931_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5932_));
AND2X2 AND2X2_1711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5933_));
AND2X2 AND2X2_1712 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5935_), .B(AES_CORE_DATAPATH__abc_16009_new_n5936_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5937_));
AND2X2 AND2X2_1713 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5940_), .B(AES_CORE_DATAPATH__abc_16009_new_n5922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5941_));
AND2X2 AND2X2_1714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5939_), .B(AES_CORE_DATAPATH__abc_16009_new_n5942_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5943_));
AND2X2 AND2X2_1715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5945_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5946_));
AND2X2 AND2X2_1716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5944_), .B(AES_CORE_DATAPATH__abc_16009_new_n5946_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5947_));
AND2X2 AND2X2_1717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5949_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n5950_));
AND2X2 AND2X2_1718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5948_), .B(AES_CORE_DATAPATH__abc_16009_new_n5950_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5951_));
AND2X2 AND2X2_1719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5952_));
AND2X2 AND2X2_172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2586_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2587_));
AND2X2 AND2X2_1720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5954_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5955_));
AND2X2 AND2X2_1721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3560_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5956_));
AND2X2 AND2X2_1722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5958_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5959_));
AND2X2 AND2X2_1723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5961_));
AND2X2 AND2X2_1724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5962_));
AND2X2 AND2X2_1725 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5963_));
AND2X2 AND2X2_1726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n5964_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5965_));
AND2X2 AND2X2_1727 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3592_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5966_));
AND2X2 AND2X2_1728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5967_));
AND2X2 AND2X2_1729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5969_));
AND2X2 AND2X2_173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2585_), .B(AES_CORE_DATAPATH__abc_16009_new_n2587_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2588_));
AND2X2 AND2X2_1730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5969_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5970_));
AND2X2 AND2X2_1731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5971_));
AND2X2 AND2X2_1732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5974_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5975_));
AND2X2 AND2X2_1733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5973_), .B(AES_CORE_DATAPATH__abc_16009_new_n5975_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5976_));
AND2X2 AND2X2_1734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5977_));
AND2X2 AND2X2_1735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5979_), .B(AES_CORE_DATAPATH__abc_16009_new_n5980_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5981_));
AND2X2 AND2X2_1736 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3583_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5984_));
AND2X2 AND2X2_1737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5984_), .B(AES_CORE_DATAPATH__abc_16009_new_n5983_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5985_));
AND2X2 AND2X2_1738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5988_), .B(AES_CORE_DATAPATH__abc_16009_new_n5989_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5990_));
AND2X2 AND2X2_1739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5982_), .B(AES_CORE_DATAPATH__abc_16009_new_n5992_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5993_));
AND2X2 AND2X2_174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2589_));
AND2X2 AND2X2_1740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5995_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5996_));
AND2X2 AND2X2_1741 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5994_), .B(AES_CORE_DATAPATH__abc_16009_new_n5996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5997_));
AND2X2 AND2X2_1742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5999_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6000_));
AND2X2 AND2X2_1743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5998_), .B(AES_CORE_DATAPATH__abc_16009_new_n6000_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6001_));
AND2X2 AND2X2_1744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6002_));
AND2X2 AND2X2_1745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6004_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6005_));
AND2X2 AND2X2_1746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3592_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6006_));
AND2X2 AND2X2_1747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6008_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6009_));
AND2X2 AND2X2_1748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6011_));
AND2X2 AND2X2_1749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6012_));
AND2X2 AND2X2_175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2591_));
AND2X2 AND2X2_1750 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6013_));
AND2X2 AND2X2_1751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6015_));
AND2X2 AND2X2_1752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3624_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6016_));
AND2X2 AND2X2_1753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6017_));
AND2X2 AND2X2_1754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6019_));
AND2X2 AND2X2_1755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6019_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6020_));
AND2X2 AND2X2_1756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6021_));
AND2X2 AND2X2_1757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6024_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6025_));
AND2X2 AND2X2_1758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6023_), .B(AES_CORE_DATAPATH__abc_16009_new_n6025_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6026_));
AND2X2 AND2X2_1759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6027_));
AND2X2 AND2X2_176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2591_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2592_));
AND2X2 AND2X2_1760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6029_), .B(AES_CORE_DATAPATH__abc_16009_new_n6030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6031_));
AND2X2 AND2X2_1761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3615_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6034_));
AND2X2 AND2X2_1762 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6034_), .B(AES_CORE_DATAPATH__abc_16009_new_n6033_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6035_));
AND2X2 AND2X2_1763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6038_), .B(AES_CORE_DATAPATH__abc_16009_new_n6039_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6040_));
AND2X2 AND2X2_1764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6032_), .B(AES_CORE_DATAPATH__abc_16009_new_n6042_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6043_));
AND2X2 AND2X2_1765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6045_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6046_));
AND2X2 AND2X2_1766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6044_), .B(AES_CORE_DATAPATH__abc_16009_new_n6046_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6047_));
AND2X2 AND2X2_1767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6049_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6050_));
AND2X2 AND2X2_1768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6048_), .B(AES_CORE_DATAPATH__abc_16009_new_n6050_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6051_));
AND2X2 AND2X2_1769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6052_));
AND2X2 AND2X2_177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2593_));
AND2X2 AND2X2_1770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6054_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6055_));
AND2X2 AND2X2_1771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3624_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6056_));
AND2X2 AND2X2_1772 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6058_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6059_));
AND2X2 AND2X2_1773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6061_));
AND2X2 AND2X2_1774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6062_));
AND2X2 AND2X2_1775 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6063_));
AND2X2 AND2X2_1776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6064_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6065_));
AND2X2 AND2X2_1777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3656_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6066_));
AND2X2 AND2X2_1778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6067_));
AND2X2 AND2X2_1779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6069_));
AND2X2 AND2X2_178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2596_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2597_));
AND2X2 AND2X2_1780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6069_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6070_));
AND2X2 AND2X2_1781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6071_));
AND2X2 AND2X2_1782 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6074_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6075_));
AND2X2 AND2X2_1783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6073_), .B(AES_CORE_DATAPATH__abc_16009_new_n6075_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6076_));
AND2X2 AND2X2_1784 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6077_));
AND2X2 AND2X2_1785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6079_), .B(AES_CORE_DATAPATH__abc_16009_new_n6080_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6081_));
AND2X2 AND2X2_1786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3647_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6084_));
AND2X2 AND2X2_1787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6084_), .B(AES_CORE_DATAPATH__abc_16009_new_n6083_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6085_));
AND2X2 AND2X2_1788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6088_), .B(AES_CORE_DATAPATH__abc_16009_new_n6089_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6090_));
AND2X2 AND2X2_1789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6082_), .B(AES_CORE_DATAPATH__abc_16009_new_n6092_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6093_));
AND2X2 AND2X2_179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2595_), .B(AES_CORE_DATAPATH__abc_16009_new_n2597_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2598_));
AND2X2 AND2X2_1790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6095_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6096_));
AND2X2 AND2X2_1791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6094_), .B(AES_CORE_DATAPATH__abc_16009_new_n6096_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6097_));
AND2X2 AND2X2_1792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6099_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6100_));
AND2X2 AND2X2_1793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6098_), .B(AES_CORE_DATAPATH__abc_16009_new_n6100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6101_));
AND2X2 AND2X2_1794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6102_));
AND2X2 AND2X2_1795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6104_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6105_));
AND2X2 AND2X2_1796 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3656_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6106_));
AND2X2 AND2X2_1797 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6108_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6109_));
AND2X2 AND2X2_1798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6111_));
AND2X2 AND2X2_1799 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6112_));
AND2X2 AND2X2_18 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n74_), .B(\op_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n93_));
AND2X2 AND2X2_180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2599_));
AND2X2 AND2X2_1800 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6113_));
AND2X2 AND2X2_1801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6114_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6115_));
AND2X2 AND2X2_1802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3679_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6117_));
AND2X2 AND2X2_1803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6117_), .B(AES_CORE_DATAPATH__abc_16009_new_n6116_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6118_));
AND2X2 AND2X2_1804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6120_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6121_));
AND2X2 AND2X2_1805 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6125_));
AND2X2 AND2X2_1806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6125_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6126_));
AND2X2 AND2X2_1807 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6127_));
AND2X2 AND2X2_1808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6130_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6131_));
AND2X2 AND2X2_1809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6129_), .B(AES_CORE_DATAPATH__abc_16009_new_n6131_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6132_));
AND2X2 AND2X2_181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2601_));
AND2X2 AND2X2_1810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6133_));
AND2X2 AND2X2_1811 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6135_), .B(AES_CORE_DATAPATH__abc_16009_new_n6136_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6137_));
AND2X2 AND2X2_1812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6140_), .B(AES_CORE_DATAPATH__abc_16009_new_n6122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6141_));
AND2X2 AND2X2_1813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6139_), .B(AES_CORE_DATAPATH__abc_16009_new_n6142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6143_));
AND2X2 AND2X2_1814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6145_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6146_));
AND2X2 AND2X2_1815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6144_), .B(AES_CORE_DATAPATH__abc_16009_new_n6146_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6147_));
AND2X2 AND2X2_1816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6149_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6150_));
AND2X2 AND2X2_1817 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6148_), .B(AES_CORE_DATAPATH__abc_16009_new_n6150_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6151_));
AND2X2 AND2X2_1818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6152_));
AND2X2 AND2X2_1819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6154_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6155_));
AND2X2 AND2X2_182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2601_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2602_));
AND2X2 AND2X2_1820 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3688_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6156_));
AND2X2 AND2X2_1821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6158_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6159_));
AND2X2 AND2X2_1822 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6161_));
AND2X2 AND2X2_1823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6162_));
AND2X2 AND2X2_1824 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6163_));
AND2X2 AND2X2_1825 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6164_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6165_));
AND2X2 AND2X2_1826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3720_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6166_));
AND2X2 AND2X2_1827 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6167_));
AND2X2 AND2X2_1828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6169_));
AND2X2 AND2X2_1829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6169_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6170_));
AND2X2 AND2X2_183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2603_));
AND2X2 AND2X2_1830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6171_));
AND2X2 AND2X2_1831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6174_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6175_));
AND2X2 AND2X2_1832 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6173_), .B(AES_CORE_DATAPATH__abc_16009_new_n6175_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6176_));
AND2X2 AND2X2_1833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6177_));
AND2X2 AND2X2_1834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6179_), .B(AES_CORE_DATAPATH__abc_16009_new_n6180_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6181_));
AND2X2 AND2X2_1835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3711_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6184_));
AND2X2 AND2X2_1836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6184_), .B(AES_CORE_DATAPATH__abc_16009_new_n6183_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6185_));
AND2X2 AND2X2_1837 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6188_), .B(AES_CORE_DATAPATH__abc_16009_new_n6189_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6190_));
AND2X2 AND2X2_1838 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6182_), .B(AES_CORE_DATAPATH__abc_16009_new_n6192_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6193_));
AND2X2 AND2X2_1839 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6195_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6196_));
AND2X2 AND2X2_184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2606_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2607_));
AND2X2 AND2X2_1840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6194_), .B(AES_CORE_DATAPATH__abc_16009_new_n6196_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6197_));
AND2X2 AND2X2_1841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6199_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6200_));
AND2X2 AND2X2_1842 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6198_), .B(AES_CORE_DATAPATH__abc_16009_new_n6200_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6201_));
AND2X2 AND2X2_1843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6202_));
AND2X2 AND2X2_1844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6204_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6205_));
AND2X2 AND2X2_1845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3720_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6206_));
AND2X2 AND2X2_1846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6208_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6209_));
AND2X2 AND2X2_1847 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6211_));
AND2X2 AND2X2_1848 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6212_));
AND2X2 AND2X2_1849 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6213_));
AND2X2 AND2X2_185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2605_), .B(AES_CORE_DATAPATH__abc_16009_new_n2607_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2608_));
AND2X2 AND2X2_1850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6214_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6215_));
AND2X2 AND2X2_1851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3743_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6217_));
AND2X2 AND2X2_1852 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6217_), .B(AES_CORE_DATAPATH__abc_16009_new_n6216_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6218_));
AND2X2 AND2X2_1853 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6220_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6221_));
AND2X2 AND2X2_1854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6225_));
AND2X2 AND2X2_1855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6225_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6226_));
AND2X2 AND2X2_1856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6227_));
AND2X2 AND2X2_1857 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6230_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6231_));
AND2X2 AND2X2_1858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6229_), .B(AES_CORE_DATAPATH__abc_16009_new_n6231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6232_));
AND2X2 AND2X2_1859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6233_));
AND2X2 AND2X2_186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2609_));
AND2X2 AND2X2_1860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6235_), .B(AES_CORE_DATAPATH__abc_16009_new_n6236_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6237_));
AND2X2 AND2X2_1861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6240_), .B(AES_CORE_DATAPATH__abc_16009_new_n6222_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6241_));
AND2X2 AND2X2_1862 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6239_), .B(AES_CORE_DATAPATH__abc_16009_new_n6242_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6243_));
AND2X2 AND2X2_1863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6245_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6246_));
AND2X2 AND2X2_1864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6244_), .B(AES_CORE_DATAPATH__abc_16009_new_n6246_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6247_));
AND2X2 AND2X2_1865 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6249_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6250_));
AND2X2 AND2X2_1866 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6248_), .B(AES_CORE_DATAPATH__abc_16009_new_n6250_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6251_));
AND2X2 AND2X2_1867 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6252_));
AND2X2 AND2X2_1868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6254_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6255_));
AND2X2 AND2X2_1869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3752_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6256_));
AND2X2 AND2X2_187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2611_));
AND2X2 AND2X2_1870 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6258_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6259_));
AND2X2 AND2X2_1871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6261_));
AND2X2 AND2X2_1872 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6262_));
AND2X2 AND2X2_1873 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6263_));
AND2X2 AND2X2_1874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6264_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6265_));
AND2X2 AND2X2_1875 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3784_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6266_));
AND2X2 AND2X2_1876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6267_));
AND2X2 AND2X2_1877 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6269_));
AND2X2 AND2X2_1878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6269_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6270_));
AND2X2 AND2X2_1879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6271_));
AND2X2 AND2X2_188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2611_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2612_));
AND2X2 AND2X2_1880 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6274_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6275_));
AND2X2 AND2X2_1881 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6273_), .B(AES_CORE_DATAPATH__abc_16009_new_n6275_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6276_));
AND2X2 AND2X2_1882 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6277_));
AND2X2 AND2X2_1883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6279_), .B(AES_CORE_DATAPATH__abc_16009_new_n6280_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6281_));
AND2X2 AND2X2_1884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3775_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6284_));
AND2X2 AND2X2_1885 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6284_), .B(AES_CORE_DATAPATH__abc_16009_new_n6283_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6285_));
AND2X2 AND2X2_1886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6288_), .B(AES_CORE_DATAPATH__abc_16009_new_n6289_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6290_));
AND2X2 AND2X2_1887 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6282_), .B(AES_CORE_DATAPATH__abc_16009_new_n6292_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6293_));
AND2X2 AND2X2_1888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6295_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6296_));
AND2X2 AND2X2_1889 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6294_), .B(AES_CORE_DATAPATH__abc_16009_new_n6296_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6297_));
AND2X2 AND2X2_189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2613_));
AND2X2 AND2X2_1890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6299_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6300_));
AND2X2 AND2X2_1891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6298_), .B(AES_CORE_DATAPATH__abc_16009_new_n6300_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6301_));
AND2X2 AND2X2_1892 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6302_));
AND2X2 AND2X2_1893 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6304_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6305_));
AND2X2 AND2X2_1894 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3784_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6306_));
AND2X2 AND2X2_1895 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6308_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6309_));
AND2X2 AND2X2_1896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6311_));
AND2X2 AND2X2_1897 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6312_));
AND2X2 AND2X2_1898 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6313_));
AND2X2 AND2X2_1899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6314_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6315_));
AND2X2 AND2X2_19 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n93_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n92_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n94_));
AND2X2 AND2X2_190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2616_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2617_));
AND2X2 AND2X2_1900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3807_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6317_));
AND2X2 AND2X2_1901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6317_), .B(AES_CORE_DATAPATH__abc_16009_new_n6316_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6318_));
AND2X2 AND2X2_1902 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6320_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6321_));
AND2X2 AND2X2_1903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6325_));
AND2X2 AND2X2_1904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6325_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6326_));
AND2X2 AND2X2_1905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6327_));
AND2X2 AND2X2_1906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6330_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6331_));
AND2X2 AND2X2_1907 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6329_), .B(AES_CORE_DATAPATH__abc_16009_new_n6331_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6332_));
AND2X2 AND2X2_1908 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6333_));
AND2X2 AND2X2_1909 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6335_), .B(AES_CORE_DATAPATH__abc_16009_new_n6336_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6337_));
AND2X2 AND2X2_191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2615_), .B(AES_CORE_DATAPATH__abc_16009_new_n2617_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2618_));
AND2X2 AND2X2_1910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6340_), .B(AES_CORE_DATAPATH__abc_16009_new_n6322_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6341_));
AND2X2 AND2X2_1911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6339_), .B(AES_CORE_DATAPATH__abc_16009_new_n6342_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6343_));
AND2X2 AND2X2_1912 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6345_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6346_));
AND2X2 AND2X2_1913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6344_), .B(AES_CORE_DATAPATH__abc_16009_new_n6346_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6347_));
AND2X2 AND2X2_1914 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6349_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6350_));
AND2X2 AND2X2_1915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6348_), .B(AES_CORE_DATAPATH__abc_16009_new_n6350_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6351_));
AND2X2 AND2X2_1916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6352_));
AND2X2 AND2X2_1917 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6354_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6355_));
AND2X2 AND2X2_1918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3816_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6356_));
AND2X2 AND2X2_1919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6358_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6359_));
AND2X2 AND2X2_192 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2619_));
AND2X2 AND2X2_1920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6361_));
AND2X2 AND2X2_1921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6362_));
AND2X2 AND2X2_1922 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6363_));
AND2X2 AND2X2_1923 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6364_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6365_));
AND2X2 AND2X2_1924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3848_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6366_));
AND2X2 AND2X2_1925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6367_));
AND2X2 AND2X2_1926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6369_));
AND2X2 AND2X2_1927 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6369_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6370_));
AND2X2 AND2X2_1928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6371_));
AND2X2 AND2X2_1929 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6374_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6375_));
AND2X2 AND2X2_193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2621_));
AND2X2 AND2X2_1930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6373_), .B(AES_CORE_DATAPATH__abc_16009_new_n6375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6376_));
AND2X2 AND2X2_1931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6377_));
AND2X2 AND2X2_1932 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6379_), .B(AES_CORE_DATAPATH__abc_16009_new_n6380_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6381_));
AND2X2 AND2X2_1933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3839_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6384_));
AND2X2 AND2X2_1934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6384_), .B(AES_CORE_DATAPATH__abc_16009_new_n6383_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6385_));
AND2X2 AND2X2_1935 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6388_), .B(AES_CORE_DATAPATH__abc_16009_new_n6389_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6390_));
AND2X2 AND2X2_1936 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6382_), .B(AES_CORE_DATAPATH__abc_16009_new_n6392_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6393_));
AND2X2 AND2X2_1937 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6395_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6396_));
AND2X2 AND2X2_1938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6394_), .B(AES_CORE_DATAPATH__abc_16009_new_n6396_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6397_));
AND2X2 AND2X2_1939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6399_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6400_));
AND2X2 AND2X2_194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2621_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2622_));
AND2X2 AND2X2_1940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6398_), .B(AES_CORE_DATAPATH__abc_16009_new_n6400_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6401_));
AND2X2 AND2X2_1941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6402_));
AND2X2 AND2X2_1942 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6404_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6405_));
AND2X2 AND2X2_1943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3848_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6406_));
AND2X2 AND2X2_1944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6408_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6409_));
AND2X2 AND2X2_1945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6411_));
AND2X2 AND2X2_1946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6412_));
AND2X2 AND2X2_1947 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6413_));
AND2X2 AND2X2_1948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6414_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6415_));
AND2X2 AND2X2_1949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3871_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6417_));
AND2X2 AND2X2_195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2623_));
AND2X2 AND2X2_1950 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6417_), .B(AES_CORE_DATAPATH__abc_16009_new_n6416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6418_));
AND2X2 AND2X2_1951 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6420_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6421_));
AND2X2 AND2X2_1952 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6425_));
AND2X2 AND2X2_1953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6425_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6426_));
AND2X2 AND2X2_1954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6427_));
AND2X2 AND2X2_1955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6430_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6431_));
AND2X2 AND2X2_1956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6429_), .B(AES_CORE_DATAPATH__abc_16009_new_n6431_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6432_));
AND2X2 AND2X2_1957 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6433_));
AND2X2 AND2X2_1958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6435_), .B(AES_CORE_DATAPATH__abc_16009_new_n6436_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6437_));
AND2X2 AND2X2_1959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6440_), .B(AES_CORE_DATAPATH__abc_16009_new_n6422_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6441_));
AND2X2 AND2X2_196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2626_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2627_));
AND2X2 AND2X2_1960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6439_), .B(AES_CORE_DATAPATH__abc_16009_new_n6442_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6443_));
AND2X2 AND2X2_1961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6445_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6446_));
AND2X2 AND2X2_1962 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6444_), .B(AES_CORE_DATAPATH__abc_16009_new_n6446_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6447_));
AND2X2 AND2X2_1963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6449_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6450_));
AND2X2 AND2X2_1964 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6448_), .B(AES_CORE_DATAPATH__abc_16009_new_n6450_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6451_));
AND2X2 AND2X2_1965 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6452_));
AND2X2 AND2X2_1966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6454_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6455_));
AND2X2 AND2X2_1967 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3880_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6456_));
AND2X2 AND2X2_1968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6458_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6459_));
AND2X2 AND2X2_1969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6461_));
AND2X2 AND2X2_197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2625_), .B(AES_CORE_DATAPATH__abc_16009_new_n2627_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2628_));
AND2X2 AND2X2_1970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6462_));
AND2X2 AND2X2_1971 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6463_));
AND2X2 AND2X2_1972 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6464_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6465_));
AND2X2 AND2X2_1973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3912_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6466_));
AND2X2 AND2X2_1974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6467_));
AND2X2 AND2X2_1975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6469_));
AND2X2 AND2X2_1976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6469_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6470_));
AND2X2 AND2X2_1977 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6471_));
AND2X2 AND2X2_1978 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6474_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6475_));
AND2X2 AND2X2_1979 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6473_), .B(AES_CORE_DATAPATH__abc_16009_new_n6475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6476_));
AND2X2 AND2X2_198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2629_));
AND2X2 AND2X2_1980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6477_));
AND2X2 AND2X2_1981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6479_), .B(AES_CORE_DATAPATH__abc_16009_new_n6480_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6481_));
AND2X2 AND2X2_1982 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3903_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6484_));
AND2X2 AND2X2_1983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6484_), .B(AES_CORE_DATAPATH__abc_16009_new_n6483_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6485_));
AND2X2 AND2X2_1984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6488_), .B(AES_CORE_DATAPATH__abc_16009_new_n6489_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6490_));
AND2X2 AND2X2_1985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6482_), .B(AES_CORE_DATAPATH__abc_16009_new_n6492_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6493_));
AND2X2 AND2X2_1986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6495_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6496_));
AND2X2 AND2X2_1987 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6494_), .B(AES_CORE_DATAPATH__abc_16009_new_n6496_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6497_));
AND2X2 AND2X2_1988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6499_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6500_));
AND2X2 AND2X2_1989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6498_), .B(AES_CORE_DATAPATH__abc_16009_new_n6500_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6501_));
AND2X2 AND2X2_199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2631_));
AND2X2 AND2X2_1990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6502_));
AND2X2 AND2X2_1991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6504_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6505_));
AND2X2 AND2X2_1992 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3912_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6506_));
AND2X2 AND2X2_1993 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6508_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6509_));
AND2X2 AND2X2_1994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6511_));
AND2X2 AND2X2_1995 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6512_));
AND2X2 AND2X2_1996 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6513_));
AND2X2 AND2X2_1997 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6514_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6515_));
AND2X2 AND2X2_1998 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3935_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6517_));
AND2X2 AND2X2_1999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6517_), .B(AES_CORE_DATAPATH__abc_16009_new_n6516_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6518_));
AND2X2 AND2X2_2 ( .A(_abc_15574_new_n13_), .B(_abc_15574_new_n11_), .Y(AES_CORE_DATAPATH_col_en_host_0_));
AND2X2 AND2X2_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n94_), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n95_));
AND2X2 AND2X2_200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2631_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2632_));
AND2X2 AND2X2_2000 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6520_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6521_));
AND2X2 AND2X2_2001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6525_));
AND2X2 AND2X2_2002 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6525_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6526_));
AND2X2 AND2X2_2003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6527_));
AND2X2 AND2X2_2004 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6530_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6531_));
AND2X2 AND2X2_2005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6529_), .B(AES_CORE_DATAPATH__abc_16009_new_n6531_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6532_));
AND2X2 AND2X2_2006 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6533_));
AND2X2 AND2X2_2007 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6535_), .B(AES_CORE_DATAPATH__abc_16009_new_n6536_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6537_));
AND2X2 AND2X2_2008 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6540_), .B(AES_CORE_DATAPATH__abc_16009_new_n6522_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6541_));
AND2X2 AND2X2_2009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6539_), .B(AES_CORE_DATAPATH__abc_16009_new_n6542_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6543_));
AND2X2 AND2X2_201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2633_));
AND2X2 AND2X2_2010 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6545_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6546_));
AND2X2 AND2X2_2011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6544_), .B(AES_CORE_DATAPATH__abc_16009_new_n6546_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6547_));
AND2X2 AND2X2_2012 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6549_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6550_));
AND2X2 AND2X2_2013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6548_), .B(AES_CORE_DATAPATH__abc_16009_new_n6550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6551_));
AND2X2 AND2X2_2014 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6552_));
AND2X2 AND2X2_2015 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6554_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6555_));
AND2X2 AND2X2_2016 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3944_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6556_));
AND2X2 AND2X2_2017 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6558_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6559_));
AND2X2 AND2X2_2018 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6561_));
AND2X2 AND2X2_2019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6562_));
AND2X2 AND2X2_202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2636_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2637_));
AND2X2 AND2X2_2020 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6563_));
AND2X2 AND2X2_2021 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6565_));
AND2X2 AND2X2_2022 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3976_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6566_));
AND2X2 AND2X2_2023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6567_));
AND2X2 AND2X2_2024 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6569_));
AND2X2 AND2X2_2025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6569_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6570_));
AND2X2 AND2X2_2026 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6571_));
AND2X2 AND2X2_2027 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6574_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6575_));
AND2X2 AND2X2_2028 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6573_), .B(AES_CORE_DATAPATH__abc_16009_new_n6575_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6576_));
AND2X2 AND2X2_2029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6577_));
AND2X2 AND2X2_203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2635_), .B(AES_CORE_DATAPATH__abc_16009_new_n2637_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2638_));
AND2X2 AND2X2_2030 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6579_), .B(AES_CORE_DATAPATH__abc_16009_new_n6580_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6581_));
AND2X2 AND2X2_2031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3967_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6584_));
AND2X2 AND2X2_2032 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6584_), .B(AES_CORE_DATAPATH__abc_16009_new_n6583_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6585_));
AND2X2 AND2X2_2033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6588_), .B(AES_CORE_DATAPATH__abc_16009_new_n6589_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6590_));
AND2X2 AND2X2_2034 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6582_), .B(AES_CORE_DATAPATH__abc_16009_new_n6592_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6593_));
AND2X2 AND2X2_2035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6595_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6596_));
AND2X2 AND2X2_2036 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6594_), .B(AES_CORE_DATAPATH__abc_16009_new_n6596_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6597_));
AND2X2 AND2X2_2037 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6599_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6600_));
AND2X2 AND2X2_2038 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6598_), .B(AES_CORE_DATAPATH__abc_16009_new_n6600_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6601_));
AND2X2 AND2X2_2039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6602_));
AND2X2 AND2X2_204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2639_));
AND2X2 AND2X2_2040 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6604_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6605_));
AND2X2 AND2X2_2041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3976_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6606_));
AND2X2 AND2X2_2042 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6608_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6609_));
AND2X2 AND2X2_2043 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6611_));
AND2X2 AND2X2_2044 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6612_));
AND2X2 AND2X2_2045 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6613_));
AND2X2 AND2X2_2046 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6614_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6615_));
AND2X2 AND2X2_2047 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3999_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6617_));
AND2X2 AND2X2_2048 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6617_), .B(AES_CORE_DATAPATH__abc_16009_new_n6616_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6618_));
AND2X2 AND2X2_2049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6620_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6621_));
AND2X2 AND2X2_205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2641_));
AND2X2 AND2X2_2050 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6625_));
AND2X2 AND2X2_2051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6625_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6626_));
AND2X2 AND2X2_2052 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6627_));
AND2X2 AND2X2_2053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6630_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6631_));
AND2X2 AND2X2_2054 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6629_), .B(AES_CORE_DATAPATH__abc_16009_new_n6631_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6632_));
AND2X2 AND2X2_2055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6633_));
AND2X2 AND2X2_2056 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6635_), .B(AES_CORE_DATAPATH__abc_16009_new_n6636_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6637_));
AND2X2 AND2X2_2057 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6640_), .B(AES_CORE_DATAPATH__abc_16009_new_n6622_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6641_));
AND2X2 AND2X2_2058 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6639_), .B(AES_CORE_DATAPATH__abc_16009_new_n6642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6643_));
AND2X2 AND2X2_2059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6645_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6646_));
AND2X2 AND2X2_206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2641_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2642_));
AND2X2 AND2X2_2060 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6644_), .B(AES_CORE_DATAPATH__abc_16009_new_n6646_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6647_));
AND2X2 AND2X2_2061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6649_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6650_));
AND2X2 AND2X2_2062 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6648_), .B(AES_CORE_DATAPATH__abc_16009_new_n6650_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6651_));
AND2X2 AND2X2_2063 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6652_));
AND2X2 AND2X2_2064 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6654_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6655_));
AND2X2 AND2X2_2065 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4008_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6656_));
AND2X2 AND2X2_2066 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6658_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6659_));
AND2X2 AND2X2_2067 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6661_));
AND2X2 AND2X2_2068 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6662_));
AND2X2 AND2X2_2069 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6663_));
AND2X2 AND2X2_207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2643_));
AND2X2 AND2X2_2070 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6664_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6665_));
AND2X2 AND2X2_2071 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4031_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6667_));
AND2X2 AND2X2_2072 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6667_), .B(AES_CORE_DATAPATH__abc_16009_new_n6666_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6668_));
AND2X2 AND2X2_2073 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6670_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6671_));
AND2X2 AND2X2_2074 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6675_));
AND2X2 AND2X2_2075 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6675_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6676_));
AND2X2 AND2X2_2076 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6677_));
AND2X2 AND2X2_2077 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6680_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6681_));
AND2X2 AND2X2_2078 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6679_), .B(AES_CORE_DATAPATH__abc_16009_new_n6681_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6682_));
AND2X2 AND2X2_2079 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6683_));
AND2X2 AND2X2_208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2646_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2647_));
AND2X2 AND2X2_2080 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6685_), .B(AES_CORE_DATAPATH__abc_16009_new_n6686_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6687_));
AND2X2 AND2X2_2081 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6690_), .B(AES_CORE_DATAPATH__abc_16009_new_n6672_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6691_));
AND2X2 AND2X2_2082 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6689_), .B(AES_CORE_DATAPATH__abc_16009_new_n6692_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6693_));
AND2X2 AND2X2_2083 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6695_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6696_));
AND2X2 AND2X2_2084 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6694_), .B(AES_CORE_DATAPATH__abc_16009_new_n6696_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6697_));
AND2X2 AND2X2_2085 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6699_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6700_));
AND2X2 AND2X2_2086 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6698_), .B(AES_CORE_DATAPATH__abc_16009_new_n6700_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6701_));
AND2X2 AND2X2_2087 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6702_));
AND2X2 AND2X2_2088 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6704_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6705_));
AND2X2 AND2X2_2089 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4040_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6706_));
AND2X2 AND2X2_209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2645_), .B(AES_CORE_DATAPATH__abc_16009_new_n2647_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2648_));
AND2X2 AND2X2_2090 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6708_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6709_));
AND2X2 AND2X2_2091 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6711_));
AND2X2 AND2X2_2092 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6712_));
AND2X2 AND2X2_2093 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6713_));
AND2X2 AND2X2_2094 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6714_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6715_));
AND2X2 AND2X2_2095 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4063_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6717_));
AND2X2 AND2X2_2096 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6717_), .B(AES_CORE_DATAPATH__abc_16009_new_n6716_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6718_));
AND2X2 AND2X2_2097 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6720_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6721_));
AND2X2 AND2X2_2098 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6725_));
AND2X2 AND2X2_2099 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6725_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6726_));
AND2X2 AND2X2_21 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n97_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_5_));
AND2X2 AND2X2_210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2649_));
AND2X2 AND2X2_2100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6727_));
AND2X2 AND2X2_2101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6730_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6731_));
AND2X2 AND2X2_2102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6729_), .B(AES_CORE_DATAPATH__abc_16009_new_n6731_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6732_));
AND2X2 AND2X2_2103 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6733_));
AND2X2 AND2X2_2104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6735_), .B(AES_CORE_DATAPATH__abc_16009_new_n6736_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6737_));
AND2X2 AND2X2_2105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6740_), .B(AES_CORE_DATAPATH__abc_16009_new_n6722_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6741_));
AND2X2 AND2X2_2106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6739_), .B(AES_CORE_DATAPATH__abc_16009_new_n6742_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6743_));
AND2X2 AND2X2_2107 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6745_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6746_));
AND2X2 AND2X2_2108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6744_), .B(AES_CORE_DATAPATH__abc_16009_new_n6746_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6747_));
AND2X2 AND2X2_2109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6749_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6750_));
AND2X2 AND2X2_211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2651_));
AND2X2 AND2X2_2110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6748_), .B(AES_CORE_DATAPATH__abc_16009_new_n6750_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6751_));
AND2X2 AND2X2_2111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6752_));
AND2X2 AND2X2_2112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6754_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6755_));
AND2X2 AND2X2_2113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4072_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6756_));
AND2X2 AND2X2_2114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6758_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6759_));
AND2X2 AND2X2_2115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6761_));
AND2X2 AND2X2_2116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6762_));
AND2X2 AND2X2_2117 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6763_));
AND2X2 AND2X2_2118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6765_));
AND2X2 AND2X2_2119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4104_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6766_));
AND2X2 AND2X2_212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2651_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2652_));
AND2X2 AND2X2_2120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6767_));
AND2X2 AND2X2_2121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6769_));
AND2X2 AND2X2_2122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6769_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6770_));
AND2X2 AND2X2_2123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6771_));
AND2X2 AND2X2_2124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6774_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6775_));
AND2X2 AND2X2_2125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6773_), .B(AES_CORE_DATAPATH__abc_16009_new_n6775_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6776_));
AND2X2 AND2X2_2126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6777_));
AND2X2 AND2X2_2127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6779_), .B(AES_CORE_DATAPATH__abc_16009_new_n6780_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6781_));
AND2X2 AND2X2_2128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4095_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6784_));
AND2X2 AND2X2_2129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6784_), .B(AES_CORE_DATAPATH__abc_16009_new_n6783_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6785_));
AND2X2 AND2X2_213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2653_));
AND2X2 AND2X2_2130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6788_), .B(AES_CORE_DATAPATH__abc_16009_new_n6789_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6790_));
AND2X2 AND2X2_2131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6782_), .B(AES_CORE_DATAPATH__abc_16009_new_n6792_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6793_));
AND2X2 AND2X2_2132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6795_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6796_));
AND2X2 AND2X2_2133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6794_), .B(AES_CORE_DATAPATH__abc_16009_new_n6796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6797_));
AND2X2 AND2X2_2134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6799_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6800_));
AND2X2 AND2X2_2135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6798_), .B(AES_CORE_DATAPATH__abc_16009_new_n6800_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6801_));
AND2X2 AND2X2_2136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6802_));
AND2X2 AND2X2_2137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6804_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6805_));
AND2X2 AND2X2_2138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4104_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6806_));
AND2X2 AND2X2_2139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6808_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6809_));
AND2X2 AND2X2_214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2656_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2657_));
AND2X2 AND2X2_2140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6811_));
AND2X2 AND2X2_2141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6812_));
AND2X2 AND2X2_2142 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6813_));
AND2X2 AND2X2_2143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6814_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6815_));
AND2X2 AND2X2_2144 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4127_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6817_));
AND2X2 AND2X2_2145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6817_), .B(AES_CORE_DATAPATH__abc_16009_new_n6816_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6818_));
AND2X2 AND2X2_2146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6820_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6821_));
AND2X2 AND2X2_2147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6825_));
AND2X2 AND2X2_2148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6825_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6826_));
AND2X2 AND2X2_2149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6827_));
AND2X2 AND2X2_215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2655_), .B(AES_CORE_DATAPATH__abc_16009_new_n2657_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2658_));
AND2X2 AND2X2_2150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6830_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6831_));
AND2X2 AND2X2_2151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6829_), .B(AES_CORE_DATAPATH__abc_16009_new_n6831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6832_));
AND2X2 AND2X2_2152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6833_));
AND2X2 AND2X2_2153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6835_), .B(AES_CORE_DATAPATH__abc_16009_new_n6836_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6837_));
AND2X2 AND2X2_2154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6840_), .B(AES_CORE_DATAPATH__abc_16009_new_n6822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6841_));
AND2X2 AND2X2_2155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6839_), .B(AES_CORE_DATAPATH__abc_16009_new_n6842_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6843_));
AND2X2 AND2X2_2156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6845_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6846_));
AND2X2 AND2X2_2157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6844_), .B(AES_CORE_DATAPATH__abc_16009_new_n6846_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6847_));
AND2X2 AND2X2_2158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6849_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6850_));
AND2X2 AND2X2_2159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6848_), .B(AES_CORE_DATAPATH__abc_16009_new_n6850_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6851_));
AND2X2 AND2X2_216 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2659_));
AND2X2 AND2X2_2160 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6852_));
AND2X2 AND2X2_2161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6854_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6855_));
AND2X2 AND2X2_2162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4136_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6856_));
AND2X2 AND2X2_2163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6858_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6859_));
AND2X2 AND2X2_2164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6861_));
AND2X2 AND2X2_2165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6862_));
AND2X2 AND2X2_2166 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6863_));
AND2X2 AND2X2_2167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6865_));
AND2X2 AND2X2_2168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4168_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6866_));
AND2X2 AND2X2_2169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6867_));
AND2X2 AND2X2_217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2661_));
AND2X2 AND2X2_2170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6869_));
AND2X2 AND2X2_2171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6869_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6870_));
AND2X2 AND2X2_2172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6871_));
AND2X2 AND2X2_2173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6874_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6875_));
AND2X2 AND2X2_2174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6873_), .B(AES_CORE_DATAPATH__abc_16009_new_n6875_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6876_));
AND2X2 AND2X2_2175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6877_));
AND2X2 AND2X2_2176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6879_), .B(AES_CORE_DATAPATH__abc_16009_new_n6880_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6881_));
AND2X2 AND2X2_2177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4159_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6884_));
AND2X2 AND2X2_2178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6884_), .B(AES_CORE_DATAPATH__abc_16009_new_n6883_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6885_));
AND2X2 AND2X2_2179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6888_), .B(AES_CORE_DATAPATH__abc_16009_new_n6889_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6890_));
AND2X2 AND2X2_218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2661_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2662_));
AND2X2 AND2X2_2180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6882_), .B(AES_CORE_DATAPATH__abc_16009_new_n6892_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6893_));
AND2X2 AND2X2_2181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6895_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6896_));
AND2X2 AND2X2_2182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6894_), .B(AES_CORE_DATAPATH__abc_16009_new_n6896_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6897_));
AND2X2 AND2X2_2183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6899_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6900_));
AND2X2 AND2X2_2184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6898_), .B(AES_CORE_DATAPATH__abc_16009_new_n6900_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6901_));
AND2X2 AND2X2_2185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6902_));
AND2X2 AND2X2_2186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6904_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6905_));
AND2X2 AND2X2_2187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4168_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6906_));
AND2X2 AND2X2_2188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6908_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6909_));
AND2X2 AND2X2_2189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6911_));
AND2X2 AND2X2_219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2663_));
AND2X2 AND2X2_2190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6912_));
AND2X2 AND2X2_2191 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6913_));
AND2X2 AND2X2_2192 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6914_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6915_));
AND2X2 AND2X2_2193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4191_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6917_));
AND2X2 AND2X2_2194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6917_), .B(AES_CORE_DATAPATH__abc_16009_new_n6916_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6918_));
AND2X2 AND2X2_2195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6920_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6921_));
AND2X2 AND2X2_2196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6925_));
AND2X2 AND2X2_2197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6925_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6926_));
AND2X2 AND2X2_2198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6927_));
AND2X2 AND2X2_2199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6930_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6931_));
AND2X2 AND2X2_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n90_), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n100_));
AND2X2 AND2X2_220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2666_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2667_));
AND2X2 AND2X2_2200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6929_), .B(AES_CORE_DATAPATH__abc_16009_new_n6931_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6932_));
AND2X2 AND2X2_2201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6933_));
AND2X2 AND2X2_2202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6935_), .B(AES_CORE_DATAPATH__abc_16009_new_n6936_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6937_));
AND2X2 AND2X2_2203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6940_), .B(AES_CORE_DATAPATH__abc_16009_new_n6922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6941_));
AND2X2 AND2X2_2204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6939_), .B(AES_CORE_DATAPATH__abc_16009_new_n6942_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6943_));
AND2X2 AND2X2_2205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6945_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6946_));
AND2X2 AND2X2_2206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6944_), .B(AES_CORE_DATAPATH__abc_16009_new_n6946_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6947_));
AND2X2 AND2X2_2207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6949_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n6950_));
AND2X2 AND2X2_2208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6948_), .B(AES_CORE_DATAPATH__abc_16009_new_n6950_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6951_));
AND2X2 AND2X2_2209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6952_));
AND2X2 AND2X2_221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2665_), .B(AES_CORE_DATAPATH__abc_16009_new_n2667_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2668_));
AND2X2 AND2X2_2210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6954_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6955_));
AND2X2 AND2X2_2211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4200_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6956_));
AND2X2 AND2X2_2212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6958_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6959_));
AND2X2 AND2X2_2213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6961_));
AND2X2 AND2X2_2214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6962_));
AND2X2 AND2X2_2215 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6963_));
AND2X2 AND2X2_2216 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n6964_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6965_));
AND2X2 AND2X2_2217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4232_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6966_));
AND2X2 AND2X2_2218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6967_));
AND2X2 AND2X2_2219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6969_));
AND2X2 AND2X2_222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2669_));
AND2X2 AND2X2_2220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6969_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6970_));
AND2X2 AND2X2_2221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6971_));
AND2X2 AND2X2_2222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6974_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6975_));
AND2X2 AND2X2_2223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6973_), .B(AES_CORE_DATAPATH__abc_16009_new_n6975_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6976_));
AND2X2 AND2X2_2224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6977_));
AND2X2 AND2X2_2225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6979_), .B(AES_CORE_DATAPATH__abc_16009_new_n6980_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6981_));
AND2X2 AND2X2_2226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4223_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6984_));
AND2X2 AND2X2_2227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6984_), .B(AES_CORE_DATAPATH__abc_16009_new_n6983_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6985_));
AND2X2 AND2X2_2228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6988_), .B(AES_CORE_DATAPATH__abc_16009_new_n6989_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6990_));
AND2X2 AND2X2_2229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6982_), .B(AES_CORE_DATAPATH__abc_16009_new_n6992_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6993_));
AND2X2 AND2X2_223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2671_));
AND2X2 AND2X2_2230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6995_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6996_));
AND2X2 AND2X2_2231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6994_), .B(AES_CORE_DATAPATH__abc_16009_new_n6996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6997_));
AND2X2 AND2X2_2232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6999_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7000_));
AND2X2 AND2X2_2233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6998_), .B(AES_CORE_DATAPATH__abc_16009_new_n7000_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7001_));
AND2X2 AND2X2_2234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7002_));
AND2X2 AND2X2_2235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7004_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7005_));
AND2X2 AND2X2_2236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4232_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7006_));
AND2X2 AND2X2_2237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7008_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7009_));
AND2X2 AND2X2_2238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7011_));
AND2X2 AND2X2_2239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7012_));
AND2X2 AND2X2_224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2671_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2672_));
AND2X2 AND2X2_2240 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7013_));
AND2X2 AND2X2_2241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7015_));
AND2X2 AND2X2_2242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4255_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7017_));
AND2X2 AND2X2_2243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7017_), .B(AES_CORE_DATAPATH__abc_16009_new_n7016_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7018_));
AND2X2 AND2X2_2244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7020_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7021_));
AND2X2 AND2X2_2245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7025_));
AND2X2 AND2X2_2246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7025_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7026_));
AND2X2 AND2X2_2247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7027_));
AND2X2 AND2X2_2248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7030_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7031_));
AND2X2 AND2X2_2249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7029_), .B(AES_CORE_DATAPATH__abc_16009_new_n7031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7032_));
AND2X2 AND2X2_225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2673_));
AND2X2 AND2X2_2250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7033_));
AND2X2 AND2X2_2251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7035_), .B(AES_CORE_DATAPATH__abc_16009_new_n7036_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7037_));
AND2X2 AND2X2_2252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7040_), .B(AES_CORE_DATAPATH__abc_16009_new_n7022_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7041_));
AND2X2 AND2X2_2253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7039_), .B(AES_CORE_DATAPATH__abc_16009_new_n7042_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7043_));
AND2X2 AND2X2_2254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7045_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7046_));
AND2X2 AND2X2_2255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7044_), .B(AES_CORE_DATAPATH__abc_16009_new_n7046_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7047_));
AND2X2 AND2X2_2256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7049_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7050_));
AND2X2 AND2X2_2257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7048_), .B(AES_CORE_DATAPATH__abc_16009_new_n7050_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7051_));
AND2X2 AND2X2_2258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7052_));
AND2X2 AND2X2_2259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7054_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7055_));
AND2X2 AND2X2_226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2676_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2677_));
AND2X2 AND2X2_2260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4264_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7056_));
AND2X2 AND2X2_2261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7058_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7059_));
AND2X2 AND2X2_2262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7061_));
AND2X2 AND2X2_2263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7062_));
AND2X2 AND2X2_2264 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7063_));
AND2X2 AND2X2_2265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7064_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7065_));
AND2X2 AND2X2_2266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4287_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7067_));
AND2X2 AND2X2_2267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7067_), .B(AES_CORE_DATAPATH__abc_16009_new_n7066_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7068_));
AND2X2 AND2X2_2268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7070_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7071_));
AND2X2 AND2X2_2269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7075_));
AND2X2 AND2X2_227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2675_), .B(AES_CORE_DATAPATH__abc_16009_new_n2677_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2678_));
AND2X2 AND2X2_2270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7075_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7076_));
AND2X2 AND2X2_2271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7077_));
AND2X2 AND2X2_2272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7080_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7081_));
AND2X2 AND2X2_2273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7079_), .B(AES_CORE_DATAPATH__abc_16009_new_n7081_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7082_));
AND2X2 AND2X2_2274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7083_));
AND2X2 AND2X2_2275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7085_), .B(AES_CORE_DATAPATH__abc_16009_new_n7086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7087_));
AND2X2 AND2X2_2276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7090_), .B(AES_CORE_DATAPATH__abc_16009_new_n7072_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7091_));
AND2X2 AND2X2_2277 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7089_), .B(AES_CORE_DATAPATH__abc_16009_new_n7092_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7093_));
AND2X2 AND2X2_2278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7095_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7096_));
AND2X2 AND2X2_2279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7094_), .B(AES_CORE_DATAPATH__abc_16009_new_n7096_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7097_));
AND2X2 AND2X2_228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2679_));
AND2X2 AND2X2_2280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7099_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7100_));
AND2X2 AND2X2_2281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7098_), .B(AES_CORE_DATAPATH__abc_16009_new_n7100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7101_));
AND2X2 AND2X2_2282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7102_));
AND2X2 AND2X2_2283 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7104_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7105_));
AND2X2 AND2X2_2284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4296_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7106_));
AND2X2 AND2X2_2285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7108_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7109_));
AND2X2 AND2X2_2286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7111_));
AND2X2 AND2X2_2287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7112_));
AND2X2 AND2X2_2288 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7113_));
AND2X2 AND2X2_2289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7114_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7115_));
AND2X2 AND2X2_229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2681_));
AND2X2 AND2X2_2290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4328_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7116_));
AND2X2 AND2X2_2291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7117_));
AND2X2 AND2X2_2292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7119_));
AND2X2 AND2X2_2293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7119_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7120_));
AND2X2 AND2X2_2294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7121_));
AND2X2 AND2X2_2295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7124_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7125_));
AND2X2 AND2X2_2296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7123_), .B(AES_CORE_DATAPATH__abc_16009_new_n7125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7126_));
AND2X2 AND2X2_2297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7127_));
AND2X2 AND2X2_2298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7129_), .B(AES_CORE_DATAPATH__abc_16009_new_n7130_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7131_));
AND2X2 AND2X2_2299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4319_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7134_));
AND2X2 AND2X2_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n99_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n100_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n101_));
AND2X2 AND2X2_230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2681_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2682_));
AND2X2 AND2X2_2300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7134_), .B(AES_CORE_DATAPATH__abc_16009_new_n7133_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7135_));
AND2X2 AND2X2_2301 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7138_), .B(AES_CORE_DATAPATH__abc_16009_new_n7139_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7140_));
AND2X2 AND2X2_2302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7132_), .B(AES_CORE_DATAPATH__abc_16009_new_n7142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7143_));
AND2X2 AND2X2_2303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7145_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7146_));
AND2X2 AND2X2_2304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7144_), .B(AES_CORE_DATAPATH__abc_16009_new_n7146_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7147_));
AND2X2 AND2X2_2305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7149_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7150_));
AND2X2 AND2X2_2306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7148_), .B(AES_CORE_DATAPATH__abc_16009_new_n7150_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7151_));
AND2X2 AND2X2_2307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7152_));
AND2X2 AND2X2_2308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7154_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7155_));
AND2X2 AND2X2_2309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4328_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7156_));
AND2X2 AND2X2_231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2683_));
AND2X2 AND2X2_2310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7158_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7159_));
AND2X2 AND2X2_2311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7161_));
AND2X2 AND2X2_2312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7162_));
AND2X2 AND2X2_2313 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7163_));
AND2X2 AND2X2_2314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7164_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7165_));
AND2X2 AND2X2_2315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4351_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7167_));
AND2X2 AND2X2_2316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7167_), .B(AES_CORE_DATAPATH__abc_16009_new_n7166_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7168_));
AND2X2 AND2X2_2317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7170_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7171_));
AND2X2 AND2X2_2318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7175_));
AND2X2 AND2X2_2319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7175_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7176_));
AND2X2 AND2X2_232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2686_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2687_));
AND2X2 AND2X2_2320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7177_));
AND2X2 AND2X2_2321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7180_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7181_));
AND2X2 AND2X2_2322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7179_), .B(AES_CORE_DATAPATH__abc_16009_new_n7181_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7182_));
AND2X2 AND2X2_2323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7183_));
AND2X2 AND2X2_2324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7185_), .B(AES_CORE_DATAPATH__abc_16009_new_n7186_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7187_));
AND2X2 AND2X2_2325 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7190_), .B(AES_CORE_DATAPATH__abc_16009_new_n7172_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7191_));
AND2X2 AND2X2_2326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7189_), .B(AES_CORE_DATAPATH__abc_16009_new_n7192_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7193_));
AND2X2 AND2X2_2327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7195_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7196_));
AND2X2 AND2X2_2328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7194_), .B(AES_CORE_DATAPATH__abc_16009_new_n7196_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7197_));
AND2X2 AND2X2_2329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7199_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7200_));
AND2X2 AND2X2_233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2685_), .B(AES_CORE_DATAPATH__abc_16009_new_n2687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2688_));
AND2X2 AND2X2_2330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7198_), .B(AES_CORE_DATAPATH__abc_16009_new_n7200_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7201_));
AND2X2 AND2X2_2331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7202_));
AND2X2 AND2X2_2332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7204_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7205_));
AND2X2 AND2X2_2333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4360_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7206_));
AND2X2 AND2X2_2334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7208_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7209_));
AND2X2 AND2X2_2335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7211_));
AND2X2 AND2X2_2336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7212_));
AND2X2 AND2X2_2337 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7213_));
AND2X2 AND2X2_2338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7214_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7215_));
AND2X2 AND2X2_2339 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4392_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7216_));
AND2X2 AND2X2_234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2689_));
AND2X2 AND2X2_2340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7217_));
AND2X2 AND2X2_2341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7219_));
AND2X2 AND2X2_2342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7219_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7220_));
AND2X2 AND2X2_2343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7221_));
AND2X2 AND2X2_2344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7224_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7225_));
AND2X2 AND2X2_2345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7223_), .B(AES_CORE_DATAPATH__abc_16009_new_n7225_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7226_));
AND2X2 AND2X2_2346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7227_));
AND2X2 AND2X2_2347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7229_), .B(AES_CORE_DATAPATH__abc_16009_new_n7230_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7231_));
AND2X2 AND2X2_2348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4383_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7234_));
AND2X2 AND2X2_2349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7234_), .B(AES_CORE_DATAPATH__abc_16009_new_n7233_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7235_));
AND2X2 AND2X2_235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2691_));
AND2X2 AND2X2_2350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7238_), .B(AES_CORE_DATAPATH__abc_16009_new_n7239_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7240_));
AND2X2 AND2X2_2351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7232_), .B(AES_CORE_DATAPATH__abc_16009_new_n7242_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7243_));
AND2X2 AND2X2_2352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7245_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7246_));
AND2X2 AND2X2_2353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7244_), .B(AES_CORE_DATAPATH__abc_16009_new_n7246_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7247_));
AND2X2 AND2X2_2354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7249_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7250_));
AND2X2 AND2X2_2355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7248_), .B(AES_CORE_DATAPATH__abc_16009_new_n7250_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7251_));
AND2X2 AND2X2_2356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7252_));
AND2X2 AND2X2_2357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7254_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7255_));
AND2X2 AND2X2_2358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4392_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7256_));
AND2X2 AND2X2_2359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7258_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7259_));
AND2X2 AND2X2_236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2691_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2692_));
AND2X2 AND2X2_2360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7261_));
AND2X2 AND2X2_2361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7262_));
AND2X2 AND2X2_2362 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7263_));
AND2X2 AND2X2_2363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7264_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7265_));
AND2X2 AND2X2_2364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4424_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7266_));
AND2X2 AND2X2_2365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7267_));
AND2X2 AND2X2_2366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7269_));
AND2X2 AND2X2_2367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7269_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7270_));
AND2X2 AND2X2_2368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7271_));
AND2X2 AND2X2_2369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7274_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7275_));
AND2X2 AND2X2_237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2693_));
AND2X2 AND2X2_2370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7273_), .B(AES_CORE_DATAPATH__abc_16009_new_n7275_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7276_));
AND2X2 AND2X2_2371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7277_));
AND2X2 AND2X2_2372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7279_), .B(AES_CORE_DATAPATH__abc_16009_new_n7280_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7281_));
AND2X2 AND2X2_2373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4415_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7284_));
AND2X2 AND2X2_2374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7284_), .B(AES_CORE_DATAPATH__abc_16009_new_n7283_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7285_));
AND2X2 AND2X2_2375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7288_), .B(AES_CORE_DATAPATH__abc_16009_new_n7289_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7290_));
AND2X2 AND2X2_2376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7282_), .B(AES_CORE_DATAPATH__abc_16009_new_n7292_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7293_));
AND2X2 AND2X2_2377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7295_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7296_));
AND2X2 AND2X2_2378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7294_), .B(AES_CORE_DATAPATH__abc_16009_new_n7296_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7297_));
AND2X2 AND2X2_2379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7299_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7300_));
AND2X2 AND2X2_238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2696_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2697_));
AND2X2 AND2X2_2380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7298_), .B(AES_CORE_DATAPATH__abc_16009_new_n7300_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7301_));
AND2X2 AND2X2_2381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7302_));
AND2X2 AND2X2_2382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7304_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7305_));
AND2X2 AND2X2_2383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4424_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7306_));
AND2X2 AND2X2_2384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7308_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7309_));
AND2X2 AND2X2_2385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5739_), .B(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7311_));
AND2X2 AND2X2_2386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7312_));
AND2X2 AND2X2_2387 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7313_));
AND2X2 AND2X2_2388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7314_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7315_));
AND2X2 AND2X2_2389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4447_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7317_));
AND2X2 AND2X2_239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2695_), .B(AES_CORE_DATAPATH__abc_16009_new_n2697_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2698_));
AND2X2 AND2X2_2390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7317_), .B(AES_CORE_DATAPATH__abc_16009_new_n7316_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7318_));
AND2X2 AND2X2_2391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7320_), .B(AES_CORE_DATAPATH__abc_16009_new_n5759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7321_));
AND2X2 AND2X2_2392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_bkp_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7325_));
AND2X2 AND2X2_2393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7325_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7326_));
AND2X2 AND2X2_2394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_bkp_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7327_));
AND2X2 AND2X2_2395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7330_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7331_));
AND2X2 AND2X2_2396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7329_), .B(AES_CORE_DATAPATH__abc_16009_new_n7331_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7332_));
AND2X2 AND2X2_2397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_bkp_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7333_));
AND2X2 AND2X2_2398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7335_), .B(AES_CORE_DATAPATH__abc_16009_new_n7336_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7337_));
AND2X2 AND2X2_2399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7340_), .B(AES_CORE_DATAPATH__abc_16009_new_n7322_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7341_));
AND2X2 AND2X2_24 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_));
AND2X2 AND2X2_240 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2699_));
AND2X2 AND2X2_2400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7339_), .B(AES_CORE_DATAPATH__abc_16009_new_n7342_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7343_));
AND2X2 AND2X2_2401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7345_), .B(AES_CORE_DATAPATH__abc_16009_new_n5793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7346_));
AND2X2 AND2X2_2402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7344_), .B(AES_CORE_DATAPATH__abc_16009_new_n7346_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7347_));
AND2X2 AND2X2_2403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7349_), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n7350_));
AND2X2 AND2X2_2404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7348_), .B(AES_CORE_DATAPATH__abc_16009_new_n7350_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7351_));
AND2X2 AND2X2_2405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7352_));
AND2X2 AND2X2_2406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7354_), .B(AES_CORE_DATAPATH__abc_16009_new_n5756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7355_));
AND2X2 AND2X2_2407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4456_), .B(AES_CORE_DATAPATH__abc_16009_new_n5754_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7356_));
AND2X2 AND2X2_2408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7358_), .B(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7359_));
AND2X2 AND2X2_2409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7361_));
AND2X2 AND2X2_241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2701_));
AND2X2 AND2X2_2410 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7362_));
AND2X2 AND2X2_2411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4561_), .B(AES_CORE_DATAPATH__abc_16009_new_n7365_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7366_));
AND2X2 AND2X2_2412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7364_), .B(AES_CORE_DATAPATH__abc_16009_new_n7366_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7367_));
AND2X2 AND2X2_2413 ( .A(\bus_in[0] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7368_));
AND2X2 AND2X2_2414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7369_));
AND2X2 AND2X2_2415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7372_), .B(AES_CORE_DATAPATH__abc_16009_new_n7371_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7373_));
AND2X2 AND2X2_2416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7374_), .B(AES_CORE_DATAPATH__abc_16009_new_n7376_), .Y(AES_CORE_DATAPATH__0key_3__31_0__0_));
AND2X2 AND2X2_2417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7379_));
AND2X2 AND2X2_2418 ( .A(\bus_in[1] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7380_));
AND2X2 AND2X2_2419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7378_), .B(AES_CORE_DATAPATH__abc_16009_new_n7382_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7383_));
AND2X2 AND2X2_242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2701_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2702_));
AND2X2 AND2X2_2420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7384_), .B(AES_CORE_DATAPATH__abc_16009_new_n7385_), .Y(AES_CORE_DATAPATH__0key_3__31_0__1_));
AND2X2 AND2X2_2421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7388_));
AND2X2 AND2X2_2422 ( .A(\bus_in[2] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7389_));
AND2X2 AND2X2_2423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7387_), .B(AES_CORE_DATAPATH__abc_16009_new_n7391_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7392_));
AND2X2 AND2X2_2424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7393_), .B(AES_CORE_DATAPATH__abc_16009_new_n7394_), .Y(AES_CORE_DATAPATH__0key_3__31_0__2_));
AND2X2 AND2X2_2425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7397_));
AND2X2 AND2X2_2426 ( .A(\bus_in[3] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7398_));
AND2X2 AND2X2_2427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7396_), .B(AES_CORE_DATAPATH__abc_16009_new_n7400_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7401_));
AND2X2 AND2X2_2428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7402_), .B(AES_CORE_DATAPATH__abc_16009_new_n7403_), .Y(AES_CORE_DATAPATH__0key_3__31_0__3_));
AND2X2 AND2X2_2429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7406_));
AND2X2 AND2X2_243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2703_));
AND2X2 AND2X2_2430 ( .A(\bus_in[4] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7407_));
AND2X2 AND2X2_2431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7405_), .B(AES_CORE_DATAPATH__abc_16009_new_n7409_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7410_));
AND2X2 AND2X2_2432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7410_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7411_));
AND2X2 AND2X2_2433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7412_));
AND2X2 AND2X2_2434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7415_));
AND2X2 AND2X2_2435 ( .A(\bus_in[5] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7416_));
AND2X2 AND2X2_2436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7414_), .B(AES_CORE_DATAPATH__abc_16009_new_n7418_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7419_));
AND2X2 AND2X2_2437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7419_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7420_));
AND2X2 AND2X2_2438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7421_));
AND2X2 AND2X2_2439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7424_));
AND2X2 AND2X2_244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2706_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2707_));
AND2X2 AND2X2_2440 ( .A(\bus_in[6] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7425_));
AND2X2 AND2X2_2441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7423_), .B(AES_CORE_DATAPATH__abc_16009_new_n7427_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7428_));
AND2X2 AND2X2_2442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7429_), .B(AES_CORE_DATAPATH__abc_16009_new_n7430_), .Y(AES_CORE_DATAPATH__0key_3__31_0__6_));
AND2X2 AND2X2_2443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7433_));
AND2X2 AND2X2_2444 ( .A(\bus_in[7] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7434_));
AND2X2 AND2X2_2445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7432_), .B(AES_CORE_DATAPATH__abc_16009_new_n7436_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7437_));
AND2X2 AND2X2_2446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7438_), .B(AES_CORE_DATAPATH__abc_16009_new_n7439_), .Y(AES_CORE_DATAPATH__0key_3__31_0__7_));
AND2X2 AND2X2_2447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7442_));
AND2X2 AND2X2_2448 ( .A(\bus_in[8] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7443_));
AND2X2 AND2X2_2449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7441_), .B(AES_CORE_DATAPATH__abc_16009_new_n7445_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7446_));
AND2X2 AND2X2_245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2705_), .B(AES_CORE_DATAPATH__abc_16009_new_n2707_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2708_));
AND2X2 AND2X2_2450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7446_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7447_));
AND2X2 AND2X2_2451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7448_));
AND2X2 AND2X2_2452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7451_));
AND2X2 AND2X2_2453 ( .A(\bus_in[9] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7452_));
AND2X2 AND2X2_2454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7450_), .B(AES_CORE_DATAPATH__abc_16009_new_n7454_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7455_));
AND2X2 AND2X2_2455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7455_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7456_));
AND2X2 AND2X2_2456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7457_));
AND2X2 AND2X2_2457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7460_));
AND2X2 AND2X2_2458 ( .A(\bus_in[10] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7461_));
AND2X2 AND2X2_2459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7459_), .B(AES_CORE_DATAPATH__abc_16009_new_n7463_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7464_));
AND2X2 AND2X2_246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2709_));
AND2X2 AND2X2_2460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7464_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7465_));
AND2X2 AND2X2_2461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7466_));
AND2X2 AND2X2_2462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7469_));
AND2X2 AND2X2_2463 ( .A(\bus_in[11] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7470_));
AND2X2 AND2X2_2464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7468_), .B(AES_CORE_DATAPATH__abc_16009_new_n7472_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7473_));
AND2X2 AND2X2_2465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7473_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7474_));
AND2X2 AND2X2_2466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7475_));
AND2X2 AND2X2_2467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7478_));
AND2X2 AND2X2_2468 ( .A(\bus_in[12] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7479_));
AND2X2 AND2X2_2469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7477_), .B(AES_CORE_DATAPATH__abc_16009_new_n7481_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7482_));
AND2X2 AND2X2_247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2711_));
AND2X2 AND2X2_2470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7482_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7483_));
AND2X2 AND2X2_2471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7484_));
AND2X2 AND2X2_2472 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7487_));
AND2X2 AND2X2_2473 ( .A(\bus_in[13] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7488_));
AND2X2 AND2X2_2474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7486_), .B(AES_CORE_DATAPATH__abc_16009_new_n7490_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7491_));
AND2X2 AND2X2_2475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7491_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7492_));
AND2X2 AND2X2_2476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7493_));
AND2X2 AND2X2_2477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7496_));
AND2X2 AND2X2_2478 ( .A(\bus_in[14] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7497_));
AND2X2 AND2X2_2479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7495_), .B(AES_CORE_DATAPATH__abc_16009_new_n7499_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7500_));
AND2X2 AND2X2_248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2711_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2712_));
AND2X2 AND2X2_2480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7500_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7501_));
AND2X2 AND2X2_2481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7502_));
AND2X2 AND2X2_2482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7505_));
AND2X2 AND2X2_2483 ( .A(\bus_in[15] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7506_));
AND2X2 AND2X2_2484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7504_), .B(AES_CORE_DATAPATH__abc_16009_new_n7508_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7509_));
AND2X2 AND2X2_2485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7509_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7510_));
AND2X2 AND2X2_2486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7511_));
AND2X2 AND2X2_2487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7514_));
AND2X2 AND2X2_2488 ( .A(\bus_in[16] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7515_));
AND2X2 AND2X2_2489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7513_), .B(AES_CORE_DATAPATH__abc_16009_new_n7517_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7518_));
AND2X2 AND2X2_249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2713_));
AND2X2 AND2X2_2490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7518_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7519_));
AND2X2 AND2X2_2491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7520_));
AND2X2 AND2X2_2492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7523_));
AND2X2 AND2X2_2493 ( .A(\bus_in[17] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7524_));
AND2X2 AND2X2_2494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7522_), .B(AES_CORE_DATAPATH__abc_16009_new_n7526_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7527_));
AND2X2 AND2X2_2495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7528_), .B(AES_CORE_DATAPATH__abc_16009_new_n7529_), .Y(AES_CORE_DATAPATH__0key_3__31_0__17_));
AND2X2 AND2X2_2496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7532_));
AND2X2 AND2X2_2497 ( .A(\bus_in[18] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7533_));
AND2X2 AND2X2_2498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7531_), .B(AES_CORE_DATAPATH__abc_16009_new_n7535_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7536_));
AND2X2 AND2X2_2499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7537_), .B(AES_CORE_DATAPATH__abc_16009_new_n7538_), .Y(AES_CORE_DATAPATH__0key_3__31_0__18_));
AND2X2 AND2X2_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n103_), .B(start), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_));
AND2X2 AND2X2_250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2716_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2717_));
AND2X2 AND2X2_2500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7541_));
AND2X2 AND2X2_2501 ( .A(\bus_in[19] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7542_));
AND2X2 AND2X2_2502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7540_), .B(AES_CORE_DATAPATH__abc_16009_new_n7544_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7545_));
AND2X2 AND2X2_2503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7546_), .B(AES_CORE_DATAPATH__abc_16009_new_n7547_), .Y(AES_CORE_DATAPATH__0key_3__31_0__19_));
AND2X2 AND2X2_2504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7550_));
AND2X2 AND2X2_2505 ( .A(\bus_in[20] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7551_));
AND2X2 AND2X2_2506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7549_), .B(AES_CORE_DATAPATH__abc_16009_new_n7553_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7554_));
AND2X2 AND2X2_2507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7554_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7555_));
AND2X2 AND2X2_2508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7556_));
AND2X2 AND2X2_2509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7559_));
AND2X2 AND2X2_251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2715_), .B(AES_CORE_DATAPATH__abc_16009_new_n2717_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2718_));
AND2X2 AND2X2_2510 ( .A(\bus_in[21] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7560_));
AND2X2 AND2X2_2511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7558_), .B(AES_CORE_DATAPATH__abc_16009_new_n7562_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7563_));
AND2X2 AND2X2_2512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7563_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7564_));
AND2X2 AND2X2_2513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7565_));
AND2X2 AND2X2_2514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7568_));
AND2X2 AND2X2_2515 ( .A(\bus_in[22] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7569_));
AND2X2 AND2X2_2516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7571_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7572_));
AND2X2 AND2X2_2517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7573_), .B(AES_CORE_DATAPATH__abc_16009_new_n7574_), .Y(AES_CORE_DATAPATH__0key_3__31_0__22_));
AND2X2 AND2X2_2518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7577_));
AND2X2 AND2X2_2519 ( .A(\bus_in[23] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7578_));
AND2X2 AND2X2_252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2719_));
AND2X2 AND2X2_2520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7576_), .B(AES_CORE_DATAPATH__abc_16009_new_n7580_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7581_));
AND2X2 AND2X2_2521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7582_), .B(AES_CORE_DATAPATH__abc_16009_new_n7583_), .Y(AES_CORE_DATAPATH__0key_3__31_0__23_));
AND2X2 AND2X2_2522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7586_));
AND2X2 AND2X2_2523 ( .A(\bus_in[24] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7587_));
AND2X2 AND2X2_2524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7585_), .B(AES_CORE_DATAPATH__abc_16009_new_n7589_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7590_));
AND2X2 AND2X2_2525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7591_), .B(AES_CORE_DATAPATH__abc_16009_new_n7592_), .Y(AES_CORE_DATAPATH__0key_3__31_0__24_));
AND2X2 AND2X2_2526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7595_));
AND2X2 AND2X2_2527 ( .A(\bus_in[25] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7596_));
AND2X2 AND2X2_2528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7594_), .B(AES_CORE_DATAPATH__abc_16009_new_n7598_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7599_));
AND2X2 AND2X2_2529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7600_), .B(AES_CORE_DATAPATH__abc_16009_new_n7601_), .Y(AES_CORE_DATAPATH__0key_3__31_0__25_));
AND2X2 AND2X2_253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2721_));
AND2X2 AND2X2_2530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7604_));
AND2X2 AND2X2_2531 ( .A(\bus_in[26] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7605_));
AND2X2 AND2X2_2532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7603_), .B(AES_CORE_DATAPATH__abc_16009_new_n7607_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7608_));
AND2X2 AND2X2_2533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7609_), .B(AES_CORE_DATAPATH__abc_16009_new_n7610_), .Y(AES_CORE_DATAPATH__0key_3__31_0__26_));
AND2X2 AND2X2_2534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7613_));
AND2X2 AND2X2_2535 ( .A(\bus_in[27] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7614_));
AND2X2 AND2X2_2536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7612_), .B(AES_CORE_DATAPATH__abc_16009_new_n7616_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7617_));
AND2X2 AND2X2_2537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7617_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7618_));
AND2X2 AND2X2_2538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7619_));
AND2X2 AND2X2_2539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7622_));
AND2X2 AND2X2_254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2721_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2722_));
AND2X2 AND2X2_2540 ( .A(\bus_in[28] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7623_));
AND2X2 AND2X2_2541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7621_), .B(AES_CORE_DATAPATH__abc_16009_new_n7625_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7626_));
AND2X2 AND2X2_2542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7626_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7627_));
AND2X2 AND2X2_2543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7628_));
AND2X2 AND2X2_2544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7631_));
AND2X2 AND2X2_2545 ( .A(\bus_in[29] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7632_));
AND2X2 AND2X2_2546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7630_), .B(AES_CORE_DATAPATH__abc_16009_new_n7634_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7635_));
AND2X2 AND2X2_2547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7636_), .B(AES_CORE_DATAPATH__abc_16009_new_n7637_), .Y(AES_CORE_DATAPATH__0key_3__31_0__29_));
AND2X2 AND2X2_2548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7640_));
AND2X2 AND2X2_2549 ( .A(\bus_in[30] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7641_));
AND2X2 AND2X2_255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2723_));
AND2X2 AND2X2_2550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7639_), .B(AES_CORE_DATAPATH__abc_16009_new_n7643_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7644_));
AND2X2 AND2X2_2551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7644_), .B(AES_CORE_DATAPATH__abc_16009_new_n7375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7645_));
AND2X2 AND2X2_2552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7646_));
AND2X2 AND2X2_2553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7365_), .B(AES_CORE_DATAPATH_key_host_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7649_));
AND2X2 AND2X2_2554 ( .A(\bus_in[31] ), .B(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7650_));
AND2X2 AND2X2_2555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7648_), .B(AES_CORE_DATAPATH__abc_16009_new_n7652_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7653_));
AND2X2 AND2X2_2556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7654_), .B(AES_CORE_DATAPATH__abc_16009_new_n7655_), .Y(AES_CORE_DATAPATH__0key_3__31_0__31_));
AND2X2 AND2X2_2557 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7657_));
AND2X2 AND2X2_2558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7370_), .B(AES_CORE_DATAPATH__abc_16009_new_n5155_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7658_));
AND2X2 AND2X2_2559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7660_), .B(AES_CORE_DATAPATH__abc_16009_new_n7661_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__1_));
AND2X2 AND2X2_256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2726_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2727_));
AND2X2 AND2X2_2560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7663_), .B(AES_CORE_DATAPATH__abc_16009_new_n7664_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__2_));
AND2X2 AND2X2_2561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7666_), .B(AES_CORE_DATAPATH__abc_16009_new_n7667_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__3_));
AND2X2 AND2X2_2562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7669_), .B(AES_CORE_DATAPATH__abc_16009_new_n7670_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__4_));
AND2X2 AND2X2_2563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7672_), .B(AES_CORE_DATAPATH__abc_16009_new_n7673_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__5_));
AND2X2 AND2X2_2564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7675_), .B(AES_CORE_DATAPATH__abc_16009_new_n7676_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__6_));
AND2X2 AND2X2_2565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7678_), .B(AES_CORE_DATAPATH__abc_16009_new_n7679_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__7_));
AND2X2 AND2X2_2566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7681_), .B(AES_CORE_DATAPATH__abc_16009_new_n7682_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__8_));
AND2X2 AND2X2_2567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7684_), .B(AES_CORE_DATAPATH__abc_16009_new_n7685_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__9_));
AND2X2 AND2X2_2568 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7687_), .B(AES_CORE_DATAPATH__abc_16009_new_n7688_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__10_));
AND2X2 AND2X2_2569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7690_), .B(AES_CORE_DATAPATH__abc_16009_new_n7691_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__11_));
AND2X2 AND2X2_257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2725_), .B(AES_CORE_DATAPATH__abc_16009_new_n2727_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2728_));
AND2X2 AND2X2_2570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7693_), .B(AES_CORE_DATAPATH__abc_16009_new_n7694_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__12_));
AND2X2 AND2X2_2571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7696_), .B(AES_CORE_DATAPATH__abc_16009_new_n7697_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__13_));
AND2X2 AND2X2_2572 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7699_), .B(AES_CORE_DATAPATH__abc_16009_new_n7700_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__14_));
AND2X2 AND2X2_2573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7702_), .B(AES_CORE_DATAPATH__abc_16009_new_n7703_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__15_));
AND2X2 AND2X2_2574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7705_), .B(AES_CORE_DATAPATH__abc_16009_new_n7706_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__16_));
AND2X2 AND2X2_2575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7708_), .B(AES_CORE_DATAPATH__abc_16009_new_n7709_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__17_));
AND2X2 AND2X2_2576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7711_), .B(AES_CORE_DATAPATH__abc_16009_new_n7712_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__18_));
AND2X2 AND2X2_2577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7714_), .B(AES_CORE_DATAPATH__abc_16009_new_n7715_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__19_));
AND2X2 AND2X2_2578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7717_), .B(AES_CORE_DATAPATH__abc_16009_new_n7718_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__20_));
AND2X2 AND2X2_2579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7720_), .B(AES_CORE_DATAPATH__abc_16009_new_n7721_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__21_));
AND2X2 AND2X2_258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2729_));
AND2X2 AND2X2_2580 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7723_), .B(AES_CORE_DATAPATH__abc_16009_new_n7724_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__22_));
AND2X2 AND2X2_2581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7726_), .B(AES_CORE_DATAPATH__abc_16009_new_n7727_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__23_));
AND2X2 AND2X2_2582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7729_), .B(AES_CORE_DATAPATH__abc_16009_new_n7730_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__24_));
AND2X2 AND2X2_2583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7732_), .B(AES_CORE_DATAPATH__abc_16009_new_n7733_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__25_));
AND2X2 AND2X2_2584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7735_), .B(AES_CORE_DATAPATH__abc_16009_new_n7736_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__26_));
AND2X2 AND2X2_2585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7738_), .B(AES_CORE_DATAPATH__abc_16009_new_n7739_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__27_));
AND2X2 AND2X2_2586 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7741_), .B(AES_CORE_DATAPATH__abc_16009_new_n7742_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__28_));
AND2X2 AND2X2_2587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7744_), .B(AES_CORE_DATAPATH__abc_16009_new_n7745_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__29_));
AND2X2 AND2X2_2588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7747_), .B(AES_CORE_DATAPATH__abc_16009_new_n7748_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__30_));
AND2X2 AND2X2_2589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7751_), .B(AES_CORE_DATAPATH__abc_16009_new_n7750_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__31_));
AND2X2 AND2X2_259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2731_));
AND2X2 AND2X2_2590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7754_));
AND2X2 AND2X2_2591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7755_));
AND2X2 AND2X2_2592 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7756_));
AND2X2 AND2X2_2593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7758_));
AND2X2 AND2X2_2594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7759_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7760_));
AND2X2 AND2X2_2595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7762_));
AND2X2 AND2X2_2596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7763_));
AND2X2 AND2X2_2597 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7764_));
AND2X2 AND2X2_2598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7765_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7766_));
AND2X2 AND2X2_2599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7767_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7768_));
AND2X2 AND2X2_26 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n105_));
AND2X2 AND2X2_260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2731_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2732_));
AND2X2 AND2X2_2600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7770_));
AND2X2 AND2X2_2601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7771_));
AND2X2 AND2X2_2602 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7772_));
AND2X2 AND2X2_2603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7773_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7774_));
AND2X2 AND2X2_2604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7775_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7776_));
AND2X2 AND2X2_2605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7778_));
AND2X2 AND2X2_2606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7779_));
AND2X2 AND2X2_2607 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7780_));
AND2X2 AND2X2_2608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7781_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7782_));
AND2X2 AND2X2_2609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7783_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7784_));
AND2X2 AND2X2_261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2733_));
AND2X2 AND2X2_2610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7786_));
AND2X2 AND2X2_2611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7787_));
AND2X2 AND2X2_2612 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7788_));
AND2X2 AND2X2_2613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7789_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7790_));
AND2X2 AND2X2_2614 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7791_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7792_));
AND2X2 AND2X2_2615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7794_));
AND2X2 AND2X2_2616 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7795_));
AND2X2 AND2X2_2617 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7796_));
AND2X2 AND2X2_2618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7797_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7798_));
AND2X2 AND2X2_2619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7799_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7800_));
AND2X2 AND2X2_262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2736_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2737_));
AND2X2 AND2X2_2620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7802_));
AND2X2 AND2X2_2621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7803_));
AND2X2 AND2X2_2622 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7804_));
AND2X2 AND2X2_2623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7806_));
AND2X2 AND2X2_2624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7807_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7808_));
AND2X2 AND2X2_2625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7810_));
AND2X2 AND2X2_2626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7811_));
AND2X2 AND2X2_2627 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7812_));
AND2X2 AND2X2_2628 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7814_));
AND2X2 AND2X2_2629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7815_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7816_));
AND2X2 AND2X2_263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2735_), .B(AES_CORE_DATAPATH__abc_16009_new_n2737_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2738_));
AND2X2 AND2X2_2630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7818_));
AND2X2 AND2X2_2631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7819_));
AND2X2 AND2X2_2632 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7820_));
AND2X2 AND2X2_2633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7821_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7822_));
AND2X2 AND2X2_2634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7823_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7824_));
AND2X2 AND2X2_2635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7826_));
AND2X2 AND2X2_2636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7827_));
AND2X2 AND2X2_2637 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7828_));
AND2X2 AND2X2_2638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7829_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7830_));
AND2X2 AND2X2_2639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7831_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7832_));
AND2X2 AND2X2_264 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2739_));
AND2X2 AND2X2_2640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7834_));
AND2X2 AND2X2_2641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7835_));
AND2X2 AND2X2_2642 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7836_));
AND2X2 AND2X2_2643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7837_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7838_));
AND2X2 AND2X2_2644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7839_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7840_));
AND2X2 AND2X2_2645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7842_));
AND2X2 AND2X2_2646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7843_));
AND2X2 AND2X2_2647 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7844_));
AND2X2 AND2X2_2648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7845_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7846_));
AND2X2 AND2X2_2649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7847_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7848_));
AND2X2 AND2X2_265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2741_));
AND2X2 AND2X2_2650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7850_));
AND2X2 AND2X2_2651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7851_));
AND2X2 AND2X2_2652 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7852_));
AND2X2 AND2X2_2653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7853_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7854_));
AND2X2 AND2X2_2654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7855_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7856_));
AND2X2 AND2X2_2655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7858_));
AND2X2 AND2X2_2656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7859_));
AND2X2 AND2X2_2657 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7860_));
AND2X2 AND2X2_2658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7861_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7862_));
AND2X2 AND2X2_2659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7863_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7864_));
AND2X2 AND2X2_266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2741_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2742_));
AND2X2 AND2X2_2660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7866_));
AND2X2 AND2X2_2661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7867_));
AND2X2 AND2X2_2662 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7868_));
AND2X2 AND2X2_2663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7869_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7870_));
AND2X2 AND2X2_2664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7871_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7872_));
AND2X2 AND2X2_2665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7874_));
AND2X2 AND2X2_2666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7875_));
AND2X2 AND2X2_2667 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7876_));
AND2X2 AND2X2_2668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7877_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7878_));
AND2X2 AND2X2_2669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7879_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7880_));
AND2X2 AND2X2_267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2743_));
AND2X2 AND2X2_2670 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7882_));
AND2X2 AND2X2_2671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7883_));
AND2X2 AND2X2_2672 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7884_));
AND2X2 AND2X2_2673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7885_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7886_));
AND2X2 AND2X2_2674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7887_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7888_));
AND2X2 AND2X2_2675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7890_));
AND2X2 AND2X2_2676 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7891_));
AND2X2 AND2X2_2677 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7892_));
AND2X2 AND2X2_2678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7893_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7894_));
AND2X2 AND2X2_2679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7895_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7896_));
AND2X2 AND2X2_268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2746_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2747_));
AND2X2 AND2X2_2680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7898_));
AND2X2 AND2X2_2681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7899_));
AND2X2 AND2X2_2682 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7900_));
AND2X2 AND2X2_2683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7901_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7902_));
AND2X2 AND2X2_2684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7903_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7904_));
AND2X2 AND2X2_2685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7906_));
AND2X2 AND2X2_2686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7907_));
AND2X2 AND2X2_2687 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7908_));
AND2X2 AND2X2_2688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7909_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7910_));
AND2X2 AND2X2_2689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7911_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7912_));
AND2X2 AND2X2_269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2745_), .B(AES_CORE_DATAPATH__abc_16009_new_n2747_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2748_));
AND2X2 AND2X2_2690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7914_));
AND2X2 AND2X2_2691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7915_));
AND2X2 AND2X2_2692 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7916_));
AND2X2 AND2X2_2693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7918_));
AND2X2 AND2X2_2694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7919_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7920_));
AND2X2 AND2X2_2695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7922_));
AND2X2 AND2X2_2696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7923_));
AND2X2 AND2X2_2697 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7924_));
AND2X2 AND2X2_2698 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7925_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7926_));
AND2X2 AND2X2_2699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7927_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7928_));
AND2X2 AND2X2_27 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n105_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n102_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n106_));
AND2X2 AND2X2_270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2749_));
AND2X2 AND2X2_2700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7930_));
AND2X2 AND2X2_2701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7931_));
AND2X2 AND2X2_2702 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7932_));
AND2X2 AND2X2_2703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7934_));
AND2X2 AND2X2_2704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7935_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7936_));
AND2X2 AND2X2_2705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7938_));
AND2X2 AND2X2_2706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7939_));
AND2X2 AND2X2_2707 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7940_));
AND2X2 AND2X2_2708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7941_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7942_));
AND2X2 AND2X2_2709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7943_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7944_));
AND2X2 AND2X2_271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2751_));
AND2X2 AND2X2_2710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7946_));
AND2X2 AND2X2_2711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7947_));
AND2X2 AND2X2_2712 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7948_));
AND2X2 AND2X2_2713 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7949_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7950_));
AND2X2 AND2X2_2714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7951_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7952_));
AND2X2 AND2X2_2715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7954_));
AND2X2 AND2X2_2716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7955_));
AND2X2 AND2X2_2717 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7956_));
AND2X2 AND2X2_2718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7957_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7958_));
AND2X2 AND2X2_2719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7959_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7960_));
AND2X2 AND2X2_272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2751_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2752_));
AND2X2 AND2X2_2720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7962_));
AND2X2 AND2X2_2721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7963_));
AND2X2 AND2X2_2722 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7964_));
AND2X2 AND2X2_2723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7965_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7966_));
AND2X2 AND2X2_2724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7967_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7968_));
AND2X2 AND2X2_2725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7970_));
AND2X2 AND2X2_2726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7971_));
AND2X2 AND2X2_2727 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7972_));
AND2X2 AND2X2_2728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7973_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7974_));
AND2X2 AND2X2_2729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7975_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7976_));
AND2X2 AND2X2_273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2753_));
AND2X2 AND2X2_2730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7978_));
AND2X2 AND2X2_2731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7979_));
AND2X2 AND2X2_2732 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7980_));
AND2X2 AND2X2_2733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7981_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7982_));
AND2X2 AND2X2_2734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7983_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7984_));
AND2X2 AND2X2_2735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7986_));
AND2X2 AND2X2_2736 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7987_));
AND2X2 AND2X2_2737 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7988_));
AND2X2 AND2X2_2738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7989_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7990_));
AND2X2 AND2X2_2739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7991_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7992_));
AND2X2 AND2X2_274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2756_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2757_));
AND2X2 AND2X2_2740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7994_));
AND2X2 AND2X2_2741 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7995_));
AND2X2 AND2X2_2742 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7996_));
AND2X2 AND2X2_2743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n7997_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7998_));
AND2X2 AND2X2_2744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7999_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8000_));
AND2X2 AND2X2_2745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7753_), .B(AES_CORE_DATAPATH_col_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8002_));
AND2X2 AND2X2_2746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8003_));
AND2X2 AND2X2_2747 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8004_));
AND2X2 AND2X2_2748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8005_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8006_));
AND2X2 AND2X2_2749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8007_), .B(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8008_));
AND2X2 AND2X2_275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2755_), .B(AES_CORE_DATAPATH__abc_16009_new_n2757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2758_));
AND2X2 AND2X2_2750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8011_));
AND2X2 AND2X2_2751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8012_));
AND2X2 AND2X2_2752 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8013_));
AND2X2 AND2X2_2753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8015_));
AND2X2 AND2X2_2754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8016_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8017_));
AND2X2 AND2X2_2755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8019_));
AND2X2 AND2X2_2756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8020_));
AND2X2 AND2X2_2757 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8021_));
AND2X2 AND2X2_2758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8022_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8023_));
AND2X2 AND2X2_2759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8024_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8025_));
AND2X2 AND2X2_276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2759_));
AND2X2 AND2X2_2760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8027_));
AND2X2 AND2X2_2761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8028_));
AND2X2 AND2X2_2762 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8029_));
AND2X2 AND2X2_2763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8031_));
AND2X2 AND2X2_2764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8032_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8033_));
AND2X2 AND2X2_2765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8035_));
AND2X2 AND2X2_2766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8036_));
AND2X2 AND2X2_2767 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8037_));
AND2X2 AND2X2_2768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8038_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8039_));
AND2X2 AND2X2_2769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8040_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8041_));
AND2X2 AND2X2_277 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2761_));
AND2X2 AND2X2_2770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8043_));
AND2X2 AND2X2_2771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8044_));
AND2X2 AND2X2_2772 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8045_));
AND2X2 AND2X2_2773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8046_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8047_));
AND2X2 AND2X2_2774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8048_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8049_));
AND2X2 AND2X2_2775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8051_));
AND2X2 AND2X2_2776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8052_));
AND2X2 AND2X2_2777 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8053_));
AND2X2 AND2X2_2778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8054_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8055_));
AND2X2 AND2X2_2779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8056_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8057_));
AND2X2 AND2X2_278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2761_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2762_));
AND2X2 AND2X2_2780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8059_));
AND2X2 AND2X2_2781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8060_));
AND2X2 AND2X2_2782 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8061_));
AND2X2 AND2X2_2783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8062_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8063_));
AND2X2 AND2X2_2784 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8064_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8065_));
AND2X2 AND2X2_2785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8067_));
AND2X2 AND2X2_2786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8068_));
AND2X2 AND2X2_2787 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8069_));
AND2X2 AND2X2_2788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8070_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8071_));
AND2X2 AND2X2_2789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8072_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8073_));
AND2X2 AND2X2_279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2763_));
AND2X2 AND2X2_2790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8075_));
AND2X2 AND2X2_2791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8076_));
AND2X2 AND2X2_2792 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8077_));
AND2X2 AND2X2_2793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8078_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8079_));
AND2X2 AND2X2_2794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8080_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8081_));
AND2X2 AND2X2_2795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8083_));
AND2X2 AND2X2_2796 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8084_));
AND2X2 AND2X2_2797 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8085_));
AND2X2 AND2X2_2798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8087_));
AND2X2 AND2X2_2799 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8088_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8089_));
AND2X2 AND2X2_28 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_));
AND2X2 AND2X2_280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2766_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2767_));
AND2X2 AND2X2_2800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8091_));
AND2X2 AND2X2_2801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8092_));
AND2X2 AND2X2_2802 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8093_));
AND2X2 AND2X2_2803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8094_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8095_));
AND2X2 AND2X2_2804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8096_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8097_));
AND2X2 AND2X2_2805 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8099_));
AND2X2 AND2X2_2806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8100_));
AND2X2 AND2X2_2807 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8101_));
AND2X2 AND2X2_2808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8103_));
AND2X2 AND2X2_2809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8104_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8105_));
AND2X2 AND2X2_281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2765_), .B(AES_CORE_DATAPATH__abc_16009_new_n2767_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2768_));
AND2X2 AND2X2_2810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8107_));
AND2X2 AND2X2_2811 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8108_));
AND2X2 AND2X2_2812 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8109_));
AND2X2 AND2X2_2813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8111_));
AND2X2 AND2X2_2814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8112_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8113_));
AND2X2 AND2X2_2815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8115_));
AND2X2 AND2X2_2816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8116_));
AND2X2 AND2X2_2817 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8117_));
AND2X2 AND2X2_2818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8118_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8119_));
AND2X2 AND2X2_2819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8120_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8121_));
AND2X2 AND2X2_282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2769_));
AND2X2 AND2X2_2820 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8123_));
AND2X2 AND2X2_2821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8124_));
AND2X2 AND2X2_2822 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8125_));
AND2X2 AND2X2_2823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8127_));
AND2X2 AND2X2_2824 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8128_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8129_));
AND2X2 AND2X2_2825 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8131_));
AND2X2 AND2X2_2826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8132_));
AND2X2 AND2X2_2827 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8133_));
AND2X2 AND2X2_2828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8134_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8135_));
AND2X2 AND2X2_2829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8136_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8137_));
AND2X2 AND2X2_283 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2771_));
AND2X2 AND2X2_2830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8139_));
AND2X2 AND2X2_2831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8140_));
AND2X2 AND2X2_2832 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8141_));
AND2X2 AND2X2_2833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8143_));
AND2X2 AND2X2_2834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8144_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8145_));
AND2X2 AND2X2_2835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8147_));
AND2X2 AND2X2_2836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8148_));
AND2X2 AND2X2_2837 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8149_));
AND2X2 AND2X2_2838 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8150_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8151_));
AND2X2 AND2X2_2839 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8152_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8153_));
AND2X2 AND2X2_284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2771_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2772_));
AND2X2 AND2X2_2840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8155_));
AND2X2 AND2X2_2841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8156_));
AND2X2 AND2X2_2842 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8157_));
AND2X2 AND2X2_2843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8158_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8159_));
AND2X2 AND2X2_2844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8160_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8161_));
AND2X2 AND2X2_2845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8163_));
AND2X2 AND2X2_2846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8164_));
AND2X2 AND2X2_2847 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8165_));
AND2X2 AND2X2_2848 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8166_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8167_));
AND2X2 AND2X2_2849 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8168_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8169_));
AND2X2 AND2X2_285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2773_));
AND2X2 AND2X2_2850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8171_));
AND2X2 AND2X2_2851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8172_));
AND2X2 AND2X2_2852 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8173_));
AND2X2 AND2X2_2853 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8174_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8175_));
AND2X2 AND2X2_2854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8176_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8177_));
AND2X2 AND2X2_2855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8179_));
AND2X2 AND2X2_2856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8180_));
AND2X2 AND2X2_2857 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8181_));
AND2X2 AND2X2_2858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8182_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8183_));
AND2X2 AND2X2_2859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8184_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8185_));
AND2X2 AND2X2_286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2776_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2777_));
AND2X2 AND2X2_2860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8187_));
AND2X2 AND2X2_2861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8188_));
AND2X2 AND2X2_2862 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8189_));
AND2X2 AND2X2_2863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8190_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8191_));
AND2X2 AND2X2_2864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8192_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8193_));
AND2X2 AND2X2_2865 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8195_));
AND2X2 AND2X2_2866 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8196_));
AND2X2 AND2X2_2867 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8197_));
AND2X2 AND2X2_2868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8198_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8199_));
AND2X2 AND2X2_2869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8200_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8201_));
AND2X2 AND2X2_287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2775_), .B(AES_CORE_DATAPATH__abc_16009_new_n2777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2778_));
AND2X2 AND2X2_2870 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8203_));
AND2X2 AND2X2_2871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8204_));
AND2X2 AND2X2_2872 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8205_));
AND2X2 AND2X2_2873 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8206_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8207_));
AND2X2 AND2X2_2874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8208_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8209_));
AND2X2 AND2X2_2875 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8211_));
AND2X2 AND2X2_2876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8212_));
AND2X2 AND2X2_2877 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8213_));
AND2X2 AND2X2_2878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8214_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8215_));
AND2X2 AND2X2_2879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8216_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8217_));
AND2X2 AND2X2_288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2779_));
AND2X2 AND2X2_2880 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8219_));
AND2X2 AND2X2_2881 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8220_));
AND2X2 AND2X2_2882 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8221_));
AND2X2 AND2X2_2883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8222_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8223_));
AND2X2 AND2X2_2884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8224_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8225_));
AND2X2 AND2X2_2885 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8227_));
AND2X2 AND2X2_2886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8228_));
AND2X2 AND2X2_2887 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8229_));
AND2X2 AND2X2_2888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8230_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8231_));
AND2X2 AND2X2_2889 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8232_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8233_));
AND2X2 AND2X2_289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2781_));
AND2X2 AND2X2_2890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8235_));
AND2X2 AND2X2_2891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8236_));
AND2X2 AND2X2_2892 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8237_));
AND2X2 AND2X2_2893 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8238_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8239_));
AND2X2 AND2X2_2894 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8240_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8241_));
AND2X2 AND2X2_2895 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8243_));
AND2X2 AND2X2_2896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8244_));
AND2X2 AND2X2_2897 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8245_));
AND2X2 AND2X2_2898 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8246_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8247_));
AND2X2 AND2X2_2899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8248_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8249_));
AND2X2 AND2X2_29 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT_state_12_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n108_));
AND2X2 AND2X2_290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2781_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2782_));
AND2X2 AND2X2_2900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8251_));
AND2X2 AND2X2_2901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8252_));
AND2X2 AND2X2_2902 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8253_));
AND2X2 AND2X2_2903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8254_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8255_));
AND2X2 AND2X2_2904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8256_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8257_));
AND2X2 AND2X2_2905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8010_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8259_));
AND2X2 AND2X2_2906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8260_));
AND2X2 AND2X2_2907 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8261_));
AND2X2 AND2X2_2908 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8262_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8263_));
AND2X2 AND2X2_2909 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8264_), .B(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8265_));
AND2X2 AND2X2_291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2783_));
AND2X2 AND2X2_2910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8268_));
AND2X2 AND2X2_2911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8269_));
AND2X2 AND2X2_2912 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8270_));
AND2X2 AND2X2_2913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8271_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8272_));
AND2X2 AND2X2_2914 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8273_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8274_));
AND2X2 AND2X2_2915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8276_));
AND2X2 AND2X2_2916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8277_));
AND2X2 AND2X2_2917 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8278_));
AND2X2 AND2X2_2918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8279_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8280_));
AND2X2 AND2X2_2919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8281_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8282_));
AND2X2 AND2X2_292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2786_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2787_));
AND2X2 AND2X2_2920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8284_));
AND2X2 AND2X2_2921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8285_));
AND2X2 AND2X2_2922 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8286_));
AND2X2 AND2X2_2923 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8287_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8288_));
AND2X2 AND2X2_2924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8289_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8290_));
AND2X2 AND2X2_2925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8292_));
AND2X2 AND2X2_2926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8293_));
AND2X2 AND2X2_2927 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8294_));
AND2X2 AND2X2_2928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8295_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8296_));
AND2X2 AND2X2_2929 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8297_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8298_));
AND2X2 AND2X2_293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2785_), .B(AES_CORE_DATAPATH__abc_16009_new_n2787_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2788_));
AND2X2 AND2X2_2930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8300_));
AND2X2 AND2X2_2931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8301_));
AND2X2 AND2X2_2932 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8302_));
AND2X2 AND2X2_2933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8303_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8304_));
AND2X2 AND2X2_2934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8305_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8306_));
AND2X2 AND2X2_2935 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8308_));
AND2X2 AND2X2_2936 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8309_));
AND2X2 AND2X2_2937 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8310_));
AND2X2 AND2X2_2938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8311_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8312_));
AND2X2 AND2X2_2939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8313_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8314_));
AND2X2 AND2X2_294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2789_));
AND2X2 AND2X2_2940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8316_));
AND2X2 AND2X2_2941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8317_));
AND2X2 AND2X2_2942 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8318_));
AND2X2 AND2X2_2943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8319_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8320_));
AND2X2 AND2X2_2944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8321_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8322_));
AND2X2 AND2X2_2945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8324_));
AND2X2 AND2X2_2946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8325_));
AND2X2 AND2X2_2947 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8326_));
AND2X2 AND2X2_2948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8327_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8328_));
AND2X2 AND2X2_2949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8329_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8330_));
AND2X2 AND2X2_295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2472_), .B(AES_CORE_DATAPATH_iv_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2791_));
AND2X2 AND2X2_2950 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8332_));
AND2X2 AND2X2_2951 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8333_));
AND2X2 AND2X2_2952 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8334_));
AND2X2 AND2X2_2953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8335_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8336_));
AND2X2 AND2X2_2954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8337_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8338_));
AND2X2 AND2X2_2955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8340_));
AND2X2 AND2X2_2956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8341_));
AND2X2 AND2X2_2957 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8342_));
AND2X2 AND2X2_2958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8343_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8344_));
AND2X2 AND2X2_2959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8345_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8346_));
AND2X2 AND2X2_296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2791_), .B(AES_CORE_DATAPATH__abc_16009_new_n2475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2792_));
AND2X2 AND2X2_2960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8348_));
AND2X2 AND2X2_2961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8349_));
AND2X2 AND2X2_2962 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8350_));
AND2X2 AND2X2_2963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8351_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8352_));
AND2X2 AND2X2_2964 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8353_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8354_));
AND2X2 AND2X2_2965 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8356_));
AND2X2 AND2X2_2966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8357_));
AND2X2 AND2X2_2967 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8358_));
AND2X2 AND2X2_2968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8359_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8360_));
AND2X2 AND2X2_2969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8361_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8362_));
AND2X2 AND2X2_297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .B(AES_CORE_DATAPATH_iv_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2793_));
AND2X2 AND2X2_2970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8364_));
AND2X2 AND2X2_2971 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8365_));
AND2X2 AND2X2_2972 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8366_));
AND2X2 AND2X2_2973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8368_));
AND2X2 AND2X2_2974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8369_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8370_));
AND2X2 AND2X2_2975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8372_));
AND2X2 AND2X2_2976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8373_));
AND2X2 AND2X2_2977 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8374_));
AND2X2 AND2X2_2978 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8376_));
AND2X2 AND2X2_2979 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8377_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8378_));
AND2X2 AND2X2_298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2796_), .B(AES_CORE_DATAPATH__abc_16009_new_n2484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2797_));
AND2X2 AND2X2_2980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8380_));
AND2X2 AND2X2_2981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8381_));
AND2X2 AND2X2_2982 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8382_));
AND2X2 AND2X2_2983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8383_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8384_));
AND2X2 AND2X2_2984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8385_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8386_));
AND2X2 AND2X2_2985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8388_));
AND2X2 AND2X2_2986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8389_));
AND2X2 AND2X2_2987 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8390_));
AND2X2 AND2X2_2988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8391_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8392_));
AND2X2 AND2X2_2989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8393_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8394_));
AND2X2 AND2X2_299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2795_), .B(AES_CORE_DATAPATH__abc_16009_new_n2797_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2798_));
AND2X2 AND2X2_2990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8396_));
AND2X2 AND2X2_2991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8397_));
AND2X2 AND2X2_2992 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8398_));
AND2X2 AND2X2_2993 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8399_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8400_));
AND2X2 AND2X2_2994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8401_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8402_));
AND2X2 AND2X2_2995 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8404_));
AND2X2 AND2X2_2996 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8405_));
AND2X2 AND2X2_2997 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8406_));
AND2X2 AND2X2_2998 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8407_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8408_));
AND2X2 AND2X2_2999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8409_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8410_));
AND2X2 AND2X2_3 ( .A(\addr[0] ), .B(write_en), .Y(_abc_15574_new_n15_));
AND2X2 AND2X2_30 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_));
AND2X2 AND2X2_300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2799_));
AND2X2 AND2X2_3000 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8412_));
AND2X2 AND2X2_3001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8413_));
AND2X2 AND2X2_3002 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8414_));
AND2X2 AND2X2_3003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8415_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8416_));
AND2X2 AND2X2_3004 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8417_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8418_));
AND2X2 AND2X2_3005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8420_));
AND2X2 AND2X2_3006 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8421_));
AND2X2 AND2X2_3007 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8422_));
AND2X2 AND2X2_3008 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8423_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8424_));
AND2X2 AND2X2_3009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8425_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8426_));
AND2X2 AND2X2_301 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2803_));
AND2X2 AND2X2_3010 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8428_));
AND2X2 AND2X2_3011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8429_));
AND2X2 AND2X2_3012 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8430_));
AND2X2 AND2X2_3013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8431_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8432_));
AND2X2 AND2X2_3014 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8433_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8434_));
AND2X2 AND2X2_3015 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8436_));
AND2X2 AND2X2_3016 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8437_));
AND2X2 AND2X2_3017 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8438_));
AND2X2 AND2X2_3018 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8439_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8440_));
AND2X2 AND2X2_3019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8441_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8442_));
AND2X2 AND2X2_302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2808_));
AND2X2 AND2X2_3020 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8444_));
AND2X2 AND2X2_3021 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8445_));
AND2X2 AND2X2_3022 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8446_));
AND2X2 AND2X2_3023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8447_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8448_));
AND2X2 AND2X2_3024 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8449_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8450_));
AND2X2 AND2X2_3025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8452_));
AND2X2 AND2X2_3026 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8453_));
AND2X2 AND2X2_3027 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8454_));
AND2X2 AND2X2_3028 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8456_));
AND2X2 AND2X2_3029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8457_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8458_));
AND2X2 AND2X2_303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2809_));
AND2X2 AND2X2_3030 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8460_));
AND2X2 AND2X2_3031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8461_));
AND2X2 AND2X2_3032 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8462_));
AND2X2 AND2X2_3033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8463_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8464_));
AND2X2 AND2X2_3034 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8465_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8466_));
AND2X2 AND2X2_3035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8468_));
AND2X2 AND2X2_3036 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8469_));
AND2X2 AND2X2_3037 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8470_));
AND2X2 AND2X2_3038 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8472_));
AND2X2 AND2X2_3039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8473_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8474_));
AND2X2 AND2X2_304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2810_), .B(AES_CORE_DATAPATH__abc_16009_new_n2807_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2811_));
AND2X2 AND2X2_3040 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8476_));
AND2X2 AND2X2_3041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8477_));
AND2X2 AND2X2_3042 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8478_));
AND2X2 AND2X2_3043 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8479_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8480_));
AND2X2 AND2X2_3044 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8481_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8482_));
AND2X2 AND2X2_3045 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8484_));
AND2X2 AND2X2_3046 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8485_));
AND2X2 AND2X2_3047 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8486_));
AND2X2 AND2X2_3048 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8487_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8488_));
AND2X2 AND2X2_3049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8489_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8490_));
AND2X2 AND2X2_305 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_out_sel_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2812_));
AND2X2 AND2X2_3050 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8492_));
AND2X2 AND2X2_3051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8493_));
AND2X2 AND2X2_3052 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8494_));
AND2X2 AND2X2_3053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8495_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8496_));
AND2X2 AND2X2_3054 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8497_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8498_));
AND2X2 AND2X2_3055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8500_));
AND2X2 AND2X2_3056 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8501_));
AND2X2 AND2X2_3057 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8502_));
AND2X2 AND2X2_3058 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8503_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8504_));
AND2X2 AND2X2_3059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8505_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8506_));
AND2X2 AND2X2_306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2815_));
AND2X2 AND2X2_3060 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8508_));
AND2X2 AND2X2_3061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8509_));
AND2X2 AND2X2_3062 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8510_));
AND2X2 AND2X2_3063 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8511_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8512_));
AND2X2 AND2X2_3064 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8513_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8514_));
AND2X2 AND2X2_3065 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8267_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8516_));
AND2X2 AND2X2_3066 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8517_));
AND2X2 AND2X2_3067 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8518_));
AND2X2 AND2X2_3068 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8519_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8520_));
AND2X2 AND2X2_3069 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8521_), .B(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8522_));
AND2X2 AND2X2_307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2816_));
AND2X2 AND2X2_3070 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8525_), .B(AES_CORE_DATAPATH_col_en_host_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8526_));
AND2X2 AND2X2_3071 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n8527_));
AND2X2 AND2X2_3072 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n8528_));
AND2X2 AND2X2_3073 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8528_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8529_));
AND2X2 AND2X2_3074 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8532_));
AND2X2 AND2X2_3075 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5808_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8533_));
AND2X2 AND2X2_3076 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8535_));
AND2X2 AND2X2_3077 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5858_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8536_));
AND2X2 AND2X2_3078 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8538_));
AND2X2 AND2X2_3079 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5908_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8539_));
AND2X2 AND2X2_308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2817_), .B(AES_CORE_DATAPATH__abc_16009_new_n2807_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2818_));
AND2X2 AND2X2_3080 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8541_));
AND2X2 AND2X2_3081 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5958_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8542_));
AND2X2 AND2X2_3082 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8544_));
AND2X2 AND2X2_3083 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6008_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8545_));
AND2X2 AND2X2_3084 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8547_));
AND2X2 AND2X2_3085 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6058_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8548_));
AND2X2 AND2X2_3086 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8550_));
AND2X2 AND2X2_3087 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6108_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8551_));
AND2X2 AND2X2_3088 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8553_));
AND2X2 AND2X2_3089 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6158_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8554_));
AND2X2 AND2X2_309 ( .A(AES_CORE_CONTROL_UNIT_key_out_sel_0_), .B(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n2819_));
AND2X2 AND2X2_3090 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8556_));
AND2X2 AND2X2_3091 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6208_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8557_));
AND2X2 AND2X2_3092 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8559_));
AND2X2 AND2X2_3093 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6258_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8560_));
AND2X2 AND2X2_3094 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8562_));
AND2X2 AND2X2_3095 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6308_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8563_));
AND2X2 AND2X2_3096 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8565_));
AND2X2 AND2X2_3097 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6358_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8566_));
AND2X2 AND2X2_3098 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8568_));
AND2X2 AND2X2_3099 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6408_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8569_));
AND2X2 AND2X2_31 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n112_));
AND2X2 AND2X2_310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2825_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2826_));
AND2X2 AND2X2_3100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8571_));
AND2X2 AND2X2_3101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6458_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8572_));
AND2X2 AND2X2_3102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8574_));
AND2X2 AND2X2_3103 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6508_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8575_));
AND2X2 AND2X2_3104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8577_));
AND2X2 AND2X2_3105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6558_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8578_));
AND2X2 AND2X2_3106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8580_));
AND2X2 AND2X2_3107 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6608_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8581_));
AND2X2 AND2X2_3108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8583_));
AND2X2 AND2X2_3109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6658_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8584_));
AND2X2 AND2X2_311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2814_), .B(AES_CORE_DATAPATH__abc_16009_new_n2821_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2828_));
AND2X2 AND2X2_3110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8586_));
AND2X2 AND2X2_3111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6708_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8587_));
AND2X2 AND2X2_3112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8589_));
AND2X2 AND2X2_3113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6758_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8590_));
AND2X2 AND2X2_3114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8592_));
AND2X2 AND2X2_3115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6808_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8593_));
AND2X2 AND2X2_3116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8595_));
AND2X2 AND2X2_3117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6858_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8596_));
AND2X2 AND2X2_3118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8598_));
AND2X2 AND2X2_3119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6908_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8599_));
AND2X2 AND2X2_312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2829_));
AND2X2 AND2X2_3120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8601_));
AND2X2 AND2X2_3121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6958_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8602_));
AND2X2 AND2X2_3122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8604_));
AND2X2 AND2X2_3123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7008_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8605_));
AND2X2 AND2X2_3124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8607_));
AND2X2 AND2X2_3125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7058_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8608_));
AND2X2 AND2X2_3126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8610_));
AND2X2 AND2X2_3127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7108_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8611_));
AND2X2 AND2X2_3128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8613_));
AND2X2 AND2X2_3129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7158_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8614_));
AND2X2 AND2X2_313 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2833_), .B(AES_CORE_DATAPATH__abc_16009_new_n2831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2834_));
AND2X2 AND2X2_3130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8616_));
AND2X2 AND2X2_3131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7208_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8617_));
AND2X2 AND2X2_3132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8619_));
AND2X2 AND2X2_3133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7258_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8620_));
AND2X2 AND2X2_3134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8622_));
AND2X2 AND2X2_3135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7308_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8623_));
AND2X2 AND2X2_3136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH_bkp_1_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8625_));
AND2X2 AND2X2_3137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7358_), .B(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8626_));
AND2X2 AND2X2_3138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8630_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8631_));
AND2X2 AND2X2_3139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8629_), .B(AES_CORE_DATAPATH__abc_16009_new_n8631_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8632_));
AND2X2 AND2X2_314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2835_), .B(AES_CORE_DATAPATH__abc_16009_new_n2836_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2837_));
AND2X2 AND2X2_3140 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8633_));
AND2X2 AND2X2_3141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8635_), .B(AES_CORE_DATAPATH__abc_16009_new_n8636_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__0_));
AND2X2 AND2X2_3142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8639_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8640_));
AND2X2 AND2X2_3143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8638_), .B(AES_CORE_DATAPATH__abc_16009_new_n8640_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8641_));
AND2X2 AND2X2_3144 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8642_));
AND2X2 AND2X2_3145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8644_), .B(AES_CORE_DATAPATH__abc_16009_new_n8645_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__1_));
AND2X2 AND2X2_3146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8648_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8649_));
AND2X2 AND2X2_3147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8647_), .B(AES_CORE_DATAPATH__abc_16009_new_n8649_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8650_));
AND2X2 AND2X2_3148 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8651_));
AND2X2 AND2X2_3149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8653_), .B(AES_CORE_DATAPATH__abc_16009_new_n8654_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__2_));
AND2X2 AND2X2_315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2837_), .B(AES_CORE_DATAPATH__abc_16009_new_n2821_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2838_));
AND2X2 AND2X2_3150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8657_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8658_));
AND2X2 AND2X2_3151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8656_), .B(AES_CORE_DATAPATH__abc_16009_new_n8658_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8659_));
AND2X2 AND2X2_3152 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8660_));
AND2X2 AND2X2_3153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8662_), .B(AES_CORE_DATAPATH__abc_16009_new_n8663_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__3_));
AND2X2 AND2X2_3154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8666_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8667_));
AND2X2 AND2X2_3155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8665_), .B(AES_CORE_DATAPATH__abc_16009_new_n8667_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8668_));
AND2X2 AND2X2_3156 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8669_));
AND2X2 AND2X2_3157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8671_), .B(AES_CORE_DATAPATH__abc_16009_new_n8672_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__4_));
AND2X2 AND2X2_3158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8675_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8676_));
AND2X2 AND2X2_3159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8674_), .B(AES_CORE_DATAPATH__abc_16009_new_n8676_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8677_));
AND2X2 AND2X2_316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2839_));
AND2X2 AND2X2_3160 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8678_));
AND2X2 AND2X2_3161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8680_), .B(AES_CORE_DATAPATH__abc_16009_new_n8681_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__5_));
AND2X2 AND2X2_3162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8684_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8685_));
AND2X2 AND2X2_3163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8683_), .B(AES_CORE_DATAPATH__abc_16009_new_n8685_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8686_));
AND2X2 AND2X2_3164 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8687_));
AND2X2 AND2X2_3165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8689_), .B(AES_CORE_DATAPATH__abc_16009_new_n8690_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__6_));
AND2X2 AND2X2_3166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8693_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8694_));
AND2X2 AND2X2_3167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8692_), .B(AES_CORE_DATAPATH__abc_16009_new_n8694_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8695_));
AND2X2 AND2X2_3168 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8696_));
AND2X2 AND2X2_3169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8698_), .B(AES_CORE_DATAPATH__abc_16009_new_n8699_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__7_));
AND2X2 AND2X2_317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2841_), .B(AES_CORE_DATAPATH__abc_16009_new_n2823_), .Y(\key_out[0] ));
AND2X2 AND2X2_3170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8702_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8703_));
AND2X2 AND2X2_3171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8701_), .B(AES_CORE_DATAPATH__abc_16009_new_n8703_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8704_));
AND2X2 AND2X2_3172 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8705_));
AND2X2 AND2X2_3173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8707_), .B(AES_CORE_DATAPATH__abc_16009_new_n8708_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__8_));
AND2X2 AND2X2_3174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8711_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8712_));
AND2X2 AND2X2_3175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8710_), .B(AES_CORE_DATAPATH__abc_16009_new_n8712_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8713_));
AND2X2 AND2X2_3176 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8714_));
AND2X2 AND2X2_3177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8716_), .B(AES_CORE_DATAPATH__abc_16009_new_n8717_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__9_));
AND2X2 AND2X2_3178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8720_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8721_));
AND2X2 AND2X2_3179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8719_), .B(AES_CORE_DATAPATH__abc_16009_new_n8721_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8722_));
AND2X2 AND2X2_318 ( .A(\key_out[0] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2806_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2843_));
AND2X2 AND2X2_3180 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8723_));
AND2X2 AND2X2_3181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8725_), .B(AES_CORE_DATAPATH__abc_16009_new_n8726_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__10_));
AND2X2 AND2X2_3182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8729_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8730_));
AND2X2 AND2X2_3183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8728_), .B(AES_CORE_DATAPATH__abc_16009_new_n8730_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8731_));
AND2X2 AND2X2_3184 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8732_));
AND2X2 AND2X2_3185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8734_), .B(AES_CORE_DATAPATH__abc_16009_new_n8735_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__11_));
AND2X2 AND2X2_3186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8738_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8739_));
AND2X2 AND2X2_3187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8737_), .B(AES_CORE_DATAPATH__abc_16009_new_n8739_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8740_));
AND2X2 AND2X2_3188 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8741_));
AND2X2 AND2X2_3189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8743_), .B(AES_CORE_DATAPATH__abc_16009_new_n8744_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__12_));
AND2X2 AND2X2_319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2844_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2845_));
AND2X2 AND2X2_3190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8747_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8748_));
AND2X2 AND2X2_3191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8746_), .B(AES_CORE_DATAPATH__abc_16009_new_n8748_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8749_));
AND2X2 AND2X2_3192 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8750_));
AND2X2 AND2X2_3193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8752_), .B(AES_CORE_DATAPATH__abc_16009_new_n8753_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__13_));
AND2X2 AND2X2_3194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8756_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8757_));
AND2X2 AND2X2_3195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8755_), .B(AES_CORE_DATAPATH__abc_16009_new_n8757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8758_));
AND2X2 AND2X2_3196 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8759_));
AND2X2 AND2X2_3197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8761_), .B(AES_CORE_DATAPATH__abc_16009_new_n8762_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__14_));
AND2X2 AND2X2_3198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8765_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8766_));
AND2X2 AND2X2_3199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8764_), .B(AES_CORE_DATAPATH__abc_16009_new_n8766_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8767_));
AND2X2 AND2X2_32 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n113_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n114_));
AND2X2 AND2X2_320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2847_), .B(AES_CORE_DATAPATH__abc_16009_new_n2804_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__0_));
AND2X2 AND2X2_3200 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8768_));
AND2X2 AND2X2_3201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8770_), .B(AES_CORE_DATAPATH__abc_16009_new_n8771_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__15_));
AND2X2 AND2X2_3202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8774_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8775_));
AND2X2 AND2X2_3203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8773_), .B(AES_CORE_DATAPATH__abc_16009_new_n8775_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8776_));
AND2X2 AND2X2_3204 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8777_));
AND2X2 AND2X2_3205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8779_), .B(AES_CORE_DATAPATH__abc_16009_new_n8780_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__16_));
AND2X2 AND2X2_3206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8783_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8784_));
AND2X2 AND2X2_3207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8782_), .B(AES_CORE_DATAPATH__abc_16009_new_n8784_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8785_));
AND2X2 AND2X2_3208 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8786_));
AND2X2 AND2X2_3209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8788_), .B(AES_CORE_DATAPATH__abc_16009_new_n8789_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__17_));
AND2X2 AND2X2_321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2852_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2853_));
AND2X2 AND2X2_3210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8792_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8793_));
AND2X2 AND2X2_3211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8791_), .B(AES_CORE_DATAPATH__abc_16009_new_n8793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8794_));
AND2X2 AND2X2_3212 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8795_));
AND2X2 AND2X2_3213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8797_), .B(AES_CORE_DATAPATH__abc_16009_new_n8798_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__18_));
AND2X2 AND2X2_3214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8801_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8802_));
AND2X2 AND2X2_3215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8800_), .B(AES_CORE_DATAPATH__abc_16009_new_n8802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8803_));
AND2X2 AND2X2_3216 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8804_));
AND2X2 AND2X2_3217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8806_), .B(AES_CORE_DATAPATH__abc_16009_new_n8807_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__19_));
AND2X2 AND2X2_3218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8810_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8811_));
AND2X2 AND2X2_3219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8809_), .B(AES_CORE_DATAPATH__abc_16009_new_n8811_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8812_));
AND2X2 AND2X2_322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2855_));
AND2X2 AND2X2_3220 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8813_));
AND2X2 AND2X2_3221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8815_), .B(AES_CORE_DATAPATH__abc_16009_new_n8816_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__20_));
AND2X2 AND2X2_3222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8819_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8820_));
AND2X2 AND2X2_3223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8818_), .B(AES_CORE_DATAPATH__abc_16009_new_n8820_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8821_));
AND2X2 AND2X2_3224 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8822_));
AND2X2 AND2X2_3225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8824_), .B(AES_CORE_DATAPATH__abc_16009_new_n8825_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__21_));
AND2X2 AND2X2_3226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8828_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8829_));
AND2X2 AND2X2_3227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8827_), .B(AES_CORE_DATAPATH__abc_16009_new_n8829_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8830_));
AND2X2 AND2X2_3228 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8831_));
AND2X2 AND2X2_3229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8833_), .B(AES_CORE_DATAPATH__abc_16009_new_n8834_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__22_));
AND2X2 AND2X2_323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2856_));
AND2X2 AND2X2_3230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8837_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8838_));
AND2X2 AND2X2_3231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8836_), .B(AES_CORE_DATAPATH__abc_16009_new_n8838_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8839_));
AND2X2 AND2X2_3232 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8840_));
AND2X2 AND2X2_3233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8842_), .B(AES_CORE_DATAPATH__abc_16009_new_n8843_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__23_));
AND2X2 AND2X2_3234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8846_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8847_));
AND2X2 AND2X2_3235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8845_), .B(AES_CORE_DATAPATH__abc_16009_new_n8847_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8848_));
AND2X2 AND2X2_3236 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8849_));
AND2X2 AND2X2_3237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8851_), .B(AES_CORE_DATAPATH__abc_16009_new_n8852_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__24_));
AND2X2 AND2X2_3238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8855_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8856_));
AND2X2 AND2X2_3239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8854_), .B(AES_CORE_DATAPATH__abc_16009_new_n8856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8857_));
AND2X2 AND2X2_324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2858_), .B(AES_CORE_DATAPATH__abc_16009_new_n2859_), .Y(\key_out[1] ));
AND2X2 AND2X2_3240 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8858_));
AND2X2 AND2X2_3241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8860_), .B(AES_CORE_DATAPATH__abc_16009_new_n8861_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__25_));
AND2X2 AND2X2_3242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8864_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8865_));
AND2X2 AND2X2_3243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8863_), .B(AES_CORE_DATAPATH__abc_16009_new_n8865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8866_));
AND2X2 AND2X2_3244 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8867_));
AND2X2 AND2X2_3245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8869_), .B(AES_CORE_DATAPATH__abc_16009_new_n8870_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__26_));
AND2X2 AND2X2_3246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8873_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8874_));
AND2X2 AND2X2_3247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8872_), .B(AES_CORE_DATAPATH__abc_16009_new_n8874_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8875_));
AND2X2 AND2X2_3248 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8876_));
AND2X2 AND2X2_3249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8878_), .B(AES_CORE_DATAPATH__abc_16009_new_n8879_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__27_));
AND2X2 AND2X2_325 ( .A(\key_out[1] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2850_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2861_));
AND2X2 AND2X2_3250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8882_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8883_));
AND2X2 AND2X2_3251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8881_), .B(AES_CORE_DATAPATH__abc_16009_new_n8883_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8884_));
AND2X2 AND2X2_3252 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8885_));
AND2X2 AND2X2_3253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8887_), .B(AES_CORE_DATAPATH__abc_16009_new_n8888_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__28_));
AND2X2 AND2X2_3254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8891_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8892_));
AND2X2 AND2X2_3255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8890_), .B(AES_CORE_DATAPATH__abc_16009_new_n8892_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8893_));
AND2X2 AND2X2_3256 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8894_));
AND2X2 AND2X2_3257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8896_), .B(AES_CORE_DATAPATH__abc_16009_new_n8897_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__29_));
AND2X2 AND2X2_3258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8900_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8901_));
AND2X2 AND2X2_3259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8899_), .B(AES_CORE_DATAPATH__abc_16009_new_n8901_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8902_));
AND2X2 AND2X2_326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2862_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2863_));
AND2X2 AND2X2_3260 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8903_));
AND2X2 AND2X2_3261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8905_), .B(AES_CORE_DATAPATH__abc_16009_new_n8906_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__30_));
AND2X2 AND2X2_3262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8909_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8910_));
AND2X2 AND2X2_3263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8908_), .B(AES_CORE_DATAPATH__abc_16009_new_n8910_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8911_));
AND2X2 AND2X2_3264 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8912_));
AND2X2 AND2X2_3265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8914_), .B(AES_CORE_DATAPATH__abc_16009_new_n8915_), .Y(AES_CORE_DATAPATH__0bkp_3__31_0__31_));
AND2X2 AND2X2_3266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2802_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8919_));
AND2X2 AND2X2_3267 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8924_));
AND2X2 AND2X2_3268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8924_), .B(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8925_));
AND2X2 AND2X2_3269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8926_), .B(AES_CORE_DATAPATH__abc_16009_new_n8923_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8927_));
AND2X2 AND2X2_327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2865_), .B(AES_CORE_DATAPATH__abc_16009_new_n2849_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__1_));
AND2X2 AND2X2_3270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8928_), .B(AES_CORE_DATAPATH__abc_16009_new_n8922_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__0_));
AND2X2 AND2X2_3271 ( .A(AES_CORE_DATAPATH_iv_3__0_), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8931_));
AND2X2 AND2X2_3272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8931_), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_16009_new_n8932_));
AND2X2 AND2X2_3273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8932_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8933_));
AND2X2 AND2X2_3274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8934_), .B(AES_CORE_DATAPATH__abc_16009_new_n8930_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8935_));
AND2X2 AND2X2_3275 ( .A(AES_CORE_DATAPATH_iv_3__0_), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_16009_new_n8938_));
AND2X2 AND2X2_3276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8939_), .B(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8940_));
AND2X2 AND2X2_3277 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8936_), .B(AES_CORE_DATAPATH__abc_16009_new_n8941_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__1_));
AND2X2 AND2X2_3278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8943_), .B(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8944_));
AND2X2 AND2X2_3279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8932_), .B(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8947_));
AND2X2 AND2X2_328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2870_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2871_));
AND2X2 AND2X2_3280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8947_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8948_));
AND2X2 AND2X2_3281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8949_), .B(AES_CORE_DATAPATH__abc_16009_new_n8946_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8950_));
AND2X2 AND2X2_3282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8951_), .B(AES_CORE_DATAPATH__abc_16009_new_n8945_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__2_));
AND2X2 AND2X2_3283 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8953_), .B(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8954_));
AND2X2 AND2X2_3284 ( .A(AES_CORE_DATAPATH_iv_3__2_), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8957_));
AND2X2 AND2X2_3285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8931_), .B(AES_CORE_DATAPATH__abc_16009_new_n8957_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8958_));
AND2X2 AND2X2_3286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8958_), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_16009_new_n8959_));
AND2X2 AND2X2_3287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8959_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8960_));
AND2X2 AND2X2_3288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8961_), .B(AES_CORE_DATAPATH__abc_16009_new_n8956_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8962_));
AND2X2 AND2X2_3289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8963_), .B(AES_CORE_DATAPATH__abc_16009_new_n8955_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__3_));
AND2X2 AND2X2_329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2873_));
AND2X2 AND2X2_3290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8965_), .B(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8966_));
AND2X2 AND2X2_3291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8959_), .B(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8969_));
AND2X2 AND2X2_3292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8969_), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8970_));
AND2X2 AND2X2_3293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8971_), .B(AES_CORE_DATAPATH__abc_16009_new_n8968_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8972_));
AND2X2 AND2X2_3294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8973_), .B(AES_CORE_DATAPATH__abc_16009_new_n8967_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__4_));
AND2X2 AND2X2_3295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8975_));
AND2X2 AND2X2_3296 ( .A(AES_CORE_DATAPATH_iv_3__4_), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8977_));
AND2X2 AND2X2_3297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8959_), .B(AES_CORE_DATAPATH__abc_16009_new_n8977_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8978_));
AND2X2 AND2X2_3298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8976_), .B(AES_CORE_DATAPATH__abc_16009_new_n8979_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8980_));
AND2X2 AND2X2_3299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH__abc_16009_new_n8982_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8983_));
AND2X2 AND2X2_33 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n114_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n102_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n115_));
AND2X2 AND2X2_330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2874_));
AND2X2 AND2X2_3300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8981_), .B(AES_CORE_DATAPATH__abc_16009_new_n8983_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8984_));
AND2X2 AND2X2_3301 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8986_));
AND2X2 AND2X2_3302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH__abc_16009_new_n8987_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8988_));
AND2X2 AND2X2_3303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8979_), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8989_));
AND2X2 AND2X2_3304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8978_), .B(AES_CORE_DATAPATH__abc_16009_new_n8990_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8991_));
AND2X2 AND2X2_3305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8993_), .B(AES_CORE_DATAPATH__abc_16009_new_n8988_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8994_));
AND2X2 AND2X2_3306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n8996_));
AND2X2 AND2X2_3307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8977_), .B(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8997_));
AND2X2 AND2X2_3308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8958_), .B(AES_CORE_DATAPATH__abc_16009_new_n8997_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8998_));
AND2X2 AND2X2_3309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8998_), .B(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8999_));
AND2X2 AND2X2_331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2876_), .B(AES_CORE_DATAPATH__abc_16009_new_n2877_), .Y(\key_out[2] ));
AND2X2 AND2X2_3310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9000_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9001_));
AND2X2 AND2X2_3311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9001_), .B(AES_CORE_DATAPATH__abc_16009_new_n8998_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9002_));
AND2X2 AND2X2_3312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9003_), .B(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9004_));
AND2X2 AND2X2_3313 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9005_), .B(AES_CORE_DATAPATH_iv_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9006_));
AND2X2 AND2X2_3314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9008_));
AND2X2 AND2X2_3315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8999_), .B(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9009_));
AND2X2 AND2X2_3316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9010_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9011_));
AND2X2 AND2X2_3317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9011_), .B(AES_CORE_DATAPATH__abc_16009_new_n8999_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9012_));
AND2X2 AND2X2_3318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9013_), .B(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9014_));
AND2X2 AND2X2_3319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9015_), .B(AES_CORE_DATAPATH_iv_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9016_));
AND2X2 AND2X2_332 ( .A(\key_out[2] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2868_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2879_));
AND2X2 AND2X2_3320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9020_));
AND2X2 AND2X2_3321 ( .A(AES_CORE_DATAPATH_iv_3__8_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9021_));
AND2X2 AND2X2_3322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8999_), .B(AES_CORE_DATAPATH__abc_16009_new_n9021_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9022_));
AND2X2 AND2X2_3323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9023_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9024_));
AND2X2 AND2X2_3324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9025_), .B(AES_CORE_DATAPATH__abc_16009_new_n9019_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9026_));
AND2X2 AND2X2_3325 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9027_));
AND2X2 AND2X2_3326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9029_), .B(AES_CORE_DATAPATH__abc_16009_new_n9018_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__9_));
AND2X2 AND2X2_3327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9022_), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9033_));
AND2X2 AND2X2_3328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9034_), .B(AES_CORE_DATAPATH__abc_16009_new_n9032_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9035_));
AND2X2 AND2X2_3329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9035_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9036_));
AND2X2 AND2X2_333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2880_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2881_));
AND2X2 AND2X2_3330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9037_));
AND2X2 AND2X2_3331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9038_));
AND2X2 AND2X2_3332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9041_), .B(AES_CORE_DATAPATH__abc_16009_new_n9031_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__10_));
AND2X2 AND2X2_3333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9045_));
AND2X2 AND2X2_3334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9033_), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9046_));
AND2X2 AND2X2_3335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9047_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9048_));
AND2X2 AND2X2_3336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9049_), .B(AES_CORE_DATAPATH__abc_16009_new_n9044_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9050_));
AND2X2 AND2X2_3337 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9051_));
AND2X2 AND2X2_3338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9053_), .B(AES_CORE_DATAPATH__abc_16009_new_n9043_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__11_));
AND2X2 AND2X2_3339 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9046_), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9056_));
AND2X2 AND2X2_334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2883_), .B(AES_CORE_DATAPATH__abc_16009_new_n2867_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__2_));
AND2X2 AND2X2_3340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9058_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9059_));
AND2X2 AND2X2_3341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9059_), .B(AES_CORE_DATAPATH__abc_16009_new_n9057_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9060_));
AND2X2 AND2X2_3342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9061_));
AND2X2 AND2X2_3343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9062_));
AND2X2 AND2X2_3344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9065_), .B(AES_CORE_DATAPATH__abc_16009_new_n9055_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__12_));
AND2X2 AND2X2_3345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9056_), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9068_));
AND2X2 AND2X2_3346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9070_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9071_));
AND2X2 AND2X2_3347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9071_), .B(AES_CORE_DATAPATH__abc_16009_new_n9069_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9072_));
AND2X2 AND2X2_3348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9073_));
AND2X2 AND2X2_3349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9074_));
AND2X2 AND2X2_335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2889_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2890_));
AND2X2 AND2X2_3350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9077_), .B(AES_CORE_DATAPATH__abc_16009_new_n9067_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__13_));
AND2X2 AND2X2_3351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9068_), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9080_));
AND2X2 AND2X2_3352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9082_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9083_));
AND2X2 AND2X2_3353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9083_), .B(AES_CORE_DATAPATH__abc_16009_new_n9081_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9084_));
AND2X2 AND2X2_3354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9085_));
AND2X2 AND2X2_3355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9086_));
AND2X2 AND2X2_3356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9089_), .B(AES_CORE_DATAPATH__abc_16009_new_n9079_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__14_));
AND2X2 AND2X2_3357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9080_), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9092_));
AND2X2 AND2X2_3358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9094_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9095_));
AND2X2 AND2X2_3359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9095_), .B(AES_CORE_DATAPATH__abc_16009_new_n9093_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9096_));
AND2X2 AND2X2_336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2892_));
AND2X2 AND2X2_3360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9097_));
AND2X2 AND2X2_3361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9098_));
AND2X2 AND2X2_3362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9101_), .B(AES_CORE_DATAPATH__abc_16009_new_n9091_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__15_));
AND2X2 AND2X2_3363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9092_), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9104_));
AND2X2 AND2X2_3364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9106_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9107_));
AND2X2 AND2X2_3365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9107_), .B(AES_CORE_DATAPATH__abc_16009_new_n9105_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9108_));
AND2X2 AND2X2_3366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9109_));
AND2X2 AND2X2_3367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9110_));
AND2X2 AND2X2_3368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9113_), .B(AES_CORE_DATAPATH__abc_16009_new_n9103_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__16_));
AND2X2 AND2X2_3369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9104_), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9116_));
AND2X2 AND2X2_337 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2893_));
AND2X2 AND2X2_3370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9118_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9119_));
AND2X2 AND2X2_3371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9119_), .B(AES_CORE_DATAPATH__abc_16009_new_n9117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9120_));
AND2X2 AND2X2_3372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9121_));
AND2X2 AND2X2_3373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9122_));
AND2X2 AND2X2_3374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9125_), .B(AES_CORE_DATAPATH__abc_16009_new_n9115_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__17_));
AND2X2 AND2X2_3375 ( .A(AES_CORE_DATAPATH_iv_3__17_), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9129_));
AND2X2 AND2X2_3376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9104_), .B(AES_CORE_DATAPATH__abc_16009_new_n9129_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9130_));
AND2X2 AND2X2_3377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9131_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9132_));
AND2X2 AND2X2_3378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9132_), .B(AES_CORE_DATAPATH__abc_16009_new_n9128_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9133_));
AND2X2 AND2X2_3379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9134_));
AND2X2 AND2X2_338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2895_), .B(AES_CORE_DATAPATH__abc_16009_new_n2887_), .Y(\key_out[3] ));
AND2X2 AND2X2_3380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9135_));
AND2X2 AND2X2_3381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9138_), .B(AES_CORE_DATAPATH__abc_16009_new_n9127_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__18_));
AND2X2 AND2X2_3382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9130_), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9141_));
AND2X2 AND2X2_3383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9143_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9144_));
AND2X2 AND2X2_3384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9144_), .B(AES_CORE_DATAPATH__abc_16009_new_n9142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9145_));
AND2X2 AND2X2_3385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9146_));
AND2X2 AND2X2_3386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9147_));
AND2X2 AND2X2_3387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9150_), .B(AES_CORE_DATAPATH__abc_16009_new_n9140_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__19_));
AND2X2 AND2X2_3388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9129_), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9153_));
AND2X2 AND2X2_3389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9104_), .B(AES_CORE_DATAPATH__abc_16009_new_n9153_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9154_));
AND2X2 AND2X2_339 ( .A(\key_out[3] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2897_));
AND2X2 AND2X2_3390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9154_), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9156_));
AND2X2 AND2X2_3391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9157_), .B(AES_CORE_DATAPATH__abc_16009_new_n9155_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9158_));
AND2X2 AND2X2_3392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9158_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9159_));
AND2X2 AND2X2_3393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9160_));
AND2X2 AND2X2_3394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9161_));
AND2X2 AND2X2_3395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9164_), .B(AES_CORE_DATAPATH__abc_16009_new_n9152_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__20_));
AND2X2 AND2X2_3396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9157_), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9167_));
AND2X2 AND2X2_3397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9156_), .B(AES_CORE_DATAPATH__abc_16009_new_n9168_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9169_));
AND2X2 AND2X2_3398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9170_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9171_));
AND2X2 AND2X2_3399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9172_));
AND2X2 AND2X2_34 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n118_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n119_));
AND2X2 AND2X2_340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2898_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2899_));
AND2X2 AND2X2_3400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9173_));
AND2X2 AND2X2_3401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9176_), .B(AES_CORE_DATAPATH__abc_16009_new_n9166_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__21_));
AND2X2 AND2X2_3402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9156_), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9179_));
AND2X2 AND2X2_3403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9141_), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9181_));
AND2X2 AND2X2_3404 ( .A(AES_CORE_DATAPATH_iv_3__21_), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9182_));
AND2X2 AND2X2_3405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9181_), .B(AES_CORE_DATAPATH__abc_16009_new_n9182_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9183_));
AND2X2 AND2X2_3406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9184_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9185_));
AND2X2 AND2X2_3407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9185_), .B(AES_CORE_DATAPATH__abc_16009_new_n9180_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9186_));
AND2X2 AND2X2_3408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9187_));
AND2X2 AND2X2_3409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9188_));
AND2X2 AND2X2_341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2901_), .B(AES_CORE_DATAPATH__abc_16009_new_n2885_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__3_));
AND2X2 AND2X2_3410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9191_), .B(AES_CORE_DATAPATH__abc_16009_new_n9178_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__22_));
AND2X2 AND2X2_3411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9183_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9194_));
AND2X2 AND2X2_3412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9196_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9197_));
AND2X2 AND2X2_3413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9197_), .B(AES_CORE_DATAPATH__abc_16009_new_n9195_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9198_));
AND2X2 AND2X2_3414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9199_));
AND2X2 AND2X2_3415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9200_));
AND2X2 AND2X2_3416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9203_), .B(AES_CORE_DATAPATH__abc_16009_new_n9193_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__23_));
AND2X2 AND2X2_3417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9182_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9206_));
AND2X2 AND2X2_3418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9156_), .B(AES_CORE_DATAPATH__abc_16009_new_n9206_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9207_));
AND2X2 AND2X2_3419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9207_), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9209_));
AND2X2 AND2X2_342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2907_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2908_));
AND2X2 AND2X2_3420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9210_), .B(AES_CORE_DATAPATH__abc_16009_new_n9208_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9211_));
AND2X2 AND2X2_3421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9211_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9212_));
AND2X2 AND2X2_3422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9213_));
AND2X2 AND2X2_3423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9214_));
AND2X2 AND2X2_3424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9217_), .B(AES_CORE_DATAPATH__abc_16009_new_n9205_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__24_));
AND2X2 AND2X2_3425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9210_), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9220_));
AND2X2 AND2X2_3426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9209_), .B(AES_CORE_DATAPATH__abc_16009_new_n9221_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9222_));
AND2X2 AND2X2_3427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9223_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9224_));
AND2X2 AND2X2_3428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9225_));
AND2X2 AND2X2_3429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9226_));
AND2X2 AND2X2_343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2910_));
AND2X2 AND2X2_3430 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9229_), .B(AES_CORE_DATAPATH__abc_16009_new_n9219_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__25_));
AND2X2 AND2X2_3431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9209_), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9232_));
AND2X2 AND2X2_3432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9232_), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9234_));
AND2X2 AND2X2_3433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9235_), .B(AES_CORE_DATAPATH__abc_16009_new_n9233_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9236_));
AND2X2 AND2X2_3434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9236_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9237_));
AND2X2 AND2X2_3435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9238_));
AND2X2 AND2X2_3436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9239_));
AND2X2 AND2X2_3437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9242_), .B(AES_CORE_DATAPATH__abc_16009_new_n9231_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__26_));
AND2X2 AND2X2_3438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9234_), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9246_));
AND2X2 AND2X2_3439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9247_), .B(AES_CORE_DATAPATH__abc_16009_new_n9245_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9248_));
AND2X2 AND2X2_344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2911_));
AND2X2 AND2X2_3440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9248_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9249_));
AND2X2 AND2X2_3441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9250_));
AND2X2 AND2X2_3442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9251_));
AND2X2 AND2X2_3443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9254_), .B(AES_CORE_DATAPATH__abc_16009_new_n9244_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__27_));
AND2X2 AND2X2_3444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9246_), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9258_));
AND2X2 AND2X2_3445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9259_), .B(AES_CORE_DATAPATH__abc_16009_new_n9257_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9260_));
AND2X2 AND2X2_3446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9260_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9261_));
AND2X2 AND2X2_3447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9262_));
AND2X2 AND2X2_3448 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9263_));
AND2X2 AND2X2_3449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9266_), .B(AES_CORE_DATAPATH__abc_16009_new_n9256_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__28_));
AND2X2 AND2X2_345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2913_), .B(AES_CORE_DATAPATH__abc_16009_new_n2905_), .Y(\key_out[4] ));
AND2X2 AND2X2_3450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9258_), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9270_));
AND2X2 AND2X2_3451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9271_), .B(AES_CORE_DATAPATH__abc_16009_new_n9269_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9272_));
AND2X2 AND2X2_3452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9272_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9273_));
AND2X2 AND2X2_3453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9274_));
AND2X2 AND2X2_3454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9275_));
AND2X2 AND2X2_3455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9278_), .B(AES_CORE_DATAPATH__abc_16009_new_n9268_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__29_));
AND2X2 AND2X2_3456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9270_), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9281_));
AND2X2 AND2X2_3457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9283_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9284_));
AND2X2 AND2X2_3458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9284_), .B(AES_CORE_DATAPATH__abc_16009_new_n9282_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9285_));
AND2X2 AND2X2_3459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9286_));
AND2X2 AND2X2_346 ( .A(\key_out[4] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2904_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2915_));
AND2X2 AND2X2_3460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9287_));
AND2X2 AND2X2_3461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9290_), .B(AES_CORE_DATAPATH__abc_16009_new_n9280_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__30_));
AND2X2 AND2X2_3462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9282_), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9293_));
AND2X2 AND2X2_3463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9281_), .B(AES_CORE_DATAPATH__abc_16009_new_n9294_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9295_));
AND2X2 AND2X2_3464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9296_), .B(AES_CORE_DATAPATH__abc_16009_new_n8924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9297_));
AND2X2 AND2X2_3465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8919_), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9298_));
AND2X2 AND2X2_3466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8937_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9299_));
AND2X2 AND2X2_3467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9302_), .B(AES_CORE_DATAPATH__abc_16009_new_n9292_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__31_));
AND2X2 AND2X2_3468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9306_), .B(AES_CORE_DATAPATH__abc_16009_new_n9304_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__0_));
AND2X2 AND2X2_3469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9309_), .B(AES_CORE_DATAPATH__abc_16009_new_n9308_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__1_));
AND2X2 AND2X2_347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2916_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2917_));
AND2X2 AND2X2_3470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9312_), .B(AES_CORE_DATAPATH__abc_16009_new_n9311_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__2_));
AND2X2 AND2X2_3471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9315_), .B(AES_CORE_DATAPATH__abc_16009_new_n9314_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__3_));
AND2X2 AND2X2_3472 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9318_), .B(AES_CORE_DATAPATH__abc_16009_new_n9317_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__4_));
AND2X2 AND2X2_3473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9321_), .B(AES_CORE_DATAPATH__abc_16009_new_n9320_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__5_));
AND2X2 AND2X2_3474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9324_), .B(AES_CORE_DATAPATH__abc_16009_new_n9323_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__6_));
AND2X2 AND2X2_3475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9327_), .B(AES_CORE_DATAPATH__abc_16009_new_n9326_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__7_));
AND2X2 AND2X2_3476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9330_), .B(AES_CORE_DATAPATH__abc_16009_new_n9329_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__8_));
AND2X2 AND2X2_3477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9333_), .B(AES_CORE_DATAPATH__abc_16009_new_n9332_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__9_));
AND2X2 AND2X2_3478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9336_), .B(AES_CORE_DATAPATH__abc_16009_new_n9335_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__10_));
AND2X2 AND2X2_3479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9339_), .B(AES_CORE_DATAPATH__abc_16009_new_n9338_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__11_));
AND2X2 AND2X2_348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2919_), .B(AES_CORE_DATAPATH__abc_16009_new_n2903_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__4_));
AND2X2 AND2X2_3480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9342_), .B(AES_CORE_DATAPATH__abc_16009_new_n9341_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__12_));
AND2X2 AND2X2_3481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9345_), .B(AES_CORE_DATAPATH__abc_16009_new_n9344_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__13_));
AND2X2 AND2X2_3482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9348_), .B(AES_CORE_DATAPATH__abc_16009_new_n9347_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__14_));
AND2X2 AND2X2_3483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9351_), .B(AES_CORE_DATAPATH__abc_16009_new_n9350_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__15_));
AND2X2 AND2X2_3484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9354_), .B(AES_CORE_DATAPATH__abc_16009_new_n9353_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__16_));
AND2X2 AND2X2_3485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9357_), .B(AES_CORE_DATAPATH__abc_16009_new_n9356_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__17_));
AND2X2 AND2X2_3486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9360_), .B(AES_CORE_DATAPATH__abc_16009_new_n9359_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__18_));
AND2X2 AND2X2_3487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9363_), .B(AES_CORE_DATAPATH__abc_16009_new_n9362_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__19_));
AND2X2 AND2X2_3488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9366_), .B(AES_CORE_DATAPATH__abc_16009_new_n9365_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__20_));
AND2X2 AND2X2_3489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9369_), .B(AES_CORE_DATAPATH__abc_16009_new_n9368_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__21_));
AND2X2 AND2X2_349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2925_));
AND2X2 AND2X2_3490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9372_), .B(AES_CORE_DATAPATH__abc_16009_new_n9371_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__22_));
AND2X2 AND2X2_3491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9375_), .B(AES_CORE_DATAPATH__abc_16009_new_n9374_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__23_));
AND2X2 AND2X2_3492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9378_), .B(AES_CORE_DATAPATH__abc_16009_new_n9377_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__24_));
AND2X2 AND2X2_3493 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9381_), .B(AES_CORE_DATAPATH__abc_16009_new_n9380_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__25_));
AND2X2 AND2X2_3494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9384_), .B(AES_CORE_DATAPATH__abc_16009_new_n9383_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__26_));
AND2X2 AND2X2_3495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9387_), .B(AES_CORE_DATAPATH__abc_16009_new_n9386_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__27_));
AND2X2 AND2X2_3496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9390_), .B(AES_CORE_DATAPATH__abc_16009_new_n9389_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__28_));
AND2X2 AND2X2_3497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9393_), .B(AES_CORE_DATAPATH__abc_16009_new_n9392_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__29_));
AND2X2 AND2X2_3498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9396_), .B(AES_CORE_DATAPATH__abc_16009_new_n9395_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__30_));
AND2X2 AND2X2_3499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9399_), .B(AES_CORE_DATAPATH__abc_16009_new_n9398_), .Y(AES_CORE_DATAPATH__0iv_2__31_0__31_));
AND2X2 AND2X2_35 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n119_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n117_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_1_));
AND2X2 AND2X2_350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2927_));
AND2X2 AND2X2_3500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8525_), .B(AES_CORE_DATAPATH_col_en_host_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9401_));
AND2X2 AND2X2_3501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8528_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9402_));
AND2X2 AND2X2_3502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9405_));
AND2X2 AND2X2_3503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8016_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9406_));
AND2X2 AND2X2_3504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9408_));
AND2X2 AND2X2_3505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8024_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9409_));
AND2X2 AND2X2_3506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9411_));
AND2X2 AND2X2_3507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8032_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9412_));
AND2X2 AND2X2_3508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9414_));
AND2X2 AND2X2_3509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8040_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9415_));
AND2X2 AND2X2_351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2928_));
AND2X2 AND2X2_3510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9417_));
AND2X2 AND2X2_3511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8048_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9418_));
AND2X2 AND2X2_3512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9420_));
AND2X2 AND2X2_3513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8056_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9421_));
AND2X2 AND2X2_3514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9423_));
AND2X2 AND2X2_3515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8064_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9424_));
AND2X2 AND2X2_3516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9426_));
AND2X2 AND2X2_3517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8072_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9427_));
AND2X2 AND2X2_3518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9429_));
AND2X2 AND2X2_3519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8080_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9430_));
AND2X2 AND2X2_352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2930_), .B(AES_CORE_DATAPATH__abc_16009_new_n2931_), .Y(\key_out[5] ));
AND2X2 AND2X2_3520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9432_));
AND2X2 AND2X2_3521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8088_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9433_));
AND2X2 AND2X2_3522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9435_));
AND2X2 AND2X2_3523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8096_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9436_));
AND2X2 AND2X2_3524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9438_));
AND2X2 AND2X2_3525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8104_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9439_));
AND2X2 AND2X2_3526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9441_));
AND2X2 AND2X2_3527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8112_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9442_));
AND2X2 AND2X2_3528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9444_));
AND2X2 AND2X2_3529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8120_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9445_));
AND2X2 AND2X2_353 ( .A(\key_out[5] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2933_));
AND2X2 AND2X2_3530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9447_));
AND2X2 AND2X2_3531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8128_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9448_));
AND2X2 AND2X2_3532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9450_));
AND2X2 AND2X2_3533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8136_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9451_));
AND2X2 AND2X2_3534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9453_));
AND2X2 AND2X2_3535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8144_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9454_));
AND2X2 AND2X2_3536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9456_));
AND2X2 AND2X2_3537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8152_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9457_));
AND2X2 AND2X2_3538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9459_));
AND2X2 AND2X2_3539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8160_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9460_));
AND2X2 AND2X2_354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2934_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2935_));
AND2X2 AND2X2_3540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9462_));
AND2X2 AND2X2_3541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8168_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9463_));
AND2X2 AND2X2_3542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9465_));
AND2X2 AND2X2_3543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8176_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9466_));
AND2X2 AND2X2_3544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9468_));
AND2X2 AND2X2_3545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8184_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9469_));
AND2X2 AND2X2_3546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9471_));
AND2X2 AND2X2_3547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8192_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9472_));
AND2X2 AND2X2_3548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9474_));
AND2X2 AND2X2_3549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8200_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9475_));
AND2X2 AND2X2_355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2937_), .B(AES_CORE_DATAPATH__abc_16009_new_n2921_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__5_));
AND2X2 AND2X2_3550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9477_));
AND2X2 AND2X2_3551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8208_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9478_));
AND2X2 AND2X2_3552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9480_));
AND2X2 AND2X2_3553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8216_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9481_));
AND2X2 AND2X2_3554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9483_));
AND2X2 AND2X2_3555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8224_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9484_));
AND2X2 AND2X2_3556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9486_));
AND2X2 AND2X2_3557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8232_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9487_));
AND2X2 AND2X2_3558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9489_));
AND2X2 AND2X2_3559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8240_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9490_));
AND2X2 AND2X2_356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2943_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2944_));
AND2X2 AND2X2_3560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9492_));
AND2X2 AND2X2_3561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8248_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9493_));
AND2X2 AND2X2_3562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9495_));
AND2X2 AND2X2_3563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8256_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9496_));
AND2X2 AND2X2_3564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH_bkp_1_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9498_));
AND2X2 AND2X2_3565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8264_), .B(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9499_));
AND2X2 AND2X2_3566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9502_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9503_));
AND2X2 AND2X2_3567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9501_), .B(AES_CORE_DATAPATH__abc_16009_new_n9503_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9504_));
AND2X2 AND2X2_3568 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9506_), .B(AES_CORE_DATAPATH__abc_16009_new_n9507_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__0_));
AND2X2 AND2X2_3569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9510_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9511_));
AND2X2 AND2X2_357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2946_));
AND2X2 AND2X2_3570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9509_), .B(AES_CORE_DATAPATH__abc_16009_new_n9511_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9512_));
AND2X2 AND2X2_3571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9514_), .B(AES_CORE_DATAPATH__abc_16009_new_n9515_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__1_));
AND2X2 AND2X2_3572 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9518_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9519_));
AND2X2 AND2X2_3573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9517_), .B(AES_CORE_DATAPATH__abc_16009_new_n9519_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9520_));
AND2X2 AND2X2_3574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9522_), .B(AES_CORE_DATAPATH__abc_16009_new_n9523_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__2_));
AND2X2 AND2X2_3575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9526_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9527_));
AND2X2 AND2X2_3576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9525_), .B(AES_CORE_DATAPATH__abc_16009_new_n9527_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9528_));
AND2X2 AND2X2_3577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9530_), .B(AES_CORE_DATAPATH__abc_16009_new_n9531_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__3_));
AND2X2 AND2X2_3578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9534_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9535_));
AND2X2 AND2X2_3579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9533_), .B(AES_CORE_DATAPATH__abc_16009_new_n9535_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9536_));
AND2X2 AND2X2_358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2947_));
AND2X2 AND2X2_3580 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9538_), .B(AES_CORE_DATAPATH__abc_16009_new_n9539_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__4_));
AND2X2 AND2X2_3581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9542_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9543_));
AND2X2 AND2X2_3582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9541_), .B(AES_CORE_DATAPATH__abc_16009_new_n9543_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9544_));
AND2X2 AND2X2_3583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9546_), .B(AES_CORE_DATAPATH__abc_16009_new_n9547_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__5_));
AND2X2 AND2X2_3584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9550_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9551_));
AND2X2 AND2X2_3585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9549_), .B(AES_CORE_DATAPATH__abc_16009_new_n9551_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9552_));
AND2X2 AND2X2_3586 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9554_), .B(AES_CORE_DATAPATH__abc_16009_new_n9555_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__6_));
AND2X2 AND2X2_3587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9558_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9559_));
AND2X2 AND2X2_3588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9557_), .B(AES_CORE_DATAPATH__abc_16009_new_n9559_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9560_));
AND2X2 AND2X2_3589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9562_), .B(AES_CORE_DATAPATH__abc_16009_new_n9563_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__7_));
AND2X2 AND2X2_359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2949_), .B(AES_CORE_DATAPATH__abc_16009_new_n2941_), .Y(\key_out[6] ));
AND2X2 AND2X2_3590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9566_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9567_));
AND2X2 AND2X2_3591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9565_), .B(AES_CORE_DATAPATH__abc_16009_new_n9567_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9568_));
AND2X2 AND2X2_3592 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9570_), .B(AES_CORE_DATAPATH__abc_16009_new_n9571_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__8_));
AND2X2 AND2X2_3593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9574_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9575_));
AND2X2 AND2X2_3594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9573_), .B(AES_CORE_DATAPATH__abc_16009_new_n9575_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9576_));
AND2X2 AND2X2_3595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9578_), .B(AES_CORE_DATAPATH__abc_16009_new_n9579_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__9_));
AND2X2 AND2X2_3596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9582_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9583_));
AND2X2 AND2X2_3597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9581_), .B(AES_CORE_DATAPATH__abc_16009_new_n9583_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9584_));
AND2X2 AND2X2_3598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9586_), .B(AES_CORE_DATAPATH__abc_16009_new_n9587_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__10_));
AND2X2 AND2X2_3599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9590_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9591_));
AND2X2 AND2X2_36 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_), .B(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n122_));
AND2X2 AND2X2_360 ( .A(\key_out[6] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2940_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2951_));
AND2X2 AND2X2_3600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9589_), .B(AES_CORE_DATAPATH__abc_16009_new_n9591_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9592_));
AND2X2 AND2X2_3601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9594_), .B(AES_CORE_DATAPATH__abc_16009_new_n9595_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__11_));
AND2X2 AND2X2_3602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9598_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9599_));
AND2X2 AND2X2_3603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9597_), .B(AES_CORE_DATAPATH__abc_16009_new_n9599_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9600_));
AND2X2 AND2X2_3604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9602_), .B(AES_CORE_DATAPATH__abc_16009_new_n9603_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__12_));
AND2X2 AND2X2_3605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9606_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9607_));
AND2X2 AND2X2_3606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9605_), .B(AES_CORE_DATAPATH__abc_16009_new_n9607_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9608_));
AND2X2 AND2X2_3607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9610_), .B(AES_CORE_DATAPATH__abc_16009_new_n9611_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__13_));
AND2X2 AND2X2_3608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9614_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9615_));
AND2X2 AND2X2_3609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9613_), .B(AES_CORE_DATAPATH__abc_16009_new_n9615_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9616_));
AND2X2 AND2X2_361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2952_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2953_));
AND2X2 AND2X2_3610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9618_), .B(AES_CORE_DATAPATH__abc_16009_new_n9619_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__14_));
AND2X2 AND2X2_3611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9622_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9623_));
AND2X2 AND2X2_3612 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9621_), .B(AES_CORE_DATAPATH__abc_16009_new_n9623_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9624_));
AND2X2 AND2X2_3613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9626_), .B(AES_CORE_DATAPATH__abc_16009_new_n9627_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__15_));
AND2X2 AND2X2_3614 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9630_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9631_));
AND2X2 AND2X2_3615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9629_), .B(AES_CORE_DATAPATH__abc_16009_new_n9631_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9632_));
AND2X2 AND2X2_3616 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9634_), .B(AES_CORE_DATAPATH__abc_16009_new_n9635_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__16_));
AND2X2 AND2X2_3617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9638_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9639_));
AND2X2 AND2X2_3618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9637_), .B(AES_CORE_DATAPATH__abc_16009_new_n9639_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9640_));
AND2X2 AND2X2_3619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9642_), .B(AES_CORE_DATAPATH__abc_16009_new_n9643_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__17_));
AND2X2 AND2X2_362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2955_), .B(AES_CORE_DATAPATH__abc_16009_new_n2939_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__6_));
AND2X2 AND2X2_3620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9646_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9647_));
AND2X2 AND2X2_3621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9645_), .B(AES_CORE_DATAPATH__abc_16009_new_n9647_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9648_));
AND2X2 AND2X2_3622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9650_), .B(AES_CORE_DATAPATH__abc_16009_new_n9651_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__18_));
AND2X2 AND2X2_3623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9654_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9655_));
AND2X2 AND2X2_3624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9653_), .B(AES_CORE_DATAPATH__abc_16009_new_n9655_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9656_));
AND2X2 AND2X2_3625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9658_), .B(AES_CORE_DATAPATH__abc_16009_new_n9659_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__19_));
AND2X2 AND2X2_3626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9662_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9663_));
AND2X2 AND2X2_3627 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9661_), .B(AES_CORE_DATAPATH__abc_16009_new_n9663_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9664_));
AND2X2 AND2X2_3628 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9666_), .B(AES_CORE_DATAPATH__abc_16009_new_n9667_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__20_));
AND2X2 AND2X2_3629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9670_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9671_));
AND2X2 AND2X2_363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2960_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2961_));
AND2X2 AND2X2_3630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9669_), .B(AES_CORE_DATAPATH__abc_16009_new_n9671_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9672_));
AND2X2 AND2X2_3631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9674_), .B(AES_CORE_DATAPATH__abc_16009_new_n9675_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__21_));
AND2X2 AND2X2_3632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9678_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9679_));
AND2X2 AND2X2_3633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9677_), .B(AES_CORE_DATAPATH__abc_16009_new_n9679_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9680_));
AND2X2 AND2X2_3634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9682_), .B(AES_CORE_DATAPATH__abc_16009_new_n9683_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__22_));
AND2X2 AND2X2_3635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9686_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9687_));
AND2X2 AND2X2_3636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9685_), .B(AES_CORE_DATAPATH__abc_16009_new_n9687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9688_));
AND2X2 AND2X2_3637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9690_), .B(AES_CORE_DATAPATH__abc_16009_new_n9691_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__23_));
AND2X2 AND2X2_3638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9694_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9695_));
AND2X2 AND2X2_3639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9693_), .B(AES_CORE_DATAPATH__abc_16009_new_n9695_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9696_));
AND2X2 AND2X2_364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2963_));
AND2X2 AND2X2_3640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9698_), .B(AES_CORE_DATAPATH__abc_16009_new_n9699_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__24_));
AND2X2 AND2X2_3641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9702_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9703_));
AND2X2 AND2X2_3642 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9701_), .B(AES_CORE_DATAPATH__abc_16009_new_n9703_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9704_));
AND2X2 AND2X2_3643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9706_), .B(AES_CORE_DATAPATH__abc_16009_new_n9707_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__25_));
AND2X2 AND2X2_3644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9710_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9711_));
AND2X2 AND2X2_3645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9709_), .B(AES_CORE_DATAPATH__abc_16009_new_n9711_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9712_));
AND2X2 AND2X2_3646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9714_), .B(AES_CORE_DATAPATH__abc_16009_new_n9715_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__26_));
AND2X2 AND2X2_3647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9718_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9719_));
AND2X2 AND2X2_3648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9717_), .B(AES_CORE_DATAPATH__abc_16009_new_n9719_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9720_));
AND2X2 AND2X2_3649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9722_), .B(AES_CORE_DATAPATH__abc_16009_new_n9723_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__27_));
AND2X2 AND2X2_365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2964_));
AND2X2 AND2X2_3650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9726_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9727_));
AND2X2 AND2X2_3651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9725_), .B(AES_CORE_DATAPATH__abc_16009_new_n9727_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9728_));
AND2X2 AND2X2_3652 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9730_), .B(AES_CORE_DATAPATH__abc_16009_new_n9731_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__28_));
AND2X2 AND2X2_3653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9734_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9735_));
AND2X2 AND2X2_3654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9733_), .B(AES_CORE_DATAPATH__abc_16009_new_n9735_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9736_));
AND2X2 AND2X2_3655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9738_), .B(AES_CORE_DATAPATH__abc_16009_new_n9739_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__29_));
AND2X2 AND2X2_3656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9742_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9743_));
AND2X2 AND2X2_3657 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9741_), .B(AES_CORE_DATAPATH__abc_16009_new_n9743_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9744_));
AND2X2 AND2X2_3658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9746_), .B(AES_CORE_DATAPATH__abc_16009_new_n9747_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__30_));
AND2X2 AND2X2_3659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9750_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9751_));
AND2X2 AND2X2_366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2966_), .B(AES_CORE_DATAPATH__abc_16009_new_n2967_), .Y(\key_out[7] ));
AND2X2 AND2X2_3660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9749_), .B(AES_CORE_DATAPATH__abc_16009_new_n9751_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9752_));
AND2X2 AND2X2_3661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9754_), .B(AES_CORE_DATAPATH__abc_16009_new_n9755_), .Y(AES_CORE_DATAPATH__0bkp_2__31_0__31_));
AND2X2 AND2X2_3662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9759_), .B(AES_CORE_DATAPATH__abc_16009_new_n9757_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__0_));
AND2X2 AND2X2_3663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9762_), .B(AES_CORE_DATAPATH__abc_16009_new_n9761_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__1_));
AND2X2 AND2X2_3664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9765_), .B(AES_CORE_DATAPATH__abc_16009_new_n9764_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__2_));
AND2X2 AND2X2_3665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9768_), .B(AES_CORE_DATAPATH__abc_16009_new_n9767_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__3_));
AND2X2 AND2X2_3666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9771_), .B(AES_CORE_DATAPATH__abc_16009_new_n9770_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__4_));
AND2X2 AND2X2_3667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9774_), .B(AES_CORE_DATAPATH__abc_16009_new_n9773_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__5_));
AND2X2 AND2X2_3668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9777_), .B(AES_CORE_DATAPATH__abc_16009_new_n9776_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__6_));
AND2X2 AND2X2_3669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9780_), .B(AES_CORE_DATAPATH__abc_16009_new_n9779_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__7_));
AND2X2 AND2X2_367 ( .A(\key_out[7] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2958_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2969_));
AND2X2 AND2X2_3670 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9783_), .B(AES_CORE_DATAPATH__abc_16009_new_n9782_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__8_));
AND2X2 AND2X2_3671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9786_), .B(AES_CORE_DATAPATH__abc_16009_new_n9785_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__9_));
AND2X2 AND2X2_3672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9789_), .B(AES_CORE_DATAPATH__abc_16009_new_n9788_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__10_));
AND2X2 AND2X2_3673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9792_), .B(AES_CORE_DATAPATH__abc_16009_new_n9791_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__11_));
AND2X2 AND2X2_3674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9795_), .B(AES_CORE_DATAPATH__abc_16009_new_n9794_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__12_));
AND2X2 AND2X2_3675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9798_), .B(AES_CORE_DATAPATH__abc_16009_new_n9797_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__13_));
AND2X2 AND2X2_3676 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9801_), .B(AES_CORE_DATAPATH__abc_16009_new_n9800_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__14_));
AND2X2 AND2X2_3677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9804_), .B(AES_CORE_DATAPATH__abc_16009_new_n9803_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__15_));
AND2X2 AND2X2_3678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9807_), .B(AES_CORE_DATAPATH__abc_16009_new_n9806_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__16_));
AND2X2 AND2X2_3679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9810_), .B(AES_CORE_DATAPATH__abc_16009_new_n9809_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__17_));
AND2X2 AND2X2_368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2970_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2971_));
AND2X2 AND2X2_3680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9813_), .B(AES_CORE_DATAPATH__abc_16009_new_n9812_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__18_));
AND2X2 AND2X2_3681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9816_), .B(AES_CORE_DATAPATH__abc_16009_new_n9815_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__19_));
AND2X2 AND2X2_3682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9819_), .B(AES_CORE_DATAPATH__abc_16009_new_n9818_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__20_));
AND2X2 AND2X2_3683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9822_), .B(AES_CORE_DATAPATH__abc_16009_new_n9821_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__21_));
AND2X2 AND2X2_3684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9825_), .B(AES_CORE_DATAPATH__abc_16009_new_n9824_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__22_));
AND2X2 AND2X2_3685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9828_), .B(AES_CORE_DATAPATH__abc_16009_new_n9827_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__23_));
AND2X2 AND2X2_3686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9831_), .B(AES_CORE_DATAPATH__abc_16009_new_n9830_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__24_));
AND2X2 AND2X2_3687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9834_), .B(AES_CORE_DATAPATH__abc_16009_new_n9833_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__25_));
AND2X2 AND2X2_3688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9837_), .B(AES_CORE_DATAPATH__abc_16009_new_n9836_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__26_));
AND2X2 AND2X2_3689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9840_), .B(AES_CORE_DATAPATH__abc_16009_new_n9839_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__27_));
AND2X2 AND2X2_369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2973_), .B(AES_CORE_DATAPATH__abc_16009_new_n2957_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__7_));
AND2X2 AND2X2_3690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9843_), .B(AES_CORE_DATAPATH__abc_16009_new_n9842_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__28_));
AND2X2 AND2X2_3691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9846_), .B(AES_CORE_DATAPATH__abc_16009_new_n9845_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__29_));
AND2X2 AND2X2_3692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9849_), .B(AES_CORE_DATAPATH__abc_16009_new_n9848_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__30_));
AND2X2 AND2X2_3693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9852_), .B(AES_CORE_DATAPATH__abc_16009_new_n9851_), .Y(AES_CORE_DATAPATH__0iv_1__31_0__31_));
AND2X2 AND2X2_3694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8525_), .B(AES_CORE_DATAPATH_col_en_host_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9854_));
AND2X2 AND2X2_3695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8528_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9855_));
AND2X2 AND2X2_3696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9858_));
AND2X2 AND2X2_3697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8273_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9859_));
AND2X2 AND2X2_3698 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9861_));
AND2X2 AND2X2_3699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8281_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9862_));
AND2X2 AND2X2_37 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_), .B(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n125_));
AND2X2 AND2X2_370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2975_));
AND2X2 AND2X2_3700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9864_));
AND2X2 AND2X2_3701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8289_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9865_));
AND2X2 AND2X2_3702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9867_));
AND2X2 AND2X2_3703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8297_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9868_));
AND2X2 AND2X2_3704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9870_));
AND2X2 AND2X2_3705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8305_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9871_));
AND2X2 AND2X2_3706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9873_));
AND2X2 AND2X2_3707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8313_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9874_));
AND2X2 AND2X2_3708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9876_));
AND2X2 AND2X2_3709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8321_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9877_));
AND2X2 AND2X2_371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2978_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2979_));
AND2X2 AND2X2_3710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9879_));
AND2X2 AND2X2_3711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8329_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9880_));
AND2X2 AND2X2_3712 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9882_));
AND2X2 AND2X2_3713 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8337_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9883_));
AND2X2 AND2X2_3714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9885_));
AND2X2 AND2X2_3715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8345_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9886_));
AND2X2 AND2X2_3716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9888_));
AND2X2 AND2X2_3717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8353_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9889_));
AND2X2 AND2X2_3718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9891_));
AND2X2 AND2X2_3719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8361_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9892_));
AND2X2 AND2X2_372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2981_));
AND2X2 AND2X2_3720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9894_));
AND2X2 AND2X2_3721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8369_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9895_));
AND2X2 AND2X2_3722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9897_));
AND2X2 AND2X2_3723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8377_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9898_));
AND2X2 AND2X2_3724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9900_));
AND2X2 AND2X2_3725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8385_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9901_));
AND2X2 AND2X2_3726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9903_));
AND2X2 AND2X2_3727 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8393_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9904_));
AND2X2 AND2X2_3728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9906_));
AND2X2 AND2X2_3729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8401_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9907_));
AND2X2 AND2X2_373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2982_));
AND2X2 AND2X2_3730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9909_));
AND2X2 AND2X2_3731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8409_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9910_));
AND2X2 AND2X2_3732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9912_));
AND2X2 AND2X2_3733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8417_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9913_));
AND2X2 AND2X2_3734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9915_));
AND2X2 AND2X2_3735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8425_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9916_));
AND2X2 AND2X2_3736 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9918_));
AND2X2 AND2X2_3737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8433_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9919_));
AND2X2 AND2X2_3738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9921_));
AND2X2 AND2X2_3739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8441_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9922_));
AND2X2 AND2X2_374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2984_), .B(AES_CORE_DATAPATH__abc_16009_new_n2985_), .Y(\key_out[8] ));
AND2X2 AND2X2_3740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9924_));
AND2X2 AND2X2_3741 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8449_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9925_));
AND2X2 AND2X2_3742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9927_));
AND2X2 AND2X2_3743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8457_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9928_));
AND2X2 AND2X2_3744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9930_));
AND2X2 AND2X2_3745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8465_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9931_));
AND2X2 AND2X2_3746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9933_));
AND2X2 AND2X2_3747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8473_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9934_));
AND2X2 AND2X2_3748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9936_));
AND2X2 AND2X2_3749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8481_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9937_));
AND2X2 AND2X2_375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2989_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2990_));
AND2X2 AND2X2_3750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9939_));
AND2X2 AND2X2_3751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8489_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9940_));
AND2X2 AND2X2_3752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9942_));
AND2X2 AND2X2_3753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8497_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9943_));
AND2X2 AND2X2_3754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9945_));
AND2X2 AND2X2_3755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8505_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9946_));
AND2X2 AND2X2_3756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9948_));
AND2X2 AND2X2_3757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8513_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9949_));
AND2X2 AND2X2_3758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH_bkp_1_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9951_));
AND2X2 AND2X2_3759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8521_), .B(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9952_));
AND2X2 AND2X2_376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2990_), .B(AES_CORE_DATAPATH__abc_16009_new_n2988_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2991_));
AND2X2 AND2X2_3760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9955_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9956_));
AND2X2 AND2X2_3761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9954_), .B(AES_CORE_DATAPATH__abc_16009_new_n9956_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9957_));
AND2X2 AND2X2_3762 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9959_), .B(AES_CORE_DATAPATH__abc_16009_new_n9960_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__0_));
AND2X2 AND2X2_3763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9963_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9964_));
AND2X2 AND2X2_3764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9962_), .B(AES_CORE_DATAPATH__abc_16009_new_n9964_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9965_));
AND2X2 AND2X2_3765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9967_), .B(AES_CORE_DATAPATH__abc_16009_new_n9968_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__1_));
AND2X2 AND2X2_3766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9971_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9972_));
AND2X2 AND2X2_3767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9970_), .B(AES_CORE_DATAPATH__abc_16009_new_n9972_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9973_));
AND2X2 AND2X2_3768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9975_), .B(AES_CORE_DATAPATH__abc_16009_new_n9976_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__2_));
AND2X2 AND2X2_3769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9979_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9980_));
AND2X2 AND2X2_377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n2996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2997_));
AND2X2 AND2X2_3770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9978_), .B(AES_CORE_DATAPATH__abc_16009_new_n9980_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9981_));
AND2X2 AND2X2_3771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9983_), .B(AES_CORE_DATAPATH__abc_16009_new_n9984_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__3_));
AND2X2 AND2X2_3772 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9987_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9988_));
AND2X2 AND2X2_3773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9986_), .B(AES_CORE_DATAPATH__abc_16009_new_n9988_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9989_));
AND2X2 AND2X2_3774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9991_), .B(AES_CORE_DATAPATH__abc_16009_new_n9992_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__4_));
AND2X2 AND2X2_3775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9995_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9996_));
AND2X2 AND2X2_3776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9994_), .B(AES_CORE_DATAPATH__abc_16009_new_n9996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9997_));
AND2X2 AND2X2_3777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9999_), .B(AES_CORE_DATAPATH__abc_16009_new_n10000_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__5_));
AND2X2 AND2X2_3778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10003_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10004_));
AND2X2 AND2X2_3779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10002_), .B(AES_CORE_DATAPATH__abc_16009_new_n10004_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10005_));
AND2X2 AND2X2_378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2999_));
AND2X2 AND2X2_3780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10007_), .B(AES_CORE_DATAPATH__abc_16009_new_n10008_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__6_));
AND2X2 AND2X2_3781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10011_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10012_));
AND2X2 AND2X2_3782 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10010_), .B(AES_CORE_DATAPATH__abc_16009_new_n10012_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10013_));
AND2X2 AND2X2_3783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10015_), .B(AES_CORE_DATAPATH__abc_16009_new_n10016_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__7_));
AND2X2 AND2X2_3784 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10019_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10020_));
AND2X2 AND2X2_3785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10018_), .B(AES_CORE_DATAPATH__abc_16009_new_n10020_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10021_));
AND2X2 AND2X2_3786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10023_), .B(AES_CORE_DATAPATH__abc_16009_new_n10024_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__8_));
AND2X2 AND2X2_3787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10027_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10028_));
AND2X2 AND2X2_3788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10026_), .B(AES_CORE_DATAPATH__abc_16009_new_n10028_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10029_));
AND2X2 AND2X2_3789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10031_), .B(AES_CORE_DATAPATH__abc_16009_new_n10032_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__9_));
AND2X2 AND2X2_379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3000_));
AND2X2 AND2X2_3790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10035_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10036_));
AND2X2 AND2X2_3791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10034_), .B(AES_CORE_DATAPATH__abc_16009_new_n10036_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10037_));
AND2X2 AND2X2_3792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10039_), .B(AES_CORE_DATAPATH__abc_16009_new_n10040_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__10_));
AND2X2 AND2X2_3793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10043_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10044_));
AND2X2 AND2X2_3794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10042_), .B(AES_CORE_DATAPATH__abc_16009_new_n10044_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10045_));
AND2X2 AND2X2_3795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10047_), .B(AES_CORE_DATAPATH__abc_16009_new_n10048_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__11_));
AND2X2 AND2X2_3796 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10051_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10052_));
AND2X2 AND2X2_3797 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10050_), .B(AES_CORE_DATAPATH__abc_16009_new_n10052_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10053_));
AND2X2 AND2X2_3798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10055_), .B(AES_CORE_DATAPATH__abc_16009_new_n10056_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__12_));
AND2X2 AND2X2_3799 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10059_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10060_));
AND2X2 AND2X2_38 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n129_));
AND2X2 AND2X2_380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3002_), .B(AES_CORE_DATAPATH__abc_16009_new_n3003_), .Y(\key_out[9] ));
AND2X2 AND2X2_3800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10058_), .B(AES_CORE_DATAPATH__abc_16009_new_n10060_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10061_));
AND2X2 AND2X2_3801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10063_), .B(AES_CORE_DATAPATH__abc_16009_new_n10064_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__13_));
AND2X2 AND2X2_3802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10067_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10068_));
AND2X2 AND2X2_3803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10066_), .B(AES_CORE_DATAPATH__abc_16009_new_n10068_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10069_));
AND2X2 AND2X2_3804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10071_), .B(AES_CORE_DATAPATH__abc_16009_new_n10072_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__14_));
AND2X2 AND2X2_3805 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10075_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10076_));
AND2X2 AND2X2_3806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10074_), .B(AES_CORE_DATAPATH__abc_16009_new_n10076_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10077_));
AND2X2 AND2X2_3807 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10079_), .B(AES_CORE_DATAPATH__abc_16009_new_n10080_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__15_));
AND2X2 AND2X2_3808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10083_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10084_));
AND2X2 AND2X2_3809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10082_), .B(AES_CORE_DATAPATH__abc_16009_new_n10084_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10085_));
AND2X2 AND2X2_381 ( .A(\key_out[9] ), .B(AES_CORE_DATAPATH__abc_16009_new_n2994_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3005_));
AND2X2 AND2X2_3810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10087_), .B(AES_CORE_DATAPATH__abc_16009_new_n10088_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__16_));
AND2X2 AND2X2_3811 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10091_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10092_));
AND2X2 AND2X2_3812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10090_), .B(AES_CORE_DATAPATH__abc_16009_new_n10092_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10093_));
AND2X2 AND2X2_3813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10095_), .B(AES_CORE_DATAPATH__abc_16009_new_n10096_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__17_));
AND2X2 AND2X2_3814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10099_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10100_));
AND2X2 AND2X2_3815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10098_), .B(AES_CORE_DATAPATH__abc_16009_new_n10100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10101_));
AND2X2 AND2X2_3816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10103_), .B(AES_CORE_DATAPATH__abc_16009_new_n10104_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__18_));
AND2X2 AND2X2_3817 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10107_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10108_));
AND2X2 AND2X2_3818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10106_), .B(AES_CORE_DATAPATH__abc_16009_new_n10108_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10109_));
AND2X2 AND2X2_3819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10111_), .B(AES_CORE_DATAPATH__abc_16009_new_n10112_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__19_));
AND2X2 AND2X2_382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3006_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3007_));
AND2X2 AND2X2_3820 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10115_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10116_));
AND2X2 AND2X2_3821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10114_), .B(AES_CORE_DATAPATH__abc_16009_new_n10116_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10117_));
AND2X2 AND2X2_3822 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10119_), .B(AES_CORE_DATAPATH__abc_16009_new_n10120_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__20_));
AND2X2 AND2X2_3823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10123_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10124_));
AND2X2 AND2X2_3824 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10122_), .B(AES_CORE_DATAPATH__abc_16009_new_n10124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10125_));
AND2X2 AND2X2_3825 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10127_), .B(AES_CORE_DATAPATH__abc_16009_new_n10128_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__21_));
AND2X2 AND2X2_3826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10131_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10132_));
AND2X2 AND2X2_3827 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10130_), .B(AES_CORE_DATAPATH__abc_16009_new_n10132_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10133_));
AND2X2 AND2X2_3828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10135_), .B(AES_CORE_DATAPATH__abc_16009_new_n10136_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__22_));
AND2X2 AND2X2_3829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10139_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10140_));
AND2X2 AND2X2_383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3009_), .B(AES_CORE_DATAPATH__abc_16009_new_n2993_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__9_));
AND2X2 AND2X2_3830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10138_), .B(AES_CORE_DATAPATH__abc_16009_new_n10140_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10141_));
AND2X2 AND2X2_3831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10143_), .B(AES_CORE_DATAPATH__abc_16009_new_n10144_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__23_));
AND2X2 AND2X2_3832 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10147_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10148_));
AND2X2 AND2X2_3833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10146_), .B(AES_CORE_DATAPATH__abc_16009_new_n10148_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10149_));
AND2X2 AND2X2_3834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10151_), .B(AES_CORE_DATAPATH__abc_16009_new_n10152_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__24_));
AND2X2 AND2X2_3835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10155_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10156_));
AND2X2 AND2X2_3836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10154_), .B(AES_CORE_DATAPATH__abc_16009_new_n10156_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10157_));
AND2X2 AND2X2_3837 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10159_), .B(AES_CORE_DATAPATH__abc_16009_new_n10160_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__25_));
AND2X2 AND2X2_3838 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10163_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10164_));
AND2X2 AND2X2_3839 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10162_), .B(AES_CORE_DATAPATH__abc_16009_new_n10164_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10165_));
AND2X2 AND2X2_384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3011_));
AND2X2 AND2X2_3840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10167_), .B(AES_CORE_DATAPATH__abc_16009_new_n10168_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__26_));
AND2X2 AND2X2_3841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10171_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10172_));
AND2X2 AND2X2_3842 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10170_), .B(AES_CORE_DATAPATH__abc_16009_new_n10172_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10173_));
AND2X2 AND2X2_3843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10175_), .B(AES_CORE_DATAPATH__abc_16009_new_n10176_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__27_));
AND2X2 AND2X2_3844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10179_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10180_));
AND2X2 AND2X2_3845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10178_), .B(AES_CORE_DATAPATH__abc_16009_new_n10180_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10181_));
AND2X2 AND2X2_3846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10183_), .B(AES_CORE_DATAPATH__abc_16009_new_n10184_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__28_));
AND2X2 AND2X2_3847 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10187_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10188_));
AND2X2 AND2X2_3848 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10186_), .B(AES_CORE_DATAPATH__abc_16009_new_n10188_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10189_));
AND2X2 AND2X2_3849 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10191_), .B(AES_CORE_DATAPATH__abc_16009_new_n10192_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__29_));
AND2X2 AND2X2_385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3015_));
AND2X2 AND2X2_3850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10195_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10196_));
AND2X2 AND2X2_3851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10194_), .B(AES_CORE_DATAPATH__abc_16009_new_n10196_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10197_));
AND2X2 AND2X2_3852 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10199_), .B(AES_CORE_DATAPATH__abc_16009_new_n10200_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__30_));
AND2X2 AND2X2_3853 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10203_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10204_));
AND2X2 AND2X2_3854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10202_), .B(AES_CORE_DATAPATH__abc_16009_new_n10204_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10205_));
AND2X2 AND2X2_3855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10207_), .B(AES_CORE_DATAPATH__abc_16009_new_n10208_), .Y(AES_CORE_DATAPATH__0bkp_1__31_0__31_));
AND2X2 AND2X2_3856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10212_), .B(AES_CORE_DATAPATH__abc_16009_new_n10210_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__0_));
AND2X2 AND2X2_3857 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10215_), .B(AES_CORE_DATAPATH__abc_16009_new_n10214_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__1_));
AND2X2 AND2X2_3858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10218_), .B(AES_CORE_DATAPATH__abc_16009_new_n10217_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__2_));
AND2X2 AND2X2_3859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10221_), .B(AES_CORE_DATAPATH__abc_16009_new_n10220_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__3_));
AND2X2 AND2X2_386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3017_));
AND2X2 AND2X2_3860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10224_), .B(AES_CORE_DATAPATH__abc_16009_new_n10223_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__4_));
AND2X2 AND2X2_3861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10227_), .B(AES_CORE_DATAPATH__abc_16009_new_n10226_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__5_));
AND2X2 AND2X2_3862 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10230_), .B(AES_CORE_DATAPATH__abc_16009_new_n10229_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__6_));
AND2X2 AND2X2_3863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10233_), .B(AES_CORE_DATAPATH__abc_16009_new_n10232_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__7_));
AND2X2 AND2X2_3864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10236_), .B(AES_CORE_DATAPATH__abc_16009_new_n10235_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__8_));
AND2X2 AND2X2_3865 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10239_), .B(AES_CORE_DATAPATH__abc_16009_new_n10238_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__9_));
AND2X2 AND2X2_3866 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10242_), .B(AES_CORE_DATAPATH__abc_16009_new_n10241_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__10_));
AND2X2 AND2X2_3867 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10245_), .B(AES_CORE_DATAPATH__abc_16009_new_n10244_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__11_));
AND2X2 AND2X2_3868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10248_), .B(AES_CORE_DATAPATH__abc_16009_new_n10247_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__12_));
AND2X2 AND2X2_3869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10251_), .B(AES_CORE_DATAPATH__abc_16009_new_n10250_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__13_));
AND2X2 AND2X2_387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3018_));
AND2X2 AND2X2_3870 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10254_), .B(AES_CORE_DATAPATH__abc_16009_new_n10253_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__14_));
AND2X2 AND2X2_3871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10257_), .B(AES_CORE_DATAPATH__abc_16009_new_n10256_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__15_));
AND2X2 AND2X2_3872 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10260_), .B(AES_CORE_DATAPATH__abc_16009_new_n10259_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__16_));
AND2X2 AND2X2_3873 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10263_), .B(AES_CORE_DATAPATH__abc_16009_new_n10262_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__17_));
AND2X2 AND2X2_3874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10266_), .B(AES_CORE_DATAPATH__abc_16009_new_n10265_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__18_));
AND2X2 AND2X2_3875 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10269_), .B(AES_CORE_DATAPATH__abc_16009_new_n10268_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__19_));
AND2X2 AND2X2_3876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10272_), .B(AES_CORE_DATAPATH__abc_16009_new_n10271_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__20_));
AND2X2 AND2X2_3877 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10275_), .B(AES_CORE_DATAPATH__abc_16009_new_n10274_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__21_));
AND2X2 AND2X2_3878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10278_), .B(AES_CORE_DATAPATH__abc_16009_new_n10277_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__22_));
AND2X2 AND2X2_3879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10281_), .B(AES_CORE_DATAPATH__abc_16009_new_n10280_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__23_));
AND2X2 AND2X2_388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3020_), .B(AES_CORE_DATAPATH__abc_16009_new_n3021_), .Y(\key_out[10] ));
AND2X2 AND2X2_3880 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10284_), .B(AES_CORE_DATAPATH__abc_16009_new_n10283_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__24_));
AND2X2 AND2X2_3881 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10287_), .B(AES_CORE_DATAPATH__abc_16009_new_n10286_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__25_));
AND2X2 AND2X2_3882 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10290_), .B(AES_CORE_DATAPATH__abc_16009_new_n10289_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__26_));
AND2X2 AND2X2_3883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10293_), .B(AES_CORE_DATAPATH__abc_16009_new_n10292_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__27_));
AND2X2 AND2X2_3884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10296_), .B(AES_CORE_DATAPATH__abc_16009_new_n10295_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__28_));
AND2X2 AND2X2_3885 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10299_), .B(AES_CORE_DATAPATH__abc_16009_new_n10298_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__29_));
AND2X2 AND2X2_3886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10302_), .B(AES_CORE_DATAPATH__abc_16009_new_n10301_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__30_));
AND2X2 AND2X2_3887 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10305_), .B(AES_CORE_DATAPATH__abc_16009_new_n10304_), .Y(AES_CORE_DATAPATH__0iv_0__31_0__31_));
AND2X2 AND2X2_3888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8525_), .B(AES_CORE_DATAPATH_col_en_host_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10307_));
AND2X2 AND2X2_3889 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8528_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10308_));
AND2X2 AND2X2_389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3025_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3026_));
AND2X2 AND2X2_3890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10311_));
AND2X2 AND2X2_3891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7759_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10312_));
AND2X2 AND2X2_3892 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10314_));
AND2X2 AND2X2_3893 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7767_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10315_));
AND2X2 AND2X2_3894 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10317_));
AND2X2 AND2X2_3895 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7775_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10318_));
AND2X2 AND2X2_3896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10320_));
AND2X2 AND2X2_3897 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7783_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10321_));
AND2X2 AND2X2_3898 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10323_));
AND2X2 AND2X2_3899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7791_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10324_));
AND2X2 AND2X2_39 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n127_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n129_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n130_));
AND2X2 AND2X2_390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3026_), .B(AES_CORE_DATAPATH__abc_16009_new_n3024_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3027_));
AND2X2 AND2X2_3900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10326_));
AND2X2 AND2X2_3901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7799_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10327_));
AND2X2 AND2X2_3902 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10329_));
AND2X2 AND2X2_3903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7807_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10330_));
AND2X2 AND2X2_3904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10332_));
AND2X2 AND2X2_3905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7815_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10333_));
AND2X2 AND2X2_3906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10335_));
AND2X2 AND2X2_3907 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7823_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10336_));
AND2X2 AND2X2_3908 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10338_));
AND2X2 AND2X2_3909 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7831_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10339_));
AND2X2 AND2X2_391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3032_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3033_));
AND2X2 AND2X2_3910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10341_));
AND2X2 AND2X2_3911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7839_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10342_));
AND2X2 AND2X2_3912 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10344_));
AND2X2 AND2X2_3913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7847_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10345_));
AND2X2 AND2X2_3914 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10347_));
AND2X2 AND2X2_3915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7855_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10348_));
AND2X2 AND2X2_3916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10350_));
AND2X2 AND2X2_3917 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7863_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10351_));
AND2X2 AND2X2_3918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10353_));
AND2X2 AND2X2_3919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7871_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10354_));
AND2X2 AND2X2_392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3035_));
AND2X2 AND2X2_3920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10356_));
AND2X2 AND2X2_3921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7879_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10357_));
AND2X2 AND2X2_3922 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10359_));
AND2X2 AND2X2_3923 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7887_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10360_));
AND2X2 AND2X2_3924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10362_));
AND2X2 AND2X2_3925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7895_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10363_));
AND2X2 AND2X2_3926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10365_));
AND2X2 AND2X2_3927 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7903_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10366_));
AND2X2 AND2X2_3928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10368_));
AND2X2 AND2X2_3929 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7911_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10369_));
AND2X2 AND2X2_393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3036_));
AND2X2 AND2X2_3930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10371_));
AND2X2 AND2X2_3931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7919_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10372_));
AND2X2 AND2X2_3932 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10374_));
AND2X2 AND2X2_3933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7927_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10375_));
AND2X2 AND2X2_3934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10377_));
AND2X2 AND2X2_3935 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7935_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10378_));
AND2X2 AND2X2_3936 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10380_));
AND2X2 AND2X2_3937 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7943_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10381_));
AND2X2 AND2X2_3938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10383_));
AND2X2 AND2X2_3939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7951_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10384_));
AND2X2 AND2X2_394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3038_), .B(AES_CORE_DATAPATH__abc_16009_new_n3039_), .Y(\key_out[11] ));
AND2X2 AND2X2_3940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10386_));
AND2X2 AND2X2_3941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7959_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10387_));
AND2X2 AND2X2_3942 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10389_));
AND2X2 AND2X2_3943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7967_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10390_));
AND2X2 AND2X2_3944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10392_));
AND2X2 AND2X2_3945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7975_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10393_));
AND2X2 AND2X2_3946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10395_));
AND2X2 AND2X2_3947 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7983_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10396_));
AND2X2 AND2X2_3948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10398_));
AND2X2 AND2X2_3949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7991_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10399_));
AND2X2 AND2X2_395 ( .A(\key_out[11] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3041_));
AND2X2 AND2X2_3950 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10401_));
AND2X2 AND2X2_3951 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7999_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10402_));
AND2X2 AND2X2_3952 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH_bkp_1_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10404_));
AND2X2 AND2X2_3953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8007_), .B(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10405_));
AND2X2 AND2X2_3954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10408_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10409_));
AND2X2 AND2X2_3955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10407_), .B(AES_CORE_DATAPATH__abc_16009_new_n10409_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10410_));
AND2X2 AND2X2_3956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10412_), .B(AES_CORE_DATAPATH__abc_16009_new_n10413_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__0_));
AND2X2 AND2X2_3957 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10416_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10417_));
AND2X2 AND2X2_3958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10415_), .B(AES_CORE_DATAPATH__abc_16009_new_n10417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10418_));
AND2X2 AND2X2_3959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10420_), .B(AES_CORE_DATAPATH__abc_16009_new_n10421_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__1_));
AND2X2 AND2X2_396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3042_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3043_));
AND2X2 AND2X2_3960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10424_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10425_));
AND2X2 AND2X2_3961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10423_), .B(AES_CORE_DATAPATH__abc_16009_new_n10425_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10426_));
AND2X2 AND2X2_3962 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10428_), .B(AES_CORE_DATAPATH__abc_16009_new_n10429_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__2_));
AND2X2 AND2X2_3963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10432_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10433_));
AND2X2 AND2X2_3964 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10431_), .B(AES_CORE_DATAPATH__abc_16009_new_n10433_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10434_));
AND2X2 AND2X2_3965 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10436_), .B(AES_CORE_DATAPATH__abc_16009_new_n10437_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__3_));
AND2X2 AND2X2_3966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10440_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10441_));
AND2X2 AND2X2_3967 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10439_), .B(AES_CORE_DATAPATH__abc_16009_new_n10441_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10442_));
AND2X2 AND2X2_3968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10444_), .B(AES_CORE_DATAPATH__abc_16009_new_n10445_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__4_));
AND2X2 AND2X2_3969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10448_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10449_));
AND2X2 AND2X2_397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3045_), .B(AES_CORE_DATAPATH__abc_16009_new_n3029_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__11_));
AND2X2 AND2X2_3970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10447_), .B(AES_CORE_DATAPATH__abc_16009_new_n10449_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10450_));
AND2X2 AND2X2_3971 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10452_), .B(AES_CORE_DATAPATH__abc_16009_new_n10453_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__5_));
AND2X2 AND2X2_3972 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10456_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10457_));
AND2X2 AND2X2_3973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10455_), .B(AES_CORE_DATAPATH__abc_16009_new_n10457_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10458_));
AND2X2 AND2X2_3974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10460_), .B(AES_CORE_DATAPATH__abc_16009_new_n10461_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__6_));
AND2X2 AND2X2_3975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10464_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10465_));
AND2X2 AND2X2_3976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10463_), .B(AES_CORE_DATAPATH__abc_16009_new_n10465_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10466_));
AND2X2 AND2X2_3977 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10468_), .B(AES_CORE_DATAPATH__abc_16009_new_n10469_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__7_));
AND2X2 AND2X2_3978 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10472_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10473_));
AND2X2 AND2X2_3979 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10471_), .B(AES_CORE_DATAPATH__abc_16009_new_n10473_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10474_));
AND2X2 AND2X2_398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3050_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3051_));
AND2X2 AND2X2_3980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10476_), .B(AES_CORE_DATAPATH__abc_16009_new_n10477_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__8_));
AND2X2 AND2X2_3981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10480_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10481_));
AND2X2 AND2X2_3982 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10479_), .B(AES_CORE_DATAPATH__abc_16009_new_n10481_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10482_));
AND2X2 AND2X2_3983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10484_), .B(AES_CORE_DATAPATH__abc_16009_new_n10485_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__9_));
AND2X2 AND2X2_3984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10488_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10489_));
AND2X2 AND2X2_3985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10487_), .B(AES_CORE_DATAPATH__abc_16009_new_n10489_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10490_));
AND2X2 AND2X2_3986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10492_), .B(AES_CORE_DATAPATH__abc_16009_new_n10493_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__10_));
AND2X2 AND2X2_3987 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10496_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10497_));
AND2X2 AND2X2_3988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10495_), .B(AES_CORE_DATAPATH__abc_16009_new_n10497_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10498_));
AND2X2 AND2X2_3989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10500_), .B(AES_CORE_DATAPATH__abc_16009_new_n10501_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__11_));
AND2X2 AND2X2_399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3053_));
AND2X2 AND2X2_3990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10504_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10505_));
AND2X2 AND2X2_3991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10503_), .B(AES_CORE_DATAPATH__abc_16009_new_n10505_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10506_));
AND2X2 AND2X2_3992 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10508_), .B(AES_CORE_DATAPATH__abc_16009_new_n10509_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__12_));
AND2X2 AND2X2_3993 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10512_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10513_));
AND2X2 AND2X2_3994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10511_), .B(AES_CORE_DATAPATH__abc_16009_new_n10513_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10514_));
AND2X2 AND2X2_3995 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10516_), .B(AES_CORE_DATAPATH__abc_16009_new_n10517_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__13_));
AND2X2 AND2X2_3996 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10520_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10521_));
AND2X2 AND2X2_3997 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10519_), .B(AES_CORE_DATAPATH__abc_16009_new_n10521_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10522_));
AND2X2 AND2X2_3998 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10524_), .B(AES_CORE_DATAPATH__abc_16009_new_n10525_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__14_));
AND2X2 AND2X2_3999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10528_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10529_));
AND2X2 AND2X2_4 ( .A(_abc_15574_new_n15_), .B(_abc_15574_new_n11_), .Y(AES_CORE_DATAPATH_col_en_host_1_));
AND2X2 AND2X2_40 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n130_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n131_));
AND2X2 AND2X2_400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3054_));
AND2X2 AND2X2_4000 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10527_), .B(AES_CORE_DATAPATH__abc_16009_new_n10529_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10530_));
AND2X2 AND2X2_4001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10532_), .B(AES_CORE_DATAPATH__abc_16009_new_n10533_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__15_));
AND2X2 AND2X2_4002 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10536_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10537_));
AND2X2 AND2X2_4003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10535_), .B(AES_CORE_DATAPATH__abc_16009_new_n10537_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10538_));
AND2X2 AND2X2_4004 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10540_), .B(AES_CORE_DATAPATH__abc_16009_new_n10541_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__16_));
AND2X2 AND2X2_4005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10544_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10545_));
AND2X2 AND2X2_4006 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10543_), .B(AES_CORE_DATAPATH__abc_16009_new_n10545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10546_));
AND2X2 AND2X2_4007 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10548_), .B(AES_CORE_DATAPATH__abc_16009_new_n10549_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__17_));
AND2X2 AND2X2_4008 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10552_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10553_));
AND2X2 AND2X2_4009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10551_), .B(AES_CORE_DATAPATH__abc_16009_new_n10553_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10554_));
AND2X2 AND2X2_401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3056_), .B(AES_CORE_DATAPATH__abc_16009_new_n3057_), .Y(\key_out[12] ));
AND2X2 AND2X2_4010 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10556_), .B(AES_CORE_DATAPATH__abc_16009_new_n10557_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__18_));
AND2X2 AND2X2_4011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10560_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10561_));
AND2X2 AND2X2_4012 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10559_), .B(AES_CORE_DATAPATH__abc_16009_new_n10561_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10562_));
AND2X2 AND2X2_4013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10564_), .B(AES_CORE_DATAPATH__abc_16009_new_n10565_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__19_));
AND2X2 AND2X2_4014 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10568_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10569_));
AND2X2 AND2X2_4015 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10567_), .B(AES_CORE_DATAPATH__abc_16009_new_n10569_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10570_));
AND2X2 AND2X2_4016 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10572_), .B(AES_CORE_DATAPATH__abc_16009_new_n10573_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__20_));
AND2X2 AND2X2_4017 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10576_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10577_));
AND2X2 AND2X2_4018 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10575_), .B(AES_CORE_DATAPATH__abc_16009_new_n10577_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10578_));
AND2X2 AND2X2_4019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10580_), .B(AES_CORE_DATAPATH__abc_16009_new_n10581_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__21_));
AND2X2 AND2X2_402 ( .A(\key_out[12] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3048_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3059_));
AND2X2 AND2X2_4020 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10584_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10585_));
AND2X2 AND2X2_4021 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10583_), .B(AES_CORE_DATAPATH__abc_16009_new_n10585_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10586_));
AND2X2 AND2X2_4022 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10588_), .B(AES_CORE_DATAPATH__abc_16009_new_n10589_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__22_));
AND2X2 AND2X2_4023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10592_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10593_));
AND2X2 AND2X2_4024 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10591_), .B(AES_CORE_DATAPATH__abc_16009_new_n10593_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10594_));
AND2X2 AND2X2_4025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10596_), .B(AES_CORE_DATAPATH__abc_16009_new_n10597_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__23_));
AND2X2 AND2X2_4026 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10600_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10601_));
AND2X2 AND2X2_4027 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10599_), .B(AES_CORE_DATAPATH__abc_16009_new_n10601_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10602_));
AND2X2 AND2X2_4028 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10604_), .B(AES_CORE_DATAPATH__abc_16009_new_n10605_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__24_));
AND2X2 AND2X2_4029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10608_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10609_));
AND2X2 AND2X2_403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3060_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3061_));
AND2X2 AND2X2_4030 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10607_), .B(AES_CORE_DATAPATH__abc_16009_new_n10609_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10610_));
AND2X2 AND2X2_4031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10612_), .B(AES_CORE_DATAPATH__abc_16009_new_n10613_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__25_));
AND2X2 AND2X2_4032 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10616_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10617_));
AND2X2 AND2X2_4033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10615_), .B(AES_CORE_DATAPATH__abc_16009_new_n10617_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10618_));
AND2X2 AND2X2_4034 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10620_), .B(AES_CORE_DATAPATH__abc_16009_new_n10621_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__26_));
AND2X2 AND2X2_4035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10624_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10625_));
AND2X2 AND2X2_4036 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10623_), .B(AES_CORE_DATAPATH__abc_16009_new_n10625_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10626_));
AND2X2 AND2X2_4037 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10628_), .B(AES_CORE_DATAPATH__abc_16009_new_n10629_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__27_));
AND2X2 AND2X2_4038 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10632_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10633_));
AND2X2 AND2X2_4039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10631_), .B(AES_CORE_DATAPATH__abc_16009_new_n10633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10634_));
AND2X2 AND2X2_404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3063_), .B(AES_CORE_DATAPATH__abc_16009_new_n3047_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__12_));
AND2X2 AND2X2_4040 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10636_), .B(AES_CORE_DATAPATH__abc_16009_new_n10637_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__28_));
AND2X2 AND2X2_4041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10640_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10641_));
AND2X2 AND2X2_4042 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10639_), .B(AES_CORE_DATAPATH__abc_16009_new_n10641_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10642_));
AND2X2 AND2X2_4043 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10644_), .B(AES_CORE_DATAPATH__abc_16009_new_n10645_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__29_));
AND2X2 AND2X2_4044 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10648_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10649_));
AND2X2 AND2X2_4045 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10647_), .B(AES_CORE_DATAPATH__abc_16009_new_n10649_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10650_));
AND2X2 AND2X2_4046 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10652_), .B(AES_CORE_DATAPATH__abc_16009_new_n10653_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__30_));
AND2X2 AND2X2_4047 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10656_), .B(AES_CORE_DATAPATH__abc_16009_new_n2802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10657_));
AND2X2 AND2X2_4048 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10655_), .B(AES_CORE_DATAPATH__abc_16009_new_n10657_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10658_));
AND2X2 AND2X2_4049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10660_), .B(AES_CORE_DATAPATH__abc_16009_new_n10661_), .Y(AES_CORE_DATAPATH__0bkp_0__31_0__31_));
AND2X2 AND2X2_405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3069_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3070_));
AND2X2 AND2X2_4050 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10664_), .B(AES_CORE_DATAPATH__abc_16009_new_n10663_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__0_));
AND2X2 AND2X2_4051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10667_), .B(AES_CORE_DATAPATH__abc_16009_new_n10666_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__1_));
AND2X2 AND2X2_4052 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10670_), .B(AES_CORE_DATAPATH__abc_16009_new_n10669_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__2_));
AND2X2 AND2X2_4053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10673_), .B(AES_CORE_DATAPATH__abc_16009_new_n10672_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__3_));
AND2X2 AND2X2_4054 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10676_), .B(AES_CORE_DATAPATH__abc_16009_new_n10675_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__0_));
AND2X2 AND2X2_4055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10679_), .B(AES_CORE_DATAPATH__abc_16009_new_n10678_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__1_));
AND2X2 AND2X2_4056 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10682_), .B(AES_CORE_DATAPATH__abc_16009_new_n10681_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__2_));
AND2X2 AND2X2_4057 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10685_), .B(AES_CORE_DATAPATH__abc_16009_new_n10684_), .Y(AES_CORE_DATAPATH__0key_en_pp1_3_0__3_));
AND2X2 AND2X2_4058 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10688_), .B(AES_CORE_DATAPATH__abc_16009_new_n10687_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__0_));
AND2X2 AND2X2_4059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10691_), .B(AES_CORE_DATAPATH__abc_16009_new_n10690_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__1_));
AND2X2 AND2X2_406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3072_));
AND2X2 AND2X2_4060 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10694_), .B(AES_CORE_DATAPATH__abc_16009_new_n10693_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__2_));
AND2X2 AND2X2_4061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10697_), .B(AES_CORE_DATAPATH__abc_16009_new_n10696_), .Y(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__3_));
AND2X2 AND2X2_4062 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out));
AND2X2 AND2X2_4063 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n328_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n330_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n331_));
AND2X2 AND2X2_4064 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n333_));
AND2X2 AND2X2_4065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n334_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n336_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_));
AND2X2 AND2X2_4066 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n339_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n341_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n342_));
AND2X2 AND2X2_4067 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n344_));
AND2X2 AND2X2_4068 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n345_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n347_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_));
AND2X2 AND2X2_4069 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n350_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n352_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n353_));
AND2X2 AND2X2_407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3073_));
AND2X2 AND2X2_4070 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n355_));
AND2X2 AND2X2_4071 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n356_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n358_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_));
AND2X2 AND2X2_4072 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n361_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n363_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n364_));
AND2X2 AND2X2_4073 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n366_));
AND2X2 AND2X2_4074 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n367_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n369_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_));
AND2X2 AND2X2_4075 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n372_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n374_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n375_));
AND2X2 AND2X2_4076 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n377_));
AND2X2 AND2X2_4077 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n378_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n380_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_));
AND2X2 AND2X2_4078 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n383_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n385_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n386_));
AND2X2 AND2X2_4079 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n388_));
AND2X2 AND2X2_408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3075_), .B(AES_CORE_DATAPATH__abc_16009_new_n3067_), .Y(\key_out[13] ));
AND2X2 AND2X2_4080 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n389_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n391_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_));
AND2X2 AND2X2_4081 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n394_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n396_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n397_));
AND2X2 AND2X2_4082 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n399_));
AND2X2 AND2X2_4083 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n400_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n402_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_));
AND2X2 AND2X2_4084 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n405_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n407_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n408_));
AND2X2 AND2X2_4085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n410_));
AND2X2 AND2X2_4086 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n411_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n413_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_));
AND2X2 AND2X2_4087 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n416_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n418_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n419_));
AND2X2 AND2X2_4088 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n421_));
AND2X2 AND2X2_4089 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n422_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n424_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_));
AND2X2 AND2X2_409 ( .A(\key_out[13] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3066_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3077_));
AND2X2 AND2X2_4090 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n427_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n429_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n430_));
AND2X2 AND2X2_4091 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n432_));
AND2X2 AND2X2_4092 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n433_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n435_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_));
AND2X2 AND2X2_4093 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n438_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n440_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n441_));
AND2X2 AND2X2_4094 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n443_));
AND2X2 AND2X2_4095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n444_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n446_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_));
AND2X2 AND2X2_4096 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n449_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n451_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n452_));
AND2X2 AND2X2_4097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n454_));
AND2X2 AND2X2_4098 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n455_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n457_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_));
AND2X2 AND2X2_4099 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n460_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n462_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n463_));
AND2X2 AND2X2_41 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n133_));
AND2X2 AND2X2_410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3078_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3079_));
AND2X2 AND2X2_4100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n465_));
AND2X2 AND2X2_4101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n466_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n468_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_));
AND2X2 AND2X2_4102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n471_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n473_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n474_));
AND2X2 AND2X2_4103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n476_));
AND2X2 AND2X2_4104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n477_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n479_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_));
AND2X2 AND2X2_4105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n482_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n484_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n485_));
AND2X2 AND2X2_4106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n487_));
AND2X2 AND2X2_4107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n488_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n490_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_));
AND2X2 AND2X2_4108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n493_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n495_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n496_));
AND2X2 AND2X2_4109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n498_));
AND2X2 AND2X2_411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3081_), .B(AES_CORE_DATAPATH__abc_16009_new_n3065_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__13_));
AND2X2 AND2X2_4110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n499_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n501_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_));
AND2X2 AND2X2_4111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n504_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n506_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n507_));
AND2X2 AND2X2_4112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n509_));
AND2X2 AND2X2_4113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n510_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n512_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_));
AND2X2 AND2X2_4114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n515_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n517_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n518_));
AND2X2 AND2X2_4115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n520_));
AND2X2 AND2X2_4116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n521_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n523_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_));
AND2X2 AND2X2_4117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n526_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n528_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n529_));
AND2X2 AND2X2_4118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n531_));
AND2X2 AND2X2_4119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n532_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n534_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_));
AND2X2 AND2X2_412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3087_));
AND2X2 AND2X2_4120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n537_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n539_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n540_));
AND2X2 AND2X2_4121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n542_));
AND2X2 AND2X2_4122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n543_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n545_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_));
AND2X2 AND2X2_4123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n548_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n550_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n551_));
AND2X2 AND2X2_4124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n553_));
AND2X2 AND2X2_4125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n554_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n556_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_));
AND2X2 AND2X2_4126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n559_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n561_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n562_));
AND2X2 AND2X2_4127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n564_));
AND2X2 AND2X2_4128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n565_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n567_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_));
AND2X2 AND2X2_4129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n570_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n572_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n573_));
AND2X2 AND2X2_413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3089_));
AND2X2 AND2X2_4130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n575_));
AND2X2 AND2X2_4131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n578_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_));
AND2X2 AND2X2_4132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n581_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n583_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n584_));
AND2X2 AND2X2_4133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n586_));
AND2X2 AND2X2_4134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n587_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n589_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_));
AND2X2 AND2X2_4135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n592_));
AND2X2 AND2X2_4136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n593_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n591_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n594_));
AND2X2 AND2X2_4137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n595_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n596_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n597_));
AND2X2 AND2X2_4138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n599_));
AND2X2 AND2X2_4139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n600_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n601_));
AND2X2 AND2X2_414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3090_));
AND2X2 AND2X2_4140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n602_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n597_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n603_));
AND2X2 AND2X2_4141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n605_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n607_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n608_));
AND2X2 AND2X2_4142 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n609_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n610_));
AND2X2 AND2X2_4143 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n611_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n594_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n612_));
AND2X2 AND2X2_4144 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n610_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n613_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n614_));
AND2X2 AND2X2_4145 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n617_));
AND2X2 AND2X2_4146 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n618_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n616_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n619_));
AND2X2 AND2X2_4147 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n597_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n600_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n622_));
AND2X2 AND2X2_4148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n596_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n623_));
AND2X2 AND2X2_4149 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n625_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n623_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n626_));
AND2X2 AND2X2_415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3092_), .B(AES_CORE_DATAPATH__abc_16009_new_n3093_), .Y(\key_out[14] ));
AND2X2 AND2X2_4150 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n623_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n595_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n629_));
AND2X2 AND2X2_4151 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n596_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n600_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n630_));
AND2X2 AND2X2_4152 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n595_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n631_));
AND2X2 AND2X2_4153 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n630_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n631_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n632_));
AND2X2 AND2X2_4154 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n628_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n634_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n635_));
AND2X2 AND2X2_4155 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n635_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n621_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n636_));
AND2X2 AND2X2_4156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n639_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n640_));
AND2X2 AND2X2_4157 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n640_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n620_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n641_));
AND2X2 AND2X2_4158 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n643_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n637_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n644_));
AND2X2 AND2X2_4159 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n645_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n619_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n646_));
AND2X2 AND2X2_416 ( .A(\key_out[14] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3084_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3095_));
AND2X2 AND2X2_4160 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n649_));
AND2X2 AND2X2_4161 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n650_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n648_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n651_));
AND2X2 AND2X2_4162 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n654_));
AND2X2 AND2X2_4163 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n655_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n656_));
AND2X2 AND2X2_4164 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n656_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n654_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n657_));
AND2X2 AND2X2_4165 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n659_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n660_));
AND2X2 AND2X2_4166 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n661_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n658_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n662_));
AND2X2 AND2X2_4167 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n600_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n663_));
AND2X2 AND2X2_4168 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n625_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n663_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n664_));
AND2X2 AND2X2_4169 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n667_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n668_));
AND2X2 AND2X2_417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3096_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3097_));
AND2X2 AND2X2_4170 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n669_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n665_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n670_));
AND2X2 AND2X2_4171 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n625_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n630_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n673_));
AND2X2 AND2X2_4172 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n597_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n677_));
AND2X2 AND2X2_4173 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n678_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n676_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n679_));
AND2X2 AND2X2_4174 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n680_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n675_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n681_));
AND2X2 AND2X2_4175 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n682_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n672_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n683_));
AND2X2 AND2X2_4176 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n683_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n684_));
AND2X2 AND2X2_4177 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n684_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n652_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n685_));
AND2X2 AND2X2_4178 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n681_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n686_));
AND2X2 AND2X2_4179 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n671_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n653_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n687_));
AND2X2 AND2X2_418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3099_), .B(AES_CORE_DATAPATH__abc_16009_new_n3083_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__14_));
AND2X2 AND2X2_4180 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n689_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n651_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n690_));
AND2X2 AND2X2_4181 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n693_));
AND2X2 AND2X2_4182 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n694_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n692_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n695_));
AND2X2 AND2X2_4183 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n656_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n663_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n697_));
AND2X2 AND2X2_4184 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n625_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n654_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n699_));
AND2X2 AND2X2_4185 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n698_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n700_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n701_));
AND2X2 AND2X2_4186 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n701_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n702_));
AND2X2 AND2X2_4187 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n703_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n704_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n705_));
AND2X2 AND2X2_4188 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n705_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n706_));
AND2X2 AND2X2_4189 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n706_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n696_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n707_));
AND2X2 AND2X2_419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3105_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3106_));
AND2X2 AND2X2_4190 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n710_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n695_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n711_));
AND2X2 AND2X2_4191 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n714_));
AND2X2 AND2X2_4192 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n715_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n713_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n716_));
AND2X2 AND2X2_4193 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n623_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n656_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n718_));
AND2X2 AND2X2_4194 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n660_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n719_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n720_));
AND2X2 AND2X2_4195 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n630_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n656_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n721_));
AND2X2 AND2X2_4196 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n668_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n722_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n723_));
AND2X2 AND2X2_4197 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n725_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n717_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n726_));
AND2X2 AND2X2_4198 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n724_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n727_));
AND2X2 AND2X2_4199 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n728_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n729_));
AND2X2 AND2X2_42 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n135_));
AND2X2 AND2X2_420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3108_));
AND2X2 AND2X2_4200 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n730_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n716_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n731_));
AND2X2 AND2X2_4201 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n729_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n732_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n733_));
AND2X2 AND2X2_4202 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n736_));
AND2X2 AND2X2_4203 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n737_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n735_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n738_));
AND2X2 AND2X2_4204 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n661_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n722_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n741_));
AND2X2 AND2X2_4205 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n669_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n719_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n742_));
AND2X2 AND2X2_4206 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n747_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n746_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n748_));
AND2X2 AND2X2_4207 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n749_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n744_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n750_));
AND2X2 AND2X2_4208 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n750_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n751_));
AND2X2 AND2X2_4209 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n751_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n739_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n752_));
AND2X2 AND2X2_421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3109_));
AND2X2 AND2X2_4210 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n748_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n753_));
AND2X2 AND2X2_4211 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n743_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n740_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n754_));
AND2X2 AND2X2_4212 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n756_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n738_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n757_));
AND2X2 AND2X2_4213 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n760_));
AND2X2 AND2X2_4214 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n761_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n759_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n762_));
AND2X2 AND2X2_4215 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n764_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n765_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n766_));
AND2X2 AND2X2_4216 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n766_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n767_));
AND2X2 AND2X2_4217 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n768_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n769_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n770_));
AND2X2 AND2X2_4218 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n770_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n771_));
AND2X2 AND2X2_4219 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n771_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n763_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n772_));
AND2X2 AND2X2_422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3111_), .B(AES_CORE_DATAPATH__abc_16009_new_n3103_), .Y(\key_out[15] ));
AND2X2 AND2X2_4220 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n773_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n762_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n774_));
AND2X2 AND2X2_4221 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n777_));
AND2X2 AND2X2_4222 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n778_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n776_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n779_));
AND2X2 AND2X2_4223 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n782_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n781_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n783_));
AND2X2 AND2X2_4224 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n784_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n785_));
AND2X2 AND2X2_4225 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n786_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n787_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n788_));
AND2X2 AND2X2_4226 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n788_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n789_));
AND2X2 AND2X2_4227 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n789_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n780_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n790_));
AND2X2 AND2X2_4228 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n793_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n779_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n794_));
AND2X2 AND2X2_4229 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n797_));
AND2X2 AND2X2_423 ( .A(\key_out[15] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3113_));
AND2X2 AND2X2_4230 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n798_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n796_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_));
AND2X2 AND2X2_4231 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n800_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n801_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_));
AND2X2 AND2X2_4232 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n804_));
AND2X2 AND2X2_4233 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n803_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_));
AND2X2 AND2X2_4234 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n807_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n808_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_));
AND2X2 AND2X2_4235 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n811_));
AND2X2 AND2X2_4236 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n812_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n810_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_));
AND2X2 AND2X2_4237 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n814_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n815_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_));
AND2X2 AND2X2_4238 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n818_));
AND2X2 AND2X2_4239 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n819_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n817_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_));
AND2X2 AND2X2_424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3115_));
AND2X2 AND2X2_4240 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n821_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n822_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_));
AND2X2 AND2X2_4241 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n825_));
AND2X2 AND2X2_4242 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n826_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n824_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_));
AND2X2 AND2X2_4243 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n829_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_));
AND2X2 AND2X2_4244 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n832_));
AND2X2 AND2X2_4245 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n833_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n831_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_));
AND2X2 AND2X2_4246 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n835_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n836_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_));
AND2X2 AND2X2_4247 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n839_));
AND2X2 AND2X2_4248 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n840_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n838_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_));
AND2X2 AND2X2_4249 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n842_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n843_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_));
AND2X2 AND2X2_425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3117_), .B(AES_CORE_DATAPATH__abc_16009_new_n3101_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__15_));
AND2X2 AND2X2_4250 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n846_));
AND2X2 AND2X2_4251 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n847_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n845_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_));
AND2X2 AND2X2_4252 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n849_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n850_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_));
AND2X2 AND2X2_4253 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n853_));
AND2X2 AND2X2_4254 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n854_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n852_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_));
AND2X2 AND2X2_4255 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n856_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n857_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_));
AND2X2 AND2X2_4256 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n860_));
AND2X2 AND2X2_4257 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n861_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n859_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_));
AND2X2 AND2X2_4258 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n863_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n864_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_));
AND2X2 AND2X2_4259 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n867_));
AND2X2 AND2X2_426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3119_));
AND2X2 AND2X2_4260 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n868_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n866_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_));
AND2X2 AND2X2_4261 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n870_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n871_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_));
AND2X2 AND2X2_4262 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n874_));
AND2X2 AND2X2_4263 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n875_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n873_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_));
AND2X2 AND2X2_4264 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n877_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n878_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_));
AND2X2 AND2X2_4265 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n881_));
AND2X2 AND2X2_4266 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n882_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n880_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_));
AND2X2 AND2X2_4267 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n884_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n885_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_));
AND2X2 AND2X2_4268 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n888_));
AND2X2 AND2X2_4269 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n889_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n887_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_));
AND2X2 AND2X2_427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3123_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3124_));
AND2X2 AND2X2_4270 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n891_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n892_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_));
AND2X2 AND2X2_4271 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n895_));
AND2X2 AND2X2_4272 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n896_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n894_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_));
AND2X2 AND2X2_4273 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n898_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n899_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_));
AND2X2 AND2X2_4274 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n902_));
AND2X2 AND2X2_4275 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n903_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n901_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_));
AND2X2 AND2X2_4276 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n905_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n906_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_));
AND2X2 AND2X2_4277 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n909_));
AND2X2 AND2X2_4278 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n910_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n908_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_));
AND2X2 AND2X2_4279 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n912_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n913_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_));
AND2X2 AND2X2_428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3126_));
AND2X2 AND2X2_4280 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n916_));
AND2X2 AND2X2_4281 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n917_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n915_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_));
AND2X2 AND2X2_4282 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n919_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n920_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_));
AND2X2 AND2X2_4283 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n923_));
AND2X2 AND2X2_4284 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n924_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n922_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_));
AND2X2 AND2X2_4285 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n926_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n927_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_));
AND2X2 AND2X2_4286 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n930_));
AND2X2 AND2X2_4287 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n931_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n929_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_));
AND2X2 AND2X2_4288 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n933_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n934_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_));
AND2X2 AND2X2_4289 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n937_));
AND2X2 AND2X2_429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3127_));
AND2X2 AND2X2_4290 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n938_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n936_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_));
AND2X2 AND2X2_4291 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n940_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n941_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_));
AND2X2 AND2X2_4292 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n944_));
AND2X2 AND2X2_4293 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n945_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n943_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_));
AND2X2 AND2X2_4294 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n947_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n948_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_));
AND2X2 AND2X2_4295 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n951_));
AND2X2 AND2X2_4296 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n952_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n950_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_));
AND2X2 AND2X2_4297 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n954_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n955_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_));
AND2X2 AND2X2_4298 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n958_));
AND2X2 AND2X2_4299 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n959_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n957_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_));
AND2X2 AND2X2_43 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n136_));
AND2X2 AND2X2_430 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3129_), .B(AES_CORE_DATAPATH__abc_16009_new_n3121_), .Y(\key_out[16] ));
AND2X2 AND2X2_4300 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n961_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n962_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_));
AND2X2 AND2X2_4301 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n965_));
AND2X2 AND2X2_4302 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n966_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n964_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_));
AND2X2 AND2X2_4303 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n968_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n969_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_));
AND2X2 AND2X2_4304 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n972_));
AND2X2 AND2X2_4305 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n973_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n971_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_));
AND2X2 AND2X2_4306 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n975_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n976_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_));
AND2X2 AND2X2_4307 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n979_));
AND2X2 AND2X2_4308 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n980_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n978_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_));
AND2X2 AND2X2_4309 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n982_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n983_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_));
AND2X2 AND2X2_431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3133_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3134_));
AND2X2 AND2X2_4310 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n986_));
AND2X2 AND2X2_4311 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n987_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n985_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_));
AND2X2 AND2X2_4312 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n989_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n990_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_));
AND2X2 AND2X2_4313 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n993_));
AND2X2 AND2X2_4314 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n994_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n992_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_));
AND2X2 AND2X2_4315 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n996_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n997_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_));
AND2X2 AND2X2_4316 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1000_));
AND2X2 AND2X2_4317 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1001_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n999_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_));
AND2X2 AND2X2_4318 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1003_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1004_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_));
AND2X2 AND2X2_4319 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1007_));
AND2X2 AND2X2_432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3134_), .B(AES_CORE_DATAPATH__abc_16009_new_n3132_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3135_));
AND2X2 AND2X2_4320 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1008_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1006_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_));
AND2X2 AND2X2_4321 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1010_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1011_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_));
AND2X2 AND2X2_4322 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1014_));
AND2X2 AND2X2_4323 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1015_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1013_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_));
AND2X2 AND2X2_4324 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1017_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1018_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_));
AND2X2 AND2X2_4325 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1021_));
AND2X2 AND2X2_4326 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1022_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1020_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_96_));
AND2X2 AND2X2_4327 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1025_));
AND2X2 AND2X2_4328 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1026_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1024_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_));
AND2X2 AND2X2_4329 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1029_));
AND2X2 AND2X2_433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3141_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3142_));
AND2X2 AND2X2_4330 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1030_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1028_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_));
AND2X2 AND2X2_4331 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1033_));
AND2X2 AND2X2_4332 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1034_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1032_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_));
AND2X2 AND2X2_4333 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1037_));
AND2X2 AND2X2_4334 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1038_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1036_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_));
AND2X2 AND2X2_4335 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1041_));
AND2X2 AND2X2_4336 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1042_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1040_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_));
AND2X2 AND2X2_4337 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1045_));
AND2X2 AND2X2_4338 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1046_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1044_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_));
AND2X2 AND2X2_4339 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1049_));
AND2X2 AND2X2_434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3144_));
AND2X2 AND2X2_4340 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1050_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1048_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_));
AND2X2 AND2X2_4341 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1053_));
AND2X2 AND2X2_4342 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1054_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1052_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_));
AND2X2 AND2X2_4343 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1057_));
AND2X2 AND2X2_4344 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1058_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1056_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_));
AND2X2 AND2X2_4345 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1061_));
AND2X2 AND2X2_4346 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1062_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1060_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_));
AND2X2 AND2X2_4347 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1065_));
AND2X2 AND2X2_4348 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1066_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1064_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_));
AND2X2 AND2X2_4349 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1069_));
AND2X2 AND2X2_435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3145_));
AND2X2 AND2X2_4350 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1070_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1068_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_));
AND2X2 AND2X2_4351 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1073_));
AND2X2 AND2X2_4352 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1074_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1072_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_));
AND2X2 AND2X2_4353 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1077_));
AND2X2 AND2X2_4354 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1078_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1076_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_));
AND2X2 AND2X2_4355 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1081_));
AND2X2 AND2X2_4356 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1082_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1080_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_));
AND2X2 AND2X2_4357 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1085_));
AND2X2 AND2X2_4358 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1086_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1084_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_));
AND2X2 AND2X2_4359 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1089_));
AND2X2 AND2X2_436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3147_), .B(AES_CORE_DATAPATH__abc_16009_new_n3139_), .Y(\key_out[17] ));
AND2X2 AND2X2_4360 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1090_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1088_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_));
AND2X2 AND2X2_4361 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1093_));
AND2X2 AND2X2_4362 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1094_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1092_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_));
AND2X2 AND2X2_4363 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1097_));
AND2X2 AND2X2_4364 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1098_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1096_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_));
AND2X2 AND2X2_4365 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1101_));
AND2X2 AND2X2_4366 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1102_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1100_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_));
AND2X2 AND2X2_4367 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1105_));
AND2X2 AND2X2_4368 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1106_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1104_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_));
AND2X2 AND2X2_4369 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1109_));
AND2X2 AND2X2_437 ( .A(\key_out[17] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3138_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3149_));
AND2X2 AND2X2_4370 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1110_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1108_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_));
AND2X2 AND2X2_4371 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1113_));
AND2X2 AND2X2_4372 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1114_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1112_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_));
AND2X2 AND2X2_4373 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n609_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1116_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1117_));
AND2X2 AND2X2_4374 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n608_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1118_));
AND2X2 AND2X2_4375 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1122_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1121_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_));
AND2X2 AND2X2_4376 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1125_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1126_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_));
AND2X2 AND2X2_4377 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1129_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1130_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_));
AND2X2 AND2X2_4378 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n728_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1132_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1133_));
AND2X2 AND2X2_4379 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1134_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1135_));
AND2X2 AND2X2_438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3150_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3151_));
AND2X2 AND2X2_4380 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1138_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1139_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_));
AND2X2 AND2X2_4381 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1144_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1141_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_));
AND2X2 AND2X2_4382 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1148_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1146_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_));
AND2X2 AND2X2_4383 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1151_));
AND2X2 AND2X2_4384 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1152_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1150_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_));
AND2X2 AND2X2_4385 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1155_));
AND2X2 AND2X2_4386 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1156_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1154_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_));
AND2X2 AND2X2_4387 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1159_));
AND2X2 AND2X2_4388 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1160_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1158_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_));
AND2X2 AND2X2_4389 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1163_));
AND2X2 AND2X2_439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3153_), .B(AES_CORE_DATAPATH__abc_16009_new_n3137_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__17_));
AND2X2 AND2X2_4390 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1164_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1162_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_));
AND2X2 AND2X2_4391 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1167_));
AND2X2 AND2X2_4392 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1168_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1166_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_));
AND2X2 AND2X2_4393 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1171_));
AND2X2 AND2X2_4394 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1172_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1170_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_));
AND2X2 AND2X2_4395 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1175_));
AND2X2 AND2X2_4396 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1176_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1174_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_));
AND2X2 AND2X2_4397 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1179_));
AND2X2 AND2X2_4398 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1180_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1178_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_));
AND2X2 AND2X2_4399 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1183_));
AND2X2 AND2X2_44 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_));
AND2X2 AND2X2_440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3159_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3160_));
AND2X2 AND2X2_4400 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1184_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1182_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_));
AND2X2 AND2X2_4401 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1187_));
AND2X2 AND2X2_4402 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1188_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1186_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_));
AND2X2 AND2X2_4403 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1191_));
AND2X2 AND2X2_4404 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1192_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1190_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_));
AND2X2 AND2X2_4405 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1195_));
AND2X2 AND2X2_4406 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1196_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1194_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_));
AND2X2 AND2X2_4407 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1199_));
AND2X2 AND2X2_4408 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1200_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1198_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_));
AND2X2 AND2X2_4409 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1203_));
AND2X2 AND2X2_441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3162_));
AND2X2 AND2X2_4410 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1204_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1202_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_));
AND2X2 AND2X2_4411 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1207_));
AND2X2 AND2X2_4412 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1208_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1206_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_));
AND2X2 AND2X2_4413 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1211_));
AND2X2 AND2X2_4414 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1212_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1210_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_));
AND2X2 AND2X2_4415 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1215_));
AND2X2 AND2X2_4416 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1216_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1214_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_));
AND2X2 AND2X2_4417 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1219_));
AND2X2 AND2X2_4418 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1220_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1218_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_));
AND2X2 AND2X2_4419 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1223_));
AND2X2 AND2X2_442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3163_));
AND2X2 AND2X2_4420 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1224_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1222_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_));
AND2X2 AND2X2_4421 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1227_));
AND2X2 AND2X2_4422 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1228_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1226_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_));
AND2X2 AND2X2_4423 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1231_));
AND2X2 AND2X2_4424 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1232_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1230_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_));
AND2X2 AND2X2_4425 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1235_));
AND2X2 AND2X2_4426 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1236_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1234_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_));
AND2X2 AND2X2_4427 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1239_));
AND2X2 AND2X2_4428 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1240_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1238_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_));
AND2X2 AND2X2_4429 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1243_));
AND2X2 AND2X2_443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3165_), .B(AES_CORE_DATAPATH__abc_16009_new_n3157_), .Y(\key_out[18] ));
AND2X2 AND2X2_4430 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1244_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1242_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_));
AND2X2 AND2X2_4431 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1247_));
AND2X2 AND2X2_4432 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1248_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1246_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_));
AND2X2 AND2X2_4433 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1251_));
AND2X2 AND2X2_4434 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1252_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1250_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_));
AND2X2 AND2X2_4435 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1255_));
AND2X2 AND2X2_4436 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1256_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1254_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_));
AND2X2 AND2X2_4437 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1259_));
AND2X2 AND2X2_4438 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1260_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1258_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_));
AND2X2 AND2X2_4439 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1263_));
AND2X2 AND2X2_444 ( .A(\key_out[18] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3156_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3167_));
AND2X2 AND2X2_4440 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1264_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1262_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_));
AND2X2 AND2X2_4441 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1267_));
AND2X2 AND2X2_4442 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1268_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1266_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_));
AND2X2 AND2X2_4443 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1271_));
AND2X2 AND2X2_4444 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1272_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1270_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_));
AND2X2 AND2X2_4445 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1275_));
AND2X2 AND2X2_4446 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1276_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1274_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_));
AND2X2 AND2X2_4447 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n97_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n98_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n99_));
AND2X2 AND2X2_4448 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n100_));
AND2X2 AND2X2_4449 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n103_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n105_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n106_));
AND2X2 AND2X2_445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3168_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3169_));
AND2X2 AND2X2_4450 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n108_));
AND2X2 AND2X2_4451 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n106_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n109_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n110_));
AND2X2 AND2X2_4452 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n114_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n113_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n115_));
AND2X2 AND2X2_4453 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n117_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n112_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_));
AND2X2 AND2X2_4454 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n120_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n121_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n122_));
AND2X2 AND2X2_4455 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n123_));
AND2X2 AND2X2_4456 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n126_));
AND2X2 AND2X2_4457 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n127_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n125_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n128_));
AND2X2 AND2X2_4458 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n130_));
AND2X2 AND2X2_4459 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n131_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n129_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_));
AND2X2 AND2X2_446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3171_), .B(AES_CORE_DATAPATH__abc_16009_new_n3155_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__18_));
AND2X2 AND2X2_4460 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n134_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n136_));
AND2X2 AND2X2_4461 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n138_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n139_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n140_));
AND2X2 AND2X2_4462 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n142_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n133_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_));
AND2X2 AND2X2_4463 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n146_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n145_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_));
AND2X2 AND2X2_4464 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n137_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n148_));
AND2X2 AND2X2_4465 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n128_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n149_));
AND2X2 AND2X2_4466 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n144_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n151_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_));
AND2X2 AND2X2_4467 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n154_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n155_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_));
AND2X2 AND2X2_4468 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n153_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n157_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_));
AND2X2 AND2X2_4469 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n159_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n161_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n162_));
AND2X2 AND2X2_447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3177_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3178_));
AND2X2 AND2X2_4470 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n162_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n163_));
AND2X2 AND2X2_4471 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n164_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n165_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n166_));
AND2X2 AND2X2_4472 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n169_));
AND2X2 AND2X2_4473 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n170_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n168_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n171_));
AND2X2 AND2X2_4474 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n171_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n172_));
AND2X2 AND2X2_4475 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n174_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n176_));
AND2X2 AND2X2_4476 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n177_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n173_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n178_));
AND2X2 AND2X2_4477 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n167_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n180_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n181_));
AND2X2 AND2X2_4478 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n166_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n179_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n182_));
AND2X2 AND2X2_4479 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n186_));
AND2X2 AND2X2_448 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3180_));
AND2X2 AND2X2_4480 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n187_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n185_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_));
AND2X2 AND2X2_4481 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n189_));
AND2X2 AND2X2_4482 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n104_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n191_));
AND2X2 AND2X2_4483 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n193_));
AND2X2 AND2X2_4484 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n196_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n197_));
AND2X2 AND2X2_4485 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n198_));
AND2X2 AND2X2_4486 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n202_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n201_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_));
AND2X2 AND2X2_4487 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n200_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n204_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n205_));
AND2X2 AND2X2_4488 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n207_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n208_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_));
AND2X2 AND2X2_4489 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n210_));
AND2X2 AND2X2_449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3181_));
AND2X2 AND2X2_4490 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n211_));
AND2X2 AND2X2_4491 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n213_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n206_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n214_));
AND2X2 AND2X2_4492 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n216_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n217_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n218_));
AND2X2 AND2X2_4493 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n215_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n219_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_));
AND2X2 AND2X2_4494 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n221_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n223_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n224_));
AND2X2 AND2X2_4495 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n224_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n225_));
AND2X2 AND2X2_4496 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n226_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n227_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n228_));
AND2X2 AND2X2_4497 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n231_));
AND2X2 AND2X2_4498 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n232_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n233_));
AND2X2 AND2X2_4499 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n229_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n235_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n236_));
AND2X2 AND2X2_45 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n91_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n142_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_));
AND2X2 AND2X2_450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3183_), .B(AES_CORE_DATAPATH__abc_16009_new_n3175_), .Y(\key_out[19] ));
AND2X2 AND2X2_4500 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n228_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n234_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n237_));
AND2X2 AND2X2_4501 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n240_));
AND2X2 AND2X2_4502 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n241_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n239_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n242_));
AND2X2 AND2X2_4503 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n109_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n244_));
AND2X2 AND2X2_4504 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n243_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n246_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n247_));
AND2X2 AND2X2_4505 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n102_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n248_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n249_));
AND2X2 AND2X2_4506 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n250_));
AND2X2 AND2X2_4507 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n252_));
AND2X2 AND2X2_4508 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n254_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n253_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_));
AND2X2 AND2X2_4509 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n256_));
AND2X2 AND2X2_451 ( .A(\key_out[19] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3174_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3185_));
AND2X2 AND2X2_4510 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n257_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n258_));
AND2X2 AND2X2_4511 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n259_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n260_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n261_));
AND2X2 AND2X2_4512 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n261_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n262_));
AND2X2 AND2X2_4513 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n245_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n266_));
AND2X2 AND2X2_4514 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n242_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n267_));
AND2X2 AND2X2_4515 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n265_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n269_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n270_));
AND2X2 AND2X2_4516 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n272_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n274_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_));
AND2X2 AND2X2_4517 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n276_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n278_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n279_));
AND2X2 AND2X2_4518 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n279_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n280_));
AND2X2 AND2X2_4519 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n281_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n282_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n283_));
AND2X2 AND2X2_452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3186_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3187_));
AND2X2 AND2X2_4520 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n286_));
AND2X2 AND2X2_4521 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n287_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n288_));
AND2X2 AND2X2_4522 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n289_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n290_));
AND2X2 AND2X2_4523 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n292_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n291_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n293_));
AND2X2 AND2X2_4524 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n284_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n295_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n296_));
AND2X2 AND2X2_4525 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n283_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n294_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n297_));
AND2X2 AND2X2_4526 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n300_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n301_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n302_));
AND2X2 AND2X2_4527 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n115_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n304_));
AND2X2 AND2X2_4528 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n101_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n305_));
AND2X2 AND2X2_4529 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n307_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n303_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n308_));
AND2X2 AND2X2_453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3189_), .B(AES_CORE_DATAPATH__abc_16009_new_n3173_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__19_));
AND2X2 AND2X2_4530 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n268_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n306_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n310_));
AND2X2 AND2X2_4531 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n247_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n311_));
AND2X2 AND2X2_4532 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n309_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n313_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n314_));
AND2X2 AND2X2_4533 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n316_));
AND2X2 AND2X2_4534 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n317_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n315_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n318_));
AND2X2 AND2X2_4535 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n173_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n222_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n320_));
AND2X2 AND2X2_4536 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n322_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n319_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n323_));
AND2X2 AND2X2_4537 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n326_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n325_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n327_));
AND2X2 AND2X2_4538 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n321_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n328_));
AND2X2 AND2X2_4539 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n318_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n329_));
AND2X2 AND2X2_454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3195_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3196_));
AND2X2 AND2X2_4540 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n324_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n331_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n332_));
AND2X2 AND2X2_4541 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n334_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n335_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n336_));
AND2X2 AND2X2_4542 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n333_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n337_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_));
AND2X2 AND2X2_4543 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n339_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n341_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n342_));
AND2X2 AND2X2_4544 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n342_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n343_));
AND2X2 AND2X2_4545 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n344_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n345_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n346_));
AND2X2 AND2X2_4546 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n349_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n351_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_));
AND2X2 AND2X2_4547 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n353_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n354_));
AND2X2 AND2X2_4548 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n355_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n356_));
AND2X2 AND2X2_4549 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n347_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n358_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n359_));
AND2X2 AND2X2_455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3198_));
AND2X2 AND2X2_4550 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n346_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n357_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n360_));
AND2X2 AND2X2_4551 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n277_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n363_));
AND2X2 AND2X2_4552 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n364_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n365_));
AND2X2 AND2X2_4553 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n369_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n367_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n370_));
AND2X2 AND2X2_4554 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n171_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n371_));
AND2X2 AND2X2_4555 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n177_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n372_));
AND2X2 AND2X2_4556 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n330_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n373_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n374_));
AND2X2 AND2X2_4557 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n375_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n376_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n377_));
AND2X2 AND2X2_4558 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n323_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n377_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n378_));
AND2X2 AND2X2_4559 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n381_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n382_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n383_));
AND2X2 AND2X2_456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3199_));
AND2X2 AND2X2_4560 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n384_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n380_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n385_));
AND2X2 AND2X2_4561 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n388_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n387_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n389_));
AND2X2 AND2X2_4562 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n390_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n391_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n392_));
AND2X2 AND2X2_4563 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n386_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n393_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n394_));
AND2X2 AND2X2_4564 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n396_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n397_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n398_));
AND2X2 AND2X2_4565 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n395_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n399_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_));
AND2X2 AND2X2_4566 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n401_));
AND2X2 AND2X2_4567 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n402_));
AND2X2 AND2X2_4568 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n350_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n405_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n406_));
AND2X2 AND2X2_4569 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n407_));
AND2X2 AND2X2_457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3201_), .B(AES_CORE_DATAPATH__abc_16009_new_n3193_), .Y(\key_out[20] ));
AND2X2 AND2X2_4570 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n404_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n409_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n410_));
AND2X2 AND2X2_4571 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n403_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n408_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n411_));
AND2X2 AND2X2_4572 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n415_));
AND2X2 AND2X2_4573 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n416_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n414_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n417_));
AND2X2 AND2X2_4574 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n418_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n419_));
AND2X2 AND2X2_4575 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n417_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n420_));
AND2X2 AND2X2_4576 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n423_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n422_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n424_));
AND2X2 AND2X2_4577 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n257_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n234_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n426_));
AND2X2 AND2X2_4578 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n261_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n235_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n427_));
AND2X2 AND2X2_4579 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n425_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n429_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n430_));
AND2X2 AND2X2_458 ( .A(\key_out[20] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3192_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3203_));
AND2X2 AND2X2_4580 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n428_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n370_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n433_));
AND2X2 AND2X2_4581 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n389_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n424_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n434_));
AND2X2 AND2X2_4582 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n431_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n436_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n437_));
AND2X2 AND2X2_4583 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n435_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n432_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n439_));
AND2X2 AND2X2_4584 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n430_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n421_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n440_));
AND2X2 AND2X2_4585 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n442_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n438_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_));
AND2X2 AND2X2_4586 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n444_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n445_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n446_));
AND2X2 AND2X2_4587 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n446_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n447_));
AND2X2 AND2X2_4588 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n448_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n449_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n450_));
AND2X2 AND2X2_4589 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n451_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n452_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n453_));
AND2X2 AND2X2_459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3204_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3205_));
AND2X2 AND2X2_4590 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n457_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n454_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_));
AND2X2 AND2X2_4591 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n355_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n405_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n460_));
AND2X2 AND2X2_4592 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n461_));
AND2X2 AND2X2_4593 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n289_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n463_));
AND2X2 AND2X2_4594 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n292_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n464_));
AND2X2 AND2X2_4595 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n467_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n468_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n469_));
AND2X2 AND2X2_4596 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n473_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n470_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n474_));
AND2X2 AND2X2_4597 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n475_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n459_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n476_));
AND2X2 AND2X2_4598 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n474_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n477_));
AND2X2 AND2X2_4599 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n479_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n480_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n481_));
AND2X2 AND2X2_46 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n146_));
AND2X2 AND2X2_460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3207_), .B(AES_CORE_DATAPATH__abc_16009_new_n3191_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__20_));
AND2X2 AND2X2_4600 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n482_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n483_));
AND2X2 AND2X2_4601 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n481_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n484_));
AND2X2 AND2X2_4602 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n488_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n486_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_));
AND2X2 AND2X2_4603 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n353_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n491_));
AND2X2 AND2X2_4604 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n471_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n492_));
AND2X2 AND2X2_4605 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n495_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n496_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n497_));
AND2X2 AND2X2_4606 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n500_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n498_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_));
AND2X2 AND2X2_4607 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n502_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n503_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_));
AND2X2 AND2X2_4608 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n245_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n505_));
AND2X2 AND2X2_4609 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n242_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n98_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n506_));
AND2X2 AND2X2_461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3213_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3214_));
AND2X2 AND2X2_4610 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n509_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n511_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_));
AND2X2 AND2X2_4611 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n514_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n515_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n516_));
AND2X2 AND2X2_4612 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n513_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n517_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n518_));
AND2X2 AND2X2_4613 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n516_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n519_));
AND2X2 AND2X2_4614 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n521_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n522_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n523_));
AND2X2 AND2X2_4615 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n524_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n525_));
AND2X2 AND2X2_4616 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n523_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n526_));
AND2X2 AND2X2_4617 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n321_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n528_));
AND2X2 AND2X2_4618 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n318_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n529_));
AND2X2 AND2X2_4619 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n527_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n531_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n532_));
AND2X2 AND2X2_462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3216_));
AND2X2 AND2X2_4620 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n533_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n534_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n535_));
AND2X2 AND2X2_4621 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n537_));
AND2X2 AND2X2_4622 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n538_));
AND2X2 AND2X2_4623 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n539_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n535_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n540_));
AND2X2 AND2X2_4624 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n541_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n542_));
AND2X2 AND2X2_4625 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n544_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n545_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n546_));
AND2X2 AND2X2_4626 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n368_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n547_));
AND2X2 AND2X2_4627 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n366_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n548_));
AND2X2 AND2X2_4628 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n551_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n553_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_));
AND2X2 AND2X2_4629 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n556_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n557_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n558_));
AND2X2 AND2X2_463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3217_));
AND2X2 AND2X2_4630 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n561_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n559_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_));
AND2X2 AND2X2_4631 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n418_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n563_));
AND2X2 AND2X2_4632 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n417_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n564_));
AND2X2 AND2X2_4633 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n567_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n568_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n569_));
AND2X2 AND2X2_4634 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n570_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n571_));
AND2X2 AND2X2_4635 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n569_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n572_));
AND2X2 AND2X2_4636 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n574_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n566_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n575_));
AND2X2 AND2X2_4637 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n573_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n565_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n576_));
AND2X2 AND2X2_4638 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n373_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n578_));
AND2X2 AND2X2_4639 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n314_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n377_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n579_));
AND2X2 AND2X2_464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3219_), .B(AES_CORE_DATAPATH__abc_16009_new_n3211_), .Y(\key_out[21] ));
AND2X2 AND2X2_4640 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n580_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n581_));
AND2X2 AND2X2_4641 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n583_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n584_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n585_));
AND2X2 AND2X2_4642 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n585_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n582_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n586_));
AND2X2 AND2X2_4643 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n588_));
AND2X2 AND2X2_4644 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n471_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n350_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n589_));
AND2X2 AND2X2_4645 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n592_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n593_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n594_));
AND2X2 AND2X2_4646 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n595_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n596_));
AND2X2 AND2X2_4647 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n594_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n597_));
AND2X2 AND2X2_4648 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n599_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n591_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n600_));
AND2X2 AND2X2_4649 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n598_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n590_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n601_));
AND2X2 AND2X2_465 ( .A(\key_out[21] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3210_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3221_));
AND2X2 AND2X2_4650 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n603_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n604_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n605_));
AND2X2 AND2X2_4651 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n608_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n609_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n610_));
AND2X2 AND2X2_4652 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n606_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n611_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_));
AND2X2 AND2X2_4653 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n613_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n614_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n615_));
AND2X2 AND2X2_4654 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n137_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n616_));
AND2X2 AND2X2_4655 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n128_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n139_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n617_));
AND2X2 AND2X2_4656 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n620_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n622_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_));
AND2X2 AND2X2_4657 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n625_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n626_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n627_));
AND2X2 AND2X2_4658 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n629_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n630_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n631_));
AND2X2 AND2X2_4659 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n628_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n632_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_));
AND2X2 AND2X2_466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3222_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3223_));
AND2X2 AND2X2_4660 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n634_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n635_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n636_));
AND2X2 AND2X2_4661 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n638_));
AND2X2 AND2X2_4662 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n196_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n639_));
AND2X2 AND2X2_4663 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n641_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n637_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n642_));
AND2X2 AND2X2_4664 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n640_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n636_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n643_));
AND2X2 AND2X2_4665 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n647_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n646_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n648_));
AND2X2 AND2X2_4666 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n651_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n649_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_));
AND2X2 AND2X2_4667 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n653_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n654_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n655_));
AND2X2 AND2X2_4668 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n656_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n657_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n658_));
AND2X2 AND2X2_4669 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n660_));
AND2X2 AND2X2_467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3225_), .B(AES_CORE_DATAPATH__abc_16009_new_n3209_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__21_));
AND2X2 AND2X2_4670 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n658_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n104_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n661_));
AND2X2 AND2X2_4671 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n664_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n666_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n667_));
AND2X2 AND2X2_4672 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n669_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n670_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n671_));
AND2X2 AND2X2_4673 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n674_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n672_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_));
AND2X2 AND2X2_4674 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n248_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n676_));
AND2X2 AND2X2_4675 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n677_));
AND2X2 AND2X2_4676 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n115_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n679_));
AND2X2 AND2X2_4677 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n101_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n680_));
AND2X2 AND2X2_4678 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n682_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n678_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n683_));
AND2X2 AND2X2_4679 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n681_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n685_));
AND2X2 AND2X2_468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3232_));
AND2X2 AND2X2_4680 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n687_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n688_));
AND2X2 AND2X2_4681 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n689_));
AND2X2 AND2X2_4682 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n552_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n691_));
AND2X2 AND2X2_4683 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n546_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n692_));
AND2X2 AND2X2_4684 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n97_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n109_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n695_));
AND2X2 AND2X2_4685 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n696_));
AND2X2 AND2X2_4686 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n698_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n699_));
AND2X2 AND2X2_4687 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n697_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n678_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n700_));
AND2X2 AND2X2_4688 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n702_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n694_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n703_));
AND2X2 AND2X2_4689 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n701_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n693_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n704_));
AND2X2 AND2X2_469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3234_));
AND2X2 AND2X2_4690 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n707_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n708_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_));
AND2X2 AND2X2_4691 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n174_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n173_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n710_));
AND2X2 AND2X2_4692 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n711_));
AND2X2 AND2X2_4693 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n570_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n713_));
AND2X2 AND2X2_4694 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n569_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n714_));
AND2X2 AND2X2_4695 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n719_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n716_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_));
AND2X2 AND2X2_4696 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n723_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n722_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_));
AND2X2 AND2X2_4697 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n232_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n364_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n725_));
AND2X2 AND2X2_4698 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n726_));
AND2X2 AND2X2_4699 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n727_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n728_));
AND2X2 AND2X2_47 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_10_));
AND2X2 AND2X2_470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3235_));
AND2X2 AND2X2_4700 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n729_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n678_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n730_));
AND2X2 AND2X2_4701 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n733_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n732_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n734_));
AND2X2 AND2X2_4702 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n731_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n734_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n735_));
AND2X2 AND2X2_4703 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n736_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n737_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_));
AND2X2 AND2X2_4704 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n739_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n741_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_));
AND2X2 AND2X2_4705 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n287_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n291_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n743_));
AND2X2 AND2X2_4706 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n744_));
AND2X2 AND2X2_4707 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n745_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n746_));
AND2X2 AND2X2_4708 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n747_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n748_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n749_));
AND2X2 AND2X2_4709 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n353_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n751_));
AND2X2 AND2X2_471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3237_), .B(AES_CORE_DATAPATH__abc_16009_new_n3229_), .Y(\key_out[22] ));
AND2X2 AND2X2_4710 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n405_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n752_));
AND2X2 AND2X2_4711 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n750_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n754_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n755_));
AND2X2 AND2X2_4712 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n749_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n753_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n756_));
AND2X2 AND2X2_4713 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n759_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n760_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_));
AND2X2 AND2X2_4714 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n348_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n355_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n762_));
AND2X2 AND2X2_4715 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n763_));
AND2X2 AND2X2_4716 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n764_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n765_));
AND2X2 AND2X2_4717 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n766_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n767_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n768_));
AND2X2 AND2X2_4718 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n771_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n769_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n772_));
AND2X2 AND2X2_4719 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n775_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n774_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_));
AND2X2 AND2X2_472 ( .A(\key_out[22] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3228_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3239_));
AND2X2 AND2X2_4720 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n777_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n778_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n779_));
AND2X2 AND2X2_4721 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n780_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n781_));
AND2X2 AND2X2_4722 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n779_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n782_));
AND2X2 AND2X2_4723 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n784_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n481_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n785_));
AND2X2 AND2X2_4724 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n783_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n482_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n786_));
AND2X2 AND2X2_4725 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n475_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n788_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n789_));
AND2X2 AND2X2_4726 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n474_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n790_));
AND2X2 AND2X2_4727 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n121_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n792_));
AND2X2 AND2X2_4728 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n793_));
AND2X2 AND2X2_4729 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n795_));
AND2X2 AND2X2_473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3240_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3241_));
AND2X2 AND2X2_4730 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n106_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n248_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n796_));
AND2X2 AND2X2_4731 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n798_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n794_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n799_));
AND2X2 AND2X2_4732 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n800_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n801_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n802_));
AND2X2 AND2X2_4733 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n805_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n804_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_));
AND2X2 AND2X2_4734 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n698_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n807_));
AND2X2 AND2X2_4735 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n697_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n808_));
AND2X2 AND2X2_4736 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n810_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n658_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n811_));
AND2X2 AND2X2_4737 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n809_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n812_));
AND2X2 AND2X2_4738 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n814_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n517_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n815_));
AND2X2 AND2X2_4739 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n516_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n816_));
AND2X2 AND2X2_474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3243_), .B(AES_CORE_DATAPATH__abc_16009_new_n3227_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__22_));
AND2X2 AND2X2_4740 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n109_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n98_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n818_));
AND2X2 AND2X2_4741 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n819_));
AND2X2 AND2X2_4742 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n820_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n821_));
AND2X2 AND2X2_4743 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n822_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n823_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n824_));
AND2X2 AND2X2_4744 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n827_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n826_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n828_));
AND2X2 AND2X2_4745 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n825_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n828_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n829_));
AND2X2 AND2X2_4746 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n830_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n831_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n832_));
AND2X2 AND2X2_4747 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n834_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n835_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_));
AND2X2 AND2X2_4748 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n173_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n837_));
AND2X2 AND2X2_4749 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n838_));
AND2X2 AND2X2_475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3249_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3250_));
AND2X2 AND2X2_4750 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n839_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n840_));
AND2X2 AND2X2_4751 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n845_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n846_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n847_));
AND2X2 AND2X2_4752 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n560_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n847_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n849_));
AND2X2 AND2X2_4753 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n558_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n850_));
AND2X2 AND2X2_4754 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n364_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n852_));
AND2X2 AND2X2_4755 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n853_));
AND2X2 AND2X2_4756 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n854_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n855_));
AND2X2 AND2X2_4757 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n856_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n857_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n858_));
AND2X2 AND2X2_4758 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n418_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n860_));
AND2X2 AND2X2_4759 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n417_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n287_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n861_));
AND2X2 AND2X2_476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3252_));
AND2X2 AND2X2_4760 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n859_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n863_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n864_));
AND2X2 AND2X2_4761 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n858_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n862_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n865_));
AND2X2 AND2X2_4762 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n869_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n867_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_));
AND2X2 AND2X2_4763 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n471_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n871_));
AND2X2 AND2X2_4764 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n348_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n872_));
AND2X2 AND2X2_4765 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n291_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n875_));
AND2X2 AND2X2_4766 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n876_));
AND2X2 AND2X2_4767 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n877_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n878_));
AND2X2 AND2X2_4768 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n879_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n880_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n881_));
AND2X2 AND2X2_4769 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n882_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n874_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n883_));
AND2X2 AND2X2_477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3253_));
AND2X2 AND2X2_4770 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n881_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n873_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n884_));
AND2X2 AND2X2_4771 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n887_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n888_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_));
AND2X2 AND2X2_4772 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n355_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n350_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n890_));
AND2X2 AND2X2_4773 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n891_));
AND2X2 AND2X2_4774 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n637_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n894_));
AND2X2 AND2X2_4775 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n636_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n895_));
AND2X2 AND2X2_4776 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n899_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n897_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n900_));
AND2X2 AND2X2_4777 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n902_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n903_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_));
AND2X2 AND2X2_4778 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n139_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n905_));
AND2X2 AND2X2_4779 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n906_));
AND2X2 AND2X2_478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3255_), .B(AES_CORE_DATAPATH__abc_16009_new_n3247_), .Y(\key_out[23] ));
AND2X2 AND2X2_4780 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n907_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n908_));
AND2X2 AND2X2_4781 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n909_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n910_));
AND2X2 AND2X2_4782 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n913_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n914_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_));
AND2X2 AND2X2_4783 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n918_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n917_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_));
AND2X2 AND2X2_4784 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n920_));
AND2X2 AND2X2_4785 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n921_));
AND2X2 AND2X2_4786 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n924_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n925_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n926_));
AND2X2 AND2X2_4787 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n673_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n926_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n928_));
AND2X2 AND2X2_4788 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n671_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n929_));
AND2X2 AND2X2_4789 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n54_));
AND2X2 AND2X2_479 ( .A(\key_out[23] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3246_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3257_));
AND2X2 AND2X2_4790 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n59_));
AND2X2 AND2X2_4791 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n61_));
AND2X2 AND2X2_4792 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n63_));
AND2X2 AND2X2_4793 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n64_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n65_));
AND2X2 AND2X2_4794 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n68_));
AND2X2 AND2X2_4795 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n69_));
AND2X2 AND2X2_4796 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n71_));
AND2X2 AND2X2_4797 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n74_));
AND2X2 AND2X2_4798 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n76_));
AND2X2 AND2X2_4799 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n81_));
AND2X2 AND2X2_48 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n152_));
AND2X2 AND2X2_480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3258_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3259_));
AND2X2 AND2X2_4800 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n83_));
AND2X2 AND2X2_4801 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n84_));
AND2X2 AND2X2_4802 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n85_));
AND2X2 AND2X2_4803 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n87_));
AND2X2 AND2X2_4804 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n90_));
AND2X2 AND2X2_4805 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n91_));
AND2X2 AND2X2_4806 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n95_));
AND2X2 AND2X2_4807 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n98_));
AND2X2 AND2X2_4808 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n97_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n100_));
AND2X2 AND2X2_4809 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n103_));
AND2X2 AND2X2_481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3261_), .B(AES_CORE_DATAPATH__abc_16009_new_n3245_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__23_));
AND2X2 AND2X2_4810 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n104_));
AND2X2 AND2X2_4811 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n106_));
AND2X2 AND2X2_4812 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n107_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n108_));
AND2X2 AND2X2_4813 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n109_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n110_));
AND2X2 AND2X2_4814 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n112_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n113_));
AND2X2 AND2X2_4815 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n115_));
AND2X2 AND2X2_4816 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n117_));
AND2X2 AND2X2_4817 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n118_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n120_));
AND2X2 AND2X2_4818 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n122_));
AND2X2 AND2X2_4819 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n123_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n124_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n125_));
AND2X2 AND2X2_482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3263_));
AND2X2 AND2X2_4820 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n126_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_));
AND2X2 AND2X2_4821 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n130_));
AND2X2 AND2X2_4822 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n131_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n132_));
AND2X2 AND2X2_4823 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n130_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n133_));
AND2X2 AND2X2_4824 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n93_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n135_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n136_));
AND2X2 AND2X2_4825 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n138_));
AND2X2 AND2X2_4826 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n139_));
AND2X2 AND2X2_4827 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n144_));
AND2X2 AND2X2_4828 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n146_));
AND2X2 AND2X2_4829 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n147_));
AND2X2 AND2X2_483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3266_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3267_));
AND2X2 AND2X2_4830 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n149_));
AND2X2 AND2X2_4831 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n150_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n151_));
AND2X2 AND2X2_4832 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n154_));
AND2X2 AND2X2_4833 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n156_));
AND2X2 AND2X2_4834 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n161_));
AND2X2 AND2X2_4835 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n163_));
AND2X2 AND2X2_4836 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n164_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_));
AND2X2 AND2X2_4837 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n167_));
AND2X2 AND2X2_4838 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n168_));
AND2X2 AND2X2_4839 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n170_));
AND2X2 AND2X2_484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3269_));
AND2X2 AND2X2_4840 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n173_));
AND2X2 AND2X2_4841 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n173_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n171_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n174_));
AND2X2 AND2X2_4842 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n175_));
AND2X2 AND2X2_4843 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n177_));
AND2X2 AND2X2_4844 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n179_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n180_));
AND2X2 AND2X2_4845 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n185_));
AND2X2 AND2X2_4846 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n187_));
AND2X2 AND2X2_4847 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n189_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n191_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n192_));
AND2X2 AND2X2_4848 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n193_));
AND2X2 AND2X2_4849 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n194_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n195_));
AND2X2 AND2X2_485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3270_));
AND2X2 AND2X2_4850 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n159_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n196_));
AND2X2 AND2X2_4851 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n197_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n198_));
AND2X2 AND2X2_4852 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n200_));
AND2X2 AND2X2_4853 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n201_));
AND2X2 AND2X2_4854 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n204_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n206_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n207_));
AND2X2 AND2X2_4855 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n208_));
AND2X2 AND2X2_4856 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n209_));
AND2X2 AND2X2_4857 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n210_));
AND2X2 AND2X2_4858 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n211_));
AND2X2 AND2X2_4859 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n213_));
AND2X2 AND2X2_486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3272_), .B(AES_CORE_DATAPATH__abc_16009_new_n3273_), .Y(\key_out[24] ));
AND2X2 AND2X2_4860 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n216_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n215_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n217_));
AND2X2 AND2X2_4861 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n217_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n218_));
AND2X2 AND2X2_4862 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n220_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n222_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n223_));
AND2X2 AND2X2_4863 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n214_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n224_));
AND2X2 AND2X2_4864 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n227_));
AND2X2 AND2X2_4865 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n228_));
AND2X2 AND2X2_4866 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n229_));
AND2X2 AND2X2_4867 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n232_));
AND2X2 AND2X2_4868 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n233_));
AND2X2 AND2X2_4869 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n235_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n236_));
AND2X2 AND2X2_487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3277_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3278_));
AND2X2 AND2X2_4870 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n242_));
AND2X2 AND2X2_4871 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n238_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_));
AND2X2 AND2X2_4872 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n246_));
AND2X2 AND2X2_4873 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n249_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n250_));
AND2X2 AND2X2_4874 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n251_));
AND2X2 AND2X2_4875 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n254_));
AND2X2 AND2X2_4876 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n255_));
AND2X2 AND2X2_4877 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n258_));
AND2X2 AND2X2_4878 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n249_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n260_));
AND2X2 AND2X2_4879 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n261_));
AND2X2 AND2X2_488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3278_), .B(AES_CORE_DATAPATH__abc_16009_new_n3276_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3279_));
AND2X2 AND2X2_4880 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n264_));
AND2X2 AND2X2_4881 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n266_));
AND2X2 AND2X2_4882 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n267_));
AND2X2 AND2X2_4883 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n270_));
AND2X2 AND2X2_4884 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n271_));
AND2X2 AND2X2_4885 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n274_));
AND2X2 AND2X2_4886 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n275_));
AND2X2 AND2X2_4887 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n276_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_));
AND2X2 AND2X2_4888 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n265_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n280_));
AND2X2 AND2X2_4889 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n281_));
AND2X2 AND2X2_489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3284_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3285_));
AND2X2 AND2X2_4890 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n284_));
AND2X2 AND2X2_4891 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n285_));
AND2X2 AND2X2_4892 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n286_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n288_));
AND2X2 AND2X2_4893 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n289_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n291_));
AND2X2 AND2X2_4894 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n292_));
AND2X2 AND2X2_4895 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n279_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n295_));
AND2X2 AND2X2_4896 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n293_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n296_));
AND2X2 AND2X2_4897 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n298_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_));
AND2X2 AND2X2_4898 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n302_));
AND2X2 AND2X2_4899 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n303_));
AND2X2 AND2X2_49 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT_state_12_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n153_));
AND2X2 AND2X2_490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3287_));
AND2X2 AND2X2_4900 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n304_));
AND2X2 AND2X2_4901 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n307_));
AND2X2 AND2X2_4902 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n309_));
AND2X2 AND2X2_4903 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n310_));
AND2X2 AND2X2_4904 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n311_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n313_));
AND2X2 AND2X2_4905 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n314_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n315_));
AND2X2 AND2X2_4906 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n317_));
AND2X2 AND2X2_4907 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n319_));
AND2X2 AND2X2_4908 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n320_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n321_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_));
AND2X2 AND2X2_4909 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n323_));
AND2X2 AND2X2_491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3288_));
AND2X2 AND2X2_4910 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n324_));
AND2X2 AND2X2_4911 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n327_));
AND2X2 AND2X2_4912 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n328_));
AND2X2 AND2X2_4913 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n329_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n331_));
AND2X2 AND2X2_4914 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n334_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n335_));
AND2X2 AND2X2_4915 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n337_));
AND2X2 AND2X2_4916 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n338_));
AND2X2 AND2X2_4917 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n340_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n341_));
AND2X2 AND2X2_4918 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n342_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n345_));
AND2X2 AND2X2_4919 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n346_));
AND2X2 AND2X2_492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3290_), .B(AES_CORE_DATAPATH__abc_16009_new_n3291_), .Y(\key_out[25] ));
AND2X2 AND2X2_4920 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n347_));
AND2X2 AND2X2_4921 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n348_));
AND2X2 AND2X2_4922 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n350_));
AND2X2 AND2X2_4923 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n352_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n353_));
AND2X2 AND2X2_4924 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n354_));
AND2X2 AND2X2_4925 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n355_));
AND2X2 AND2X2_4926 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n356_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n357_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n358_));
AND2X2 AND2X2_4927 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n361_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n363_));
AND2X2 AND2X2_4928 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n363_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n360_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n364_));
AND2X2 AND2X2_4929 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n367_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_));
AND2X2 AND2X2_493 ( .A(\key_out[25] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3282_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3293_));
AND2X2 AND2X2_4930 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n370_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n372_));
AND2X2 AND2X2_4931 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n373_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_));
AND2X2 AND2X2_4932 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n376_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_));
AND2X2 AND2X2_4933 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n380_));
AND2X2 AND2X2_4934 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n381_));
AND2X2 AND2X2_4935 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n383_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n384_));
AND2X2 AND2X2_4936 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n386_));
AND2X2 AND2X2_4937 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n384_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n387_));
AND2X2 AND2X2_4938 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n389_));
AND2X2 AND2X2_4939 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n390_));
AND2X2 AND2X2_494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3295_));
AND2X2 AND2X2_4940 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n391_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n393_));
AND2X2 AND2X2_4941 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n395_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n397_));
AND2X2 AND2X2_4942 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n400_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n399_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n401_));
AND2X2 AND2X2_4943 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n398_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n402_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_));
AND2X2 AND2X2_4944 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n404_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n405_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n406_));
AND2X2 AND2X2_4945 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n409_));
AND2X2 AND2X2_4946 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n410_));
AND2X2 AND2X2_4947 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n408_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_));
AND2X2 AND2X2_4948 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n407_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n414_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_));
AND2X2 AND2X2_4949 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n417_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_));
AND2X2 AND2X2_495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3297_), .B(AES_CORE_DATAPATH__abc_16009_new_n3281_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__25_));
AND2X2 AND2X2_4950 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n421_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n422_));
AND2X2 AND2X2_4951 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n426_));
AND2X2 AND2X2_4952 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_));
AND2X2 AND2X2_4953 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n429_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n430_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_));
AND2X2 AND2X2_4954 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n432_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_));
AND2X2 AND2X2_4955 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n435_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_));
AND2X2 AND2X2_4956 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n438_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n439_));
AND2X2 AND2X2_4957 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n440_));
AND2X2 AND2X2_4958 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n442_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n445_));
AND2X2 AND2X2_4959 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n447_));
AND2X2 AND2X2_496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3302_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3303_));
AND2X2 AND2X2_4960 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n449_));
AND2X2 AND2X2_4961 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n450_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n452_));
AND2X2 AND2X2_4962 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n448_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n454_));
AND2X2 AND2X2_4963 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n455_));
AND2X2 AND2X2_4964 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n456_));
AND2X2 AND2X2_4965 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n458_));
AND2X2 AND2X2_4966 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n461_));
AND2X2 AND2X2_4967 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n462_));
AND2X2 AND2X2_4968 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n465_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n464_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n466_));
AND2X2 AND2X2_4969 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_));
AND2X2 AND2X2_497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3305_));
AND2X2 AND2X2_4970 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n469_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n470_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n471_));
AND2X2 AND2X2_4971 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n473_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n474_));
AND2X2 AND2X2_4972 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n476_));
AND2X2 AND2X2_4973 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n477_));
AND2X2 AND2X2_4974 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n478_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n480_));
AND2X2 AND2X2_4975 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n481_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n482_));
AND2X2 AND2X2_4976 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n483_));
AND2X2 AND2X2_4977 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n486_));
AND2X2 AND2X2_4978 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n487_));
AND2X2 AND2X2_4979 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n488_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n489_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n490_));
AND2X2 AND2X2_498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3306_));
AND2X2 AND2X2_4980 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n492_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n494_));
AND2X2 AND2X2_4981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n495_));
AND2X2 AND2X2_4982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n496_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n498_));
AND2X2 AND2X2_4983 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n500_));
AND2X2 AND2X2_4984 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n501_));
AND2X2 AND2X2_4985 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n504_));
AND2X2 AND2X2_4986 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n507_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n508_));
AND2X2 AND2X2_4987 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n506_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n510_));
AND2X2 AND2X2_4988 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n513_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n514_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n515_));
AND2X2 AND2X2_4989 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n516_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n512_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_));
AND2X2 AND2X2_499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3308_), .B(AES_CORE_DATAPATH__abc_16009_new_n3309_), .Y(\key_out[26] ));
AND2X2 AND2X2_4990 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n518_));
AND2X2 AND2X2_4991 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n520_));
AND2X2 AND2X2_4992 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n523_));
AND2X2 AND2X2_4993 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n524_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n525_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n526_));
AND2X2 AND2X2_4994 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n528_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n529_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n530_));
AND2X2 AND2X2_4995 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n530_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n531_));
AND2X2 AND2X2_4996 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n532_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n533_));
AND2X2 AND2X2_4997 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n537_));
AND2X2 AND2X2_4998 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n538_));
AND2X2 AND2X2_4999 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n539_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n540_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n541_));
AND2X2 AND2X2_5 ( .A(_abc_15574_new_n13_), .B(\addr[1] ), .Y(AES_CORE_DATAPATH_col_en_host_2_));
AND2X2 AND2X2_50 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n154_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_4_));
AND2X2 AND2X2_500 ( .A(\key_out[26] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3300_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3311_));
AND2X2 AND2X2_5000 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n543_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n544_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n545_));
AND2X2 AND2X2_5001 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n547_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n548_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_));
AND2X2 AND2X2_5002 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n550_));
AND2X2 AND2X2_5003 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n551_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n552_));
AND2X2 AND2X2_5004 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n554_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n555_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_));
AND2X2 AND2X2_5005 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n54_));
AND2X2 AND2X2_5006 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n59_));
AND2X2 AND2X2_5007 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n61_));
AND2X2 AND2X2_5008 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n63_));
AND2X2 AND2X2_5009 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n64_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n65_));
AND2X2 AND2X2_501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3312_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3313_));
AND2X2 AND2X2_5010 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n68_));
AND2X2 AND2X2_5011 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n69_));
AND2X2 AND2X2_5012 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n71_));
AND2X2 AND2X2_5013 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n74_));
AND2X2 AND2X2_5014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n76_));
AND2X2 AND2X2_5015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n81_));
AND2X2 AND2X2_5016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n83_));
AND2X2 AND2X2_5017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n84_));
AND2X2 AND2X2_5018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n85_));
AND2X2 AND2X2_5019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n87_));
AND2X2 AND2X2_502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3315_), .B(AES_CORE_DATAPATH__abc_16009_new_n3299_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__26_));
AND2X2 AND2X2_5020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n90_));
AND2X2 AND2X2_5021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n91_));
AND2X2 AND2X2_5022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n95_));
AND2X2 AND2X2_5023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n98_));
AND2X2 AND2X2_5024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n97_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n100_));
AND2X2 AND2X2_5025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n103_));
AND2X2 AND2X2_5026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n104_));
AND2X2 AND2X2_5027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n106_));
AND2X2 AND2X2_5028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n107_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n108_));
AND2X2 AND2X2_5029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n109_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n110_));
AND2X2 AND2X2_503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3320_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3321_));
AND2X2 AND2X2_5030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n112_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n113_));
AND2X2 AND2X2_5031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n115_));
AND2X2 AND2X2_5032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n117_));
AND2X2 AND2X2_5033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n118_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n120_));
AND2X2 AND2X2_5034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n122_));
AND2X2 AND2X2_5035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n123_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n124_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n125_));
AND2X2 AND2X2_5036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n126_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_));
AND2X2 AND2X2_5037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n130_));
AND2X2 AND2X2_5038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n131_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n132_));
AND2X2 AND2X2_5039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n130_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n133_));
AND2X2 AND2X2_504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3323_));
AND2X2 AND2X2_5040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n93_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n135_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n136_));
AND2X2 AND2X2_5041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n138_));
AND2X2 AND2X2_5042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n139_));
AND2X2 AND2X2_5043 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n144_));
AND2X2 AND2X2_5044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n146_));
AND2X2 AND2X2_5045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n147_));
AND2X2 AND2X2_5046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n149_));
AND2X2 AND2X2_5047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n150_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n151_));
AND2X2 AND2X2_5048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n154_));
AND2X2 AND2X2_5049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n156_));
AND2X2 AND2X2_505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3324_));
AND2X2 AND2X2_5050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n161_));
AND2X2 AND2X2_5051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n163_));
AND2X2 AND2X2_5052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n164_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_));
AND2X2 AND2X2_5053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n167_));
AND2X2 AND2X2_5054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n168_));
AND2X2 AND2X2_5055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n170_));
AND2X2 AND2X2_5056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n173_));
AND2X2 AND2X2_5057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n173_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n171_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n174_));
AND2X2 AND2X2_5058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n175_));
AND2X2 AND2X2_5059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n177_));
AND2X2 AND2X2_506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3326_), .B(AES_CORE_DATAPATH__abc_16009_new_n3327_), .Y(\key_out[27] ));
AND2X2 AND2X2_5060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n179_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n180_));
AND2X2 AND2X2_5061 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n185_));
AND2X2 AND2X2_5062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n187_));
AND2X2 AND2X2_5063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n189_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n191_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n192_));
AND2X2 AND2X2_5064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n193_));
AND2X2 AND2X2_5065 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n194_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n195_));
AND2X2 AND2X2_5066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n159_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n196_));
AND2X2 AND2X2_5067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n197_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n198_));
AND2X2 AND2X2_5068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n200_));
AND2X2 AND2X2_5069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n201_));
AND2X2 AND2X2_507 ( .A(\key_out[27] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3318_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3329_));
AND2X2 AND2X2_5070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n204_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n206_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n207_));
AND2X2 AND2X2_5071 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n208_));
AND2X2 AND2X2_5072 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n209_));
AND2X2 AND2X2_5073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n210_));
AND2X2 AND2X2_5074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n211_));
AND2X2 AND2X2_5075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n213_));
AND2X2 AND2X2_5076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n216_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n215_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n217_));
AND2X2 AND2X2_5077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n217_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n218_));
AND2X2 AND2X2_5078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n220_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n222_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n223_));
AND2X2 AND2X2_5079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n214_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n224_));
AND2X2 AND2X2_508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3330_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3331_));
AND2X2 AND2X2_5080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n227_));
AND2X2 AND2X2_5081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n228_));
AND2X2 AND2X2_5082 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n229_));
AND2X2 AND2X2_5083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n232_));
AND2X2 AND2X2_5084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n233_));
AND2X2 AND2X2_5085 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n235_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n236_));
AND2X2 AND2X2_5086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n242_));
AND2X2 AND2X2_5087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n238_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_));
AND2X2 AND2X2_5088 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n246_));
AND2X2 AND2X2_5089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n249_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n250_));
AND2X2 AND2X2_509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3333_), .B(AES_CORE_DATAPATH__abc_16009_new_n3317_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__27_));
AND2X2 AND2X2_5090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n251_));
AND2X2 AND2X2_5091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n254_));
AND2X2 AND2X2_5092 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n255_));
AND2X2 AND2X2_5093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n258_));
AND2X2 AND2X2_5094 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n249_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n260_));
AND2X2 AND2X2_5095 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n261_));
AND2X2 AND2X2_5096 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n264_));
AND2X2 AND2X2_5097 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n266_));
AND2X2 AND2X2_5098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n267_));
AND2X2 AND2X2_5099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n270_));
AND2X2 AND2X2_51 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n156_));
AND2X2 AND2X2_510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3335_));
AND2X2 AND2X2_5100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n271_));
AND2X2 AND2X2_5101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n274_));
AND2X2 AND2X2_5102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n275_));
AND2X2 AND2X2_5103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n276_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_));
AND2X2 AND2X2_5104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n265_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n280_));
AND2X2 AND2X2_5105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n281_));
AND2X2 AND2X2_5106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n284_));
AND2X2 AND2X2_5107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n285_));
AND2X2 AND2X2_5108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n286_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n288_));
AND2X2 AND2X2_5109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n289_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n291_));
AND2X2 AND2X2_511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3338_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3339_));
AND2X2 AND2X2_5110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n292_));
AND2X2 AND2X2_5111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n279_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n295_));
AND2X2 AND2X2_5112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n293_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n296_));
AND2X2 AND2X2_5113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n298_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_));
AND2X2 AND2X2_5114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n302_));
AND2X2 AND2X2_5115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n303_));
AND2X2 AND2X2_5116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n304_));
AND2X2 AND2X2_5117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n307_));
AND2X2 AND2X2_5118 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n309_));
AND2X2 AND2X2_5119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n310_));
AND2X2 AND2X2_512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3341_));
AND2X2 AND2X2_5120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n311_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n313_));
AND2X2 AND2X2_5121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n314_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n315_));
AND2X2 AND2X2_5122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n317_));
AND2X2 AND2X2_5123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n319_));
AND2X2 AND2X2_5124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n320_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n321_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_));
AND2X2 AND2X2_5125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n323_));
AND2X2 AND2X2_5126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n324_));
AND2X2 AND2X2_5127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n327_));
AND2X2 AND2X2_5128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n328_));
AND2X2 AND2X2_5129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n329_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n331_));
AND2X2 AND2X2_513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3342_));
AND2X2 AND2X2_5130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n334_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n335_));
AND2X2 AND2X2_5131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n337_));
AND2X2 AND2X2_5132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n338_));
AND2X2 AND2X2_5133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n340_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n341_));
AND2X2 AND2X2_5134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n342_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n345_));
AND2X2 AND2X2_5135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n346_));
AND2X2 AND2X2_5136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n347_));
AND2X2 AND2X2_5137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n348_));
AND2X2 AND2X2_5138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n350_));
AND2X2 AND2X2_5139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n352_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n353_));
AND2X2 AND2X2_514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3344_), .B(AES_CORE_DATAPATH__abc_16009_new_n3345_), .Y(\key_out[28] ));
AND2X2 AND2X2_5140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n354_));
AND2X2 AND2X2_5141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n355_));
AND2X2 AND2X2_5142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n356_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n357_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n358_));
AND2X2 AND2X2_5143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n361_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n363_));
AND2X2 AND2X2_5144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n363_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n360_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n364_));
AND2X2 AND2X2_5145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n367_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_));
AND2X2 AND2X2_5146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n370_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n372_));
AND2X2 AND2X2_5147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n373_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_));
AND2X2 AND2X2_5148 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n376_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_));
AND2X2 AND2X2_5149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n380_));
AND2X2 AND2X2_515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3349_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3350_));
AND2X2 AND2X2_5150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n381_));
AND2X2 AND2X2_5151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n383_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n384_));
AND2X2 AND2X2_5152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n386_));
AND2X2 AND2X2_5153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n384_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n387_));
AND2X2 AND2X2_5154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n389_));
AND2X2 AND2X2_5155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n390_));
AND2X2 AND2X2_5156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n391_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n393_));
AND2X2 AND2X2_5157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n395_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n397_));
AND2X2 AND2X2_5158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n400_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n399_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n401_));
AND2X2 AND2X2_5159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n398_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n402_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_));
AND2X2 AND2X2_516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3350_), .B(AES_CORE_DATAPATH__abc_16009_new_n3348_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3351_));
AND2X2 AND2X2_5160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n404_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n405_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n406_));
AND2X2 AND2X2_5161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n409_));
AND2X2 AND2X2_5162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n410_));
AND2X2 AND2X2_5163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n408_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_));
AND2X2 AND2X2_5164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n407_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n414_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_));
AND2X2 AND2X2_5165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n417_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_));
AND2X2 AND2X2_5166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n421_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n422_));
AND2X2 AND2X2_5167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n426_));
AND2X2 AND2X2_5168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_));
AND2X2 AND2X2_5169 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n429_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n430_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_));
AND2X2 AND2X2_517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3353_));
AND2X2 AND2X2_5170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n432_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_));
AND2X2 AND2X2_5171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n435_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_));
AND2X2 AND2X2_5172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n438_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n439_));
AND2X2 AND2X2_5173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n440_));
AND2X2 AND2X2_5174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n442_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n445_));
AND2X2 AND2X2_5175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n447_));
AND2X2 AND2X2_5176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n449_));
AND2X2 AND2X2_5177 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n450_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n452_));
AND2X2 AND2X2_5178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n448_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n454_));
AND2X2 AND2X2_5179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n455_));
AND2X2 AND2X2_518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3356_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3357_));
AND2X2 AND2X2_5180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n456_));
AND2X2 AND2X2_5181 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n458_));
AND2X2 AND2X2_5182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n461_));
AND2X2 AND2X2_5183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n462_));
AND2X2 AND2X2_5184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n465_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n464_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n466_));
AND2X2 AND2X2_5185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_));
AND2X2 AND2X2_5186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n469_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n470_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n471_));
AND2X2 AND2X2_5187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n473_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n474_));
AND2X2 AND2X2_5188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n476_));
AND2X2 AND2X2_5189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n477_));
AND2X2 AND2X2_519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3359_));
AND2X2 AND2X2_5190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n478_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n480_));
AND2X2 AND2X2_5191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n481_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n482_));
AND2X2 AND2X2_5192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n483_));
AND2X2 AND2X2_5193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n486_));
AND2X2 AND2X2_5194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n487_));
AND2X2 AND2X2_5195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n488_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n489_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n490_));
AND2X2 AND2X2_5196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n492_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n494_));
AND2X2 AND2X2_5197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n495_));
AND2X2 AND2X2_5198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n496_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n498_));
AND2X2 AND2X2_5199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n500_));
AND2X2 AND2X2_52 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n157_));
AND2X2 AND2X2_520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3360_));
AND2X2 AND2X2_5200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n501_));
AND2X2 AND2X2_5201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n504_));
AND2X2 AND2X2_5202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n507_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n508_));
AND2X2 AND2X2_5203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n506_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n510_));
AND2X2 AND2X2_5204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n513_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n514_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n515_));
AND2X2 AND2X2_5205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n516_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n512_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_));
AND2X2 AND2X2_5206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n518_));
AND2X2 AND2X2_5207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n520_));
AND2X2 AND2X2_5208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n523_));
AND2X2 AND2X2_5209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n524_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n525_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n526_));
AND2X2 AND2X2_521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3362_), .B(AES_CORE_DATAPATH__abc_16009_new_n3363_), .Y(\key_out[29] ));
AND2X2 AND2X2_5210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n528_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n529_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n530_));
AND2X2 AND2X2_5211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n530_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n531_));
AND2X2 AND2X2_5212 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n532_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n533_));
AND2X2 AND2X2_5213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n537_));
AND2X2 AND2X2_5214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n538_));
AND2X2 AND2X2_5215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n539_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n540_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n541_));
AND2X2 AND2X2_5216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n543_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n544_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n545_));
AND2X2 AND2X2_5217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n547_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n548_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_));
AND2X2 AND2X2_5218 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n550_));
AND2X2 AND2X2_5219 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n551_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n552_));
AND2X2 AND2X2_522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3367_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3368_));
AND2X2 AND2X2_5220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n554_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n555_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_));
AND2X2 AND2X2_5221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n54_));
AND2X2 AND2X2_5222 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n59_));
AND2X2 AND2X2_5223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n61_));
AND2X2 AND2X2_5224 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n63_));
AND2X2 AND2X2_5225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n64_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n65_));
AND2X2 AND2X2_5226 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n68_));
AND2X2 AND2X2_5227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n69_));
AND2X2 AND2X2_5228 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n71_));
AND2X2 AND2X2_5229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n74_));
AND2X2 AND2X2_523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3368_), .B(AES_CORE_DATAPATH__abc_16009_new_n3366_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3369_));
AND2X2 AND2X2_5230 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n76_));
AND2X2 AND2X2_5231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n81_));
AND2X2 AND2X2_5232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n83_));
AND2X2 AND2X2_5233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n84_));
AND2X2 AND2X2_5234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n85_));
AND2X2 AND2X2_5235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n87_));
AND2X2 AND2X2_5236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n90_));
AND2X2 AND2X2_5237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n91_));
AND2X2 AND2X2_5238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n95_));
AND2X2 AND2X2_5239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n98_));
AND2X2 AND2X2_524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3371_));
AND2X2 AND2X2_5240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n97_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n100_));
AND2X2 AND2X2_5241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n103_));
AND2X2 AND2X2_5242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n104_));
AND2X2 AND2X2_5243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n106_));
AND2X2 AND2X2_5244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n107_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n108_));
AND2X2 AND2X2_5245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n109_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n110_));
AND2X2 AND2X2_5246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n112_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n113_));
AND2X2 AND2X2_5247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n115_));
AND2X2 AND2X2_5248 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n117_));
AND2X2 AND2X2_5249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n118_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n120_));
AND2X2 AND2X2_525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3374_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3375_));
AND2X2 AND2X2_5250 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n122_));
AND2X2 AND2X2_5251 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n123_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n124_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n125_));
AND2X2 AND2X2_5252 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n126_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_));
AND2X2 AND2X2_5253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n130_));
AND2X2 AND2X2_5254 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n131_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n132_));
AND2X2 AND2X2_5255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n130_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n133_));
AND2X2 AND2X2_5256 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n93_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n135_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n136_));
AND2X2 AND2X2_5257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n138_));
AND2X2 AND2X2_5258 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n139_));
AND2X2 AND2X2_5259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n144_));
AND2X2 AND2X2_526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3377_));
AND2X2 AND2X2_5260 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n146_));
AND2X2 AND2X2_5261 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n147_));
AND2X2 AND2X2_5262 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n149_));
AND2X2 AND2X2_5263 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n150_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n151_));
AND2X2 AND2X2_5264 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n154_));
AND2X2 AND2X2_5265 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n156_));
AND2X2 AND2X2_5266 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n161_));
AND2X2 AND2X2_5267 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n163_));
AND2X2 AND2X2_5268 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n164_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_));
AND2X2 AND2X2_5269 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n167_));
AND2X2 AND2X2_527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3378_));
AND2X2 AND2X2_5270 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n168_));
AND2X2 AND2X2_5271 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n170_));
AND2X2 AND2X2_5272 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n173_));
AND2X2 AND2X2_5273 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n173_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n171_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n174_));
AND2X2 AND2X2_5274 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n175_));
AND2X2 AND2X2_5275 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n177_));
AND2X2 AND2X2_5276 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n179_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n180_));
AND2X2 AND2X2_5277 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n185_));
AND2X2 AND2X2_5278 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n187_));
AND2X2 AND2X2_5279 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n189_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n191_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n192_));
AND2X2 AND2X2_528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3380_), .B(AES_CORE_DATAPATH__abc_16009_new_n3381_), .Y(\key_out[30] ));
AND2X2 AND2X2_5280 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n193_));
AND2X2 AND2X2_5281 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n194_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n195_));
AND2X2 AND2X2_5282 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n159_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n196_));
AND2X2 AND2X2_5283 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n197_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n198_));
AND2X2 AND2X2_5284 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n200_));
AND2X2 AND2X2_5285 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n201_));
AND2X2 AND2X2_5286 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n204_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n206_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n207_));
AND2X2 AND2X2_5287 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n208_));
AND2X2 AND2X2_5288 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n209_));
AND2X2 AND2X2_5289 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n210_));
AND2X2 AND2X2_529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3385_), .B(AES_CORE_DATAPATH__abc_16009_new_n2803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3386_));
AND2X2 AND2X2_5290 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n211_));
AND2X2 AND2X2_5291 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n213_));
AND2X2 AND2X2_5292 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n216_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n215_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n217_));
AND2X2 AND2X2_5293 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n217_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n218_));
AND2X2 AND2X2_5294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n220_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n222_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n223_));
AND2X2 AND2X2_5295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n214_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n224_));
AND2X2 AND2X2_5296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n227_));
AND2X2 AND2X2_5297 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n228_));
AND2X2 AND2X2_5298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n229_));
AND2X2 AND2X2_5299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n232_));
AND2X2 AND2X2_53 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n93_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n104_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n159_));
AND2X2 AND2X2_530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3386_), .B(AES_CORE_DATAPATH__abc_16009_new_n3384_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3387_));
AND2X2 AND2X2_5300 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n233_));
AND2X2 AND2X2_5301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n235_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n236_));
AND2X2 AND2X2_5302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n242_));
AND2X2 AND2X2_5303 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n238_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_));
AND2X2 AND2X2_5304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n246_));
AND2X2 AND2X2_5305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n249_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n250_));
AND2X2 AND2X2_5306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n251_));
AND2X2 AND2X2_5307 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n254_));
AND2X2 AND2X2_5308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n255_));
AND2X2 AND2X2_5309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n258_));
AND2X2 AND2X2_531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH__abc_16009_new_n3393_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3394_));
AND2X2 AND2X2_5310 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n249_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n260_));
AND2X2 AND2X2_5311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n261_));
AND2X2 AND2X2_5312 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n264_));
AND2X2 AND2X2_5313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n266_));
AND2X2 AND2X2_5314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n267_));
AND2X2 AND2X2_5315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n270_));
AND2X2 AND2X2_5316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n271_));
AND2X2 AND2X2_5317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n274_));
AND2X2 AND2X2_5318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n275_));
AND2X2 AND2X2_5319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n276_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_));
AND2X2 AND2X2_532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2828_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3396_));
AND2X2 AND2X2_5320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n265_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n280_));
AND2X2 AND2X2_5321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n281_));
AND2X2 AND2X2_5322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n284_));
AND2X2 AND2X2_5323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n285_));
AND2X2 AND2X2_5324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n286_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n288_));
AND2X2 AND2X2_5325 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n289_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n291_));
AND2X2 AND2X2_5326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n292_));
AND2X2 AND2X2_5327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n279_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n295_));
AND2X2 AND2X2_5328 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n293_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n296_));
AND2X2 AND2X2_5329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n298_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_));
AND2X2 AND2X2_533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2838_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3397_));
AND2X2 AND2X2_5330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n302_));
AND2X2 AND2X2_5331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n303_));
AND2X2 AND2X2_5332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n304_));
AND2X2 AND2X2_5333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n307_));
AND2X2 AND2X2_5334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n309_));
AND2X2 AND2X2_5335 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n310_));
AND2X2 AND2X2_5336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n311_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n313_));
AND2X2 AND2X2_5337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n314_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n315_));
AND2X2 AND2X2_5338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n317_));
AND2X2 AND2X2_5339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n319_));
AND2X2 AND2X2_534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3399_), .B(AES_CORE_DATAPATH__abc_16009_new_n3391_), .Y(\key_out[31] ));
AND2X2 AND2X2_5340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n320_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n321_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_));
AND2X2 AND2X2_5341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n323_));
AND2X2 AND2X2_5342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n324_));
AND2X2 AND2X2_5343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n327_));
AND2X2 AND2X2_5344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n328_));
AND2X2 AND2X2_5345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n329_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n331_));
AND2X2 AND2X2_5346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n334_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n335_));
AND2X2 AND2X2_5347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n337_));
AND2X2 AND2X2_5348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n338_));
AND2X2 AND2X2_5349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n340_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n341_));
AND2X2 AND2X2_535 ( .A(\key_out[31] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3390_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3401_));
AND2X2 AND2X2_5350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n342_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n345_));
AND2X2 AND2X2_5351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n346_));
AND2X2 AND2X2_5352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n347_));
AND2X2 AND2X2_5353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n348_));
AND2X2 AND2X2_5354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n350_));
AND2X2 AND2X2_5355 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n352_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n353_));
AND2X2 AND2X2_5356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n354_));
AND2X2 AND2X2_5357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n355_));
AND2X2 AND2X2_5358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n356_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n357_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n358_));
AND2X2 AND2X2_5359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n361_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n363_));
AND2X2 AND2X2_536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3402_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3403_));
AND2X2 AND2X2_5360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n363_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n360_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n364_));
AND2X2 AND2X2_5361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n367_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_));
AND2X2 AND2X2_5362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n370_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n372_));
AND2X2 AND2X2_5363 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n373_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_));
AND2X2 AND2X2_5364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n376_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_));
AND2X2 AND2X2_5365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n380_));
AND2X2 AND2X2_5366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n381_));
AND2X2 AND2X2_5367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n383_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n384_));
AND2X2 AND2X2_5368 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n386_));
AND2X2 AND2X2_5369 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n384_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n387_));
AND2X2 AND2X2_537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3405_), .B(AES_CORE_DATAPATH__abc_16009_new_n3389_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__31_));
AND2X2 AND2X2_5370 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n389_));
AND2X2 AND2X2_5371 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n390_));
AND2X2 AND2X2_5372 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n391_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n393_));
AND2X2 AND2X2_5373 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n395_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n397_));
AND2X2 AND2X2_5374 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n400_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n399_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n401_));
AND2X2 AND2X2_5375 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n398_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n402_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_));
AND2X2 AND2X2_5376 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n404_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n405_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n406_));
AND2X2 AND2X2_5377 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n409_));
AND2X2 AND2X2_5378 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n410_));
AND2X2 AND2X2_5379 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n408_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_));
AND2X2 AND2X2_538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_rk_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3407_));
AND2X2 AND2X2_5380 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n407_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n414_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_));
AND2X2 AND2X2_5381 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n417_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_));
AND2X2 AND2X2_5382 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n421_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n422_));
AND2X2 AND2X2_5383 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n426_));
AND2X2 AND2X2_5384 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_));
AND2X2 AND2X2_5385 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n429_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n430_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_));
AND2X2 AND2X2_5386 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n432_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_));
AND2X2 AND2X2_5387 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n435_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_));
AND2X2 AND2X2_5388 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n438_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n439_));
AND2X2 AND2X2_5389 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n440_));
AND2X2 AND2X2_539 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_rk_sel_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3408_));
AND2X2 AND2X2_5390 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n442_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n445_));
AND2X2 AND2X2_5391 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n447_));
AND2X2 AND2X2_5392 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n449_));
AND2X2 AND2X2_5393 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n450_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n452_));
AND2X2 AND2X2_5394 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n448_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n454_));
AND2X2 AND2X2_5395 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n455_));
AND2X2 AND2X2_5396 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n456_));
AND2X2 AND2X2_5397 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n458_));
AND2X2 AND2X2_5398 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n461_));
AND2X2 AND2X2_5399 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n462_));
AND2X2 AND2X2_54 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n142_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_));
AND2X2 AND2X2_540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_rk_sel_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3411_));
AND2X2 AND2X2_5400 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n465_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n464_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n466_));
AND2X2 AND2X2_5401 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_));
AND2X2 AND2X2_5402 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n469_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n470_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n471_));
AND2X2 AND2X2_5403 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n473_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n474_));
AND2X2 AND2X2_5404 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n476_));
AND2X2 AND2X2_5405 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n477_));
AND2X2 AND2X2_5406 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n478_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n480_));
AND2X2 AND2X2_5407 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n481_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n482_));
AND2X2 AND2X2_5408 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n483_));
AND2X2 AND2X2_5409 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n486_));
AND2X2 AND2X2_541 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_rk_sel_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3412_));
AND2X2 AND2X2_5410 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n487_));
AND2X2 AND2X2_5411 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n488_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n489_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n490_));
AND2X2 AND2X2_5412 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n492_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n494_));
AND2X2 AND2X2_5413 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n495_));
AND2X2 AND2X2_5414 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n496_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n498_));
AND2X2 AND2X2_5415 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n500_));
AND2X2 AND2X2_5416 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n501_));
AND2X2 AND2X2_5417 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n504_));
AND2X2 AND2X2_5418 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n507_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n508_));
AND2X2 AND2X2_5419 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n506_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n510_));
AND2X2 AND2X2_542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3410_), .B(AES_CORE_DATAPATH__abc_16009_new_n3414_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3415_));
AND2X2 AND2X2_5420 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n513_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n514_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n515_));
AND2X2 AND2X2_5421 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n516_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n512_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_));
AND2X2 AND2X2_5422 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n518_));
AND2X2 AND2X2_5423 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n520_));
AND2X2 AND2X2_5424 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n523_));
AND2X2 AND2X2_5425 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n524_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n525_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n526_));
AND2X2 AND2X2_5426 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n528_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n529_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n530_));
AND2X2 AND2X2_5427 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n530_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n531_));
AND2X2 AND2X2_5428 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n532_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n533_));
AND2X2 AND2X2_5429 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n537_));
AND2X2 AND2X2_543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3420_), .B(AES_CORE_DATAPATH__abc_16009_new_n3419_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3421_));
AND2X2 AND2X2_5430 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n538_));
AND2X2 AND2X2_5431 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n539_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n540_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n541_));
AND2X2 AND2X2_5432 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n543_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n544_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n545_));
AND2X2 AND2X2_5433 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n547_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n548_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_));
AND2X2 AND2X2_5434 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n550_));
AND2X2 AND2X2_5435 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n551_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n552_));
AND2X2 AND2X2_5436 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n554_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n555_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_));
AND2X2 AND2X2_5437 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n51_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n53_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n54_));
AND2X2 AND2X2_5438 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n56_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n58_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n59_));
AND2X2 AND2X2_5439 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n61_));
AND2X2 AND2X2_544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3421_), .B(AES_CORE_DATAPATH__abc_16009_new_n3418_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3422_));
AND2X2 AND2X2_5440 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n63_));
AND2X2 AND2X2_5441 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n64_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n65_));
AND2X2 AND2X2_5442 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n68_));
AND2X2 AND2X2_5443 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n69_));
AND2X2 AND2X2_5444 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n71_));
AND2X2 AND2X2_5445 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n72_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n74_));
AND2X2 AND2X2_5446 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n76_));
AND2X2 AND2X2_5447 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n78_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n80_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n81_));
AND2X2 AND2X2_5448 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n83_));
AND2X2 AND2X2_5449 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n70_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n84_));
AND2X2 AND2X2_545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3423_));
AND2X2 AND2X2_5450 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n85_));
AND2X2 AND2X2_5451 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n87_));
AND2X2 AND2X2_5452 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n62_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n90_));
AND2X2 AND2X2_5453 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n54_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n55_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n91_));
AND2X2 AND2X2_5454 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n95_));
AND2X2 AND2X2_5455 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n98_));
AND2X2 AND2X2_5456 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n99_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n97_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n100_));
AND2X2 AND2X2_5457 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n60_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n103_));
AND2X2 AND2X2_5458 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n59_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n104_));
AND2X2 AND2X2_5459 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n73_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n106_));
AND2X2 AND2X2_546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3424_), .B(AES_CORE_DATAPATH__abc_16009_new_n3428_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3429_));
AND2X2 AND2X2_5460 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n107_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n108_));
AND2X2 AND2X2_5461 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n109_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n110_));
AND2X2 AND2X2_5462 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n111_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n112_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n113_));
AND2X2 AND2X2_5463 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n115_));
AND2X2 AND2X2_5464 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n117_));
AND2X2 AND2X2_5465 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n118_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n120_));
AND2X2 AND2X2_5466 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n122_));
AND2X2 AND2X2_5467 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n123_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n124_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n125_));
AND2X2 AND2X2_5468 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n121_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n126_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_));
AND2X2 AND2X2_5469 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n128_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n129_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n130_));
AND2X2 AND2X2_547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3421_), .B(AES_CORE_DATAPATH__abc_16009_new_n3417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3430_));
AND2X2 AND2X2_5470 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n131_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n132_));
AND2X2 AND2X2_5471 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n130_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n133_));
AND2X2 AND2X2_5472 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n93_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n135_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n136_));
AND2X2 AND2X2_5473 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n105_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n138_));
AND2X2 AND2X2_5474 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n139_));
AND2X2 AND2X2_5475 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n143_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n142_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n144_));
AND2X2 AND2X2_5476 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n114_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n67_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n146_));
AND2X2 AND2X2_5477 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n113_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n147_));
AND2X2 AND2X2_5478 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n148_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n131_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n149_));
AND2X2 AND2X2_5479 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n150_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n151_));
AND2X2 AND2X2_548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3431_));
AND2X2 AND2X2_5480 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n153_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n145_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n154_));
AND2X2 AND2X2_5481 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n156_));
AND2X2 AND2X2_5482 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n160_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n161_));
AND2X2 AND2X2_5483 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n162_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n163_));
AND2X2 AND2X2_5484 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n164_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n158_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_));
AND2X2 AND2X2_5485 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n167_));
AND2X2 AND2X2_5486 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n168_));
AND2X2 AND2X2_5487 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n170_));
AND2X2 AND2X2_5488 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n158_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n173_));
AND2X2 AND2X2_5489 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n173_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n171_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n174_));
AND2X2 AND2X2_549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3439_));
AND2X2 AND2X2_5490 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n169_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n175_));
AND2X2 AND2X2_5491 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n177_));
AND2X2 AND2X2_5492 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n178_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n179_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n180_));
AND2X2 AND2X2_5493 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n182_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n184_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n185_));
AND2X2 AND2X2_5494 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n187_));
AND2X2 AND2X2_5495 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n189_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n191_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n192_));
AND2X2 AND2X2_5496 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n174_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n193_));
AND2X2 AND2X2_5497 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n194_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n195_));
AND2X2 AND2X2_5498 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n159_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n196_));
AND2X2 AND2X2_5499 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n197_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n160_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n198_));
AND2X2 AND2X2_55 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n161_));
AND2X2 AND2X2_550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3440_), .B(AES_CORE_DATAPATH__abc_16009_new_n3436_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3441_));
AND2X2 AND2X2_5500 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n171_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n200_));
AND2X2 AND2X2_5501 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n200_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n199_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n201_));
AND2X2 AND2X2_5502 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n204_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n206_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n207_));
AND2X2 AND2X2_5503 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n208_));
AND2X2 AND2X2_5504 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n209_));
AND2X2 AND2X2_5505 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n210_));
AND2X2 AND2X2_5506 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n211_));
AND2X2 AND2X2_5507 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n213_));
AND2X2 AND2X2_5508 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n216_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n215_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n217_));
AND2X2 AND2X2_5509 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n217_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n218_));
AND2X2 AND2X2_551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3441_), .B(AES_CORE_DATAPATH__abc_16009_new_n3432_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3442_));
AND2X2 AND2X2_5510 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n220_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n222_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n223_));
AND2X2 AND2X2_5511 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n223_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n214_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n224_));
AND2X2 AND2X2_5512 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n226_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n194_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n227_));
AND2X2 AND2X2_5513 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n188_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n228_));
AND2X2 AND2X2_5514 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n229_));
AND2X2 AND2X2_5515 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n232_));
AND2X2 AND2X2_5516 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n233_));
AND2X2 AND2X2_5517 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n234_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n235_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n236_));
AND2X2 AND2X2_5518 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n241_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n239_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n242_));
AND2X2 AND2X2_5519 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n243_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n238_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_));
AND2X2 AND2X2_552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3442_), .B(AES_CORE_DATAPATH__abc_16009_new_n3429_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3443_));
AND2X2 AND2X2_5520 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n246_));
AND2X2 AND2X2_5521 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n249_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n250_));
AND2X2 AND2X2_5522 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n251_));
AND2X2 AND2X2_5523 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n254_));
AND2X2 AND2X2_5524 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n255_));
AND2X2 AND2X2_5525 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n256_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n257_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n258_));
AND2X2 AND2X2_5526 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n249_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n260_));
AND2X2 AND2X2_5527 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n261_));
AND2X2 AND2X2_5528 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n264_));
AND2X2 AND2X2_5529 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n248_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n265_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n266_));
AND2X2 AND2X2_553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3414_), .B(AES_CORE_DATAPATH__abc_16009_new_n3409_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3445_));
AND2X2 AND2X2_5530 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n267_));
AND2X2 AND2X2_5531 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n270_));
AND2X2 AND2X2_5532 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n271_));
AND2X2 AND2X2_5533 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n272_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n273_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n274_));
AND2X2 AND2X2_5534 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n275_));
AND2X2 AND2X2_5535 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n276_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n277_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_));
AND2X2 AND2X2_5536 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n265_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n259_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n280_));
AND2X2 AND2X2_5537 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n281_));
AND2X2 AND2X2_5538 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n284_));
AND2X2 AND2X2_5539 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n285_));
AND2X2 AND2X2_554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3446_));
AND2X2 AND2X2_5540 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n286_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n287_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n288_));
AND2X2 AND2X2_5541 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n290_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n289_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n291_));
AND2X2 AND2X2_5542 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n292_));
AND2X2 AND2X2_5543 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n294_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n279_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n295_));
AND2X2 AND2X2_5544 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n293_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n296_));
AND2X2 AND2X2_5545 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n300_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n298_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_));
AND2X2 AND2X2_5546 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n302_));
AND2X2 AND2X2_5547 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n186_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n303_));
AND2X2 AND2X2_5548 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n304_));
AND2X2 AND2X2_5549 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n305_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n306_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n307_));
AND2X2 AND2X2_555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3410_), .B(AES_CORE_DATAPATH__abc_16009_new_n3413_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3447_));
AND2X2 AND2X2_5550 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n309_));
AND2X2 AND2X2_5551 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n310_));
AND2X2 AND2X2_5552 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n311_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n312_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n313_));
AND2X2 AND2X2_5553 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n314_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n315_));
AND2X2 AND2X2_5554 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n317_));
AND2X2 AND2X2_5555 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n319_));
AND2X2 AND2X2_5556 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n320_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n321_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_));
AND2X2 AND2X2_5557 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n323_));
AND2X2 AND2X2_5558 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n324_));
AND2X2 AND2X2_5559 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n327_));
AND2X2 AND2X2_556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3448_));
AND2X2 AND2X2_5560 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n328_));
AND2X2 AND2X2_5561 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n329_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n330_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n331_));
AND2X2 AND2X2_5562 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n333_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n334_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n335_));
AND2X2 AND2X2_5563 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n337_));
AND2X2 AND2X2_5564 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n338_));
AND2X2 AND2X2_5565 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n339_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n340_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n341_));
AND2X2 AND2X2_5566 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n342_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n344_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n345_));
AND2X2 AND2X2_5567 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n180_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n263_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n346_));
AND2X2 AND2X2_5568 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n207_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n347_));
AND2X2 AND2X2_5569 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n348_));
AND2X2 AND2X2_557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3444_), .B(AES_CORE_DATAPATH__abc_16009_new_n3450_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3451_));
AND2X2 AND2X2_5570 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n350_));
AND2X2 AND2X2_5571 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n352_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n349_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n353_));
AND2X2 AND2X2_5572 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n354_));
AND2X2 AND2X2_5573 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n355_));
AND2X2 AND2X2_5574 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n356_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n357_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n358_));
AND2X2 AND2X2_5575 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n361_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n362_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n363_));
AND2X2 AND2X2_5576 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n363_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n360_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n364_));
AND2X2 AND2X2_5577 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n359_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n367_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_));
AND2X2 AND2X2_5578 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n370_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n371_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n372_));
AND2X2 AND2X2_5579 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n374_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n373_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_));
AND2X2 AND2X2_558 ( .A(\key_out[0] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3451_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3454_));
AND2X2 AND2X2_5580 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n369_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n376_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_));
AND2X2 AND2X2_5581 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n380_));
AND2X2 AND2X2_5582 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n381_));
AND2X2 AND2X2_5583 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n379_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n383_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n384_));
AND2X2 AND2X2_5584 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n385_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n386_));
AND2X2 AND2X2_5585 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n384_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n387_));
AND2X2 AND2X2_5586 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n389_));
AND2X2 AND2X2_5587 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n390_));
AND2X2 AND2X2_5588 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n391_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n392_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n393_));
AND2X2 AND2X2_5589 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n396_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n395_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n397_));
AND2X2 AND2X2_559 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .B(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH__abc_16009_new_n3459_));
AND2X2 AND2X2_5590 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n400_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n399_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n401_));
AND2X2 AND2X2_5591 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n398_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n402_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_));
AND2X2 AND2X2_5592 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n404_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n405_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n406_));
AND2X2 AND2X2_5593 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n409_));
AND2X2 AND2X2_5594 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n410_));
AND2X2 AND2X2_5595 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n408_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_));
AND2X2 AND2X2_5596 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n407_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n414_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_));
AND2X2 AND2X2_5597 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n417_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n418_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_));
AND2X2 AND2X2_5598 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n420_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n421_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n422_));
AND2X2 AND2X2_5599 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n424_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n425_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n426_));
AND2X2 AND2X2_56 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n111_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n163_));
AND2X2 AND2X2_560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3461_));
AND2X2 AND2X2_5600 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n423_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n427_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_));
AND2X2 AND2X2_5601 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n429_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n430_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_));
AND2X2 AND2X2_5602 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n433_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n432_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_));
AND2X2 AND2X2_5603 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n435_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n436_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_));
AND2X2 AND2X2_5604 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n438_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n439_));
AND2X2 AND2X2_5605 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n440_));
AND2X2 AND2X2_5606 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n444_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n442_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n445_));
AND2X2 AND2X2_5607 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n447_));
AND2X2 AND2X2_5608 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n449_));
AND2X2 AND2X2_5609 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n450_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n451_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n452_));
AND2X2 AND2X2_561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3458_), .B(AES_CORE_DATAPATH__abc_16009_new_n3463_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3464_));
AND2X2 AND2X2_5610 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n448_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n454_));
AND2X2 AND2X2_5611 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n454_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n455_));
AND2X2 AND2X2_5612 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n456_));
AND2X2 AND2X2_5613 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n447_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n458_));
AND2X2 AND2X2_5614 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n461_));
AND2X2 AND2X2_5615 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n446_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n462_));
AND2X2 AND2X2_5616 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n465_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n464_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n466_));
AND2X2 AND2X2_5617 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_));
AND2X2 AND2X2_5618 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n469_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n470_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n471_));
AND2X2 AND2X2_5619 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n473_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n472_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n474_));
AND2X2 AND2X2_562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3464_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3465_));
AND2X2 AND2X2_5620 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n476_));
AND2X2 AND2X2_5621 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n477_));
AND2X2 AND2X2_5622 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n478_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n480_));
AND2X2 AND2X2_5623 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n481_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n460_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n482_));
AND2X2 AND2X2_5624 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n480_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n483_));
AND2X2 AND2X2_5625 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n486_));
AND2X2 AND2X2_5626 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n487_));
AND2X2 AND2X2_5627 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n488_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n489_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n490_));
AND2X2 AND2X2_5628 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n493_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n492_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n494_));
AND2X2 AND2X2_5629 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n485_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n495_));
AND2X2 AND2X2_563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3466_));
AND2X2 AND2X2_5630 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n496_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n497_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n498_));
AND2X2 AND2X2_5631 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n453_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n500_));
AND2X2 AND2X2_5632 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n498_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n501_));
AND2X2 AND2X2_5633 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n445_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n504_));
AND2X2 AND2X2_5634 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n507_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n508_));
AND2X2 AND2X2_5635 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n506_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n510_));
AND2X2 AND2X2_5636 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n513_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n514_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n515_));
AND2X2 AND2X2_5637 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n516_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n512_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_));
AND2X2 AND2X2_5638 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n499_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n503_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n518_));
AND2X2 AND2X2_5639 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n520_));
AND2X2 AND2X2_564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3471_), .B(AES_CORE_DATAPATH__abc_16009_new_n3469_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3472_));
AND2X2 AND2X2_5640 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n523_));
AND2X2 AND2X2_5641 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n524_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n525_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n526_));
AND2X2 AND2X2_5642 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n528_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n529_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n530_));
AND2X2 AND2X2_5643 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n530_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n531_));
AND2X2 AND2X2_5644 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n532_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n509_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n533_));
AND2X2 AND2X2_5645 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n537_));
AND2X2 AND2X2_5646 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n538_));
AND2X2 AND2X2_5647 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n539_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n540_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n541_));
AND2X2 AND2X2_5648 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n543_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n544_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n545_));
AND2X2 AND2X2_5649 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n547_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n548_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_));
AND2X2 AND2X2_565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3473_));
AND2X2 AND2X2_5650 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n550_));
AND2X2 AND2X2_5651 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n551_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n552_));
AND2X2 AND2X2_5652 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n554_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n555_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_));
AND2X2 AND2X2_5653 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n67_), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_));
AND2X2 AND2X2_5654 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n69_));
AND2X2 AND2X2_5655 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n70_), .B(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_));
AND2X2 AND2X2_5656 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n72_));
AND2X2 AND2X2_5657 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n67_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n70_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_));
AND2X2 AND2X2_5658 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n75_));
AND2X2 AND2X2_5659 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_));
AND2X2 AND2X2_566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3474_));
AND2X2 AND2X2_5660 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n77_));
AND2X2 AND2X2_5661 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n80_));
AND2X2 AND2X2_5662 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n81_));
AND2X2 AND2X2_5663 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n83_));
AND2X2 AND2X2_5664 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n84_));
AND2X2 AND2X2_5665 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n87_));
AND2X2 AND2X2_5666 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n88_));
AND2X2 AND2X2_5667 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n90_));
AND2X2 AND2X2_5668 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n91_));
AND2X2 AND2X2_5669 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n94_));
AND2X2 AND2X2_567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3475_));
AND2X2 AND2X2_5670 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n95_));
AND2X2 AND2X2_5671 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n97_));
AND2X2 AND2X2_5672 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n98_));
AND2X2 AND2X2_5673 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n101_));
AND2X2 AND2X2_5674 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n102_));
AND2X2 AND2X2_5675 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n104_));
AND2X2 AND2X2_5676 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n105_));
AND2X2 AND2X2_5677 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n108_));
AND2X2 AND2X2_5678 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n109_));
AND2X2 AND2X2_5679 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n111_));
AND2X2 AND2X2_568 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3478_), .B(AES_CORE_DATAPATH__abc_16009_new_n3472_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3479_));
AND2X2 AND2X2_5680 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n112_));
AND2X2 AND2X2_5681 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n115_));
AND2X2 AND2X2_5682 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n116_));
AND2X2 AND2X2_5683 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n118_));
AND2X2 AND2X2_5684 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n119_));
AND2X2 AND2X2_5685 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n122_));
AND2X2 AND2X2_5686 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n123_));
AND2X2 AND2X2_5687 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n125_));
AND2X2 AND2X2_5688 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n126_));
AND2X2 AND2X2_5689 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n129_));
AND2X2 AND2X2_569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3482_));
AND2X2 AND2X2_5690 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n130_));
AND2X2 AND2X2_5691 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n132_));
AND2X2 AND2X2_5692 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n133_));
AND2X2 AND2X2_5693 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n136_));
AND2X2 AND2X2_5694 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n137_));
AND2X2 AND2X2_5695 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n139_));
AND2X2 AND2X2_5696 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n140_));
AND2X2 AND2X2_5697 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n143_));
AND2X2 AND2X2_5698 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n144_));
AND2X2 AND2X2_5699 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n146_));
AND2X2 AND2X2_57 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n107_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_));
AND2X2 AND2X2_570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3483_));
AND2X2 AND2X2_5700 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n147_));
AND2X2 AND2X2_5701 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n150_));
AND2X2 AND2X2_5702 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n151_));
AND2X2 AND2X2_5703 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n153_));
AND2X2 AND2X2_5704 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n154_));
AND2X2 AND2X2_5705 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n157_));
AND2X2 AND2X2_5706 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n158_));
AND2X2 AND2X2_5707 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n160_));
AND2X2 AND2X2_5708 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n161_));
AND2X2 AND2X2_5709 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n164_));
AND2X2 AND2X2_571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3481_), .B(AES_CORE_DATAPATH__abc_16009_new_n3485_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3486_));
AND2X2 AND2X2_5710 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n165_));
AND2X2 AND2X2_5711 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n167_));
AND2X2 AND2X2_5712 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n168_));
AND2X2 AND2X2_5713 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n171_));
AND2X2 AND2X2_5714 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n172_));
AND2X2 AND2X2_5715 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n174_));
AND2X2 AND2X2_5716 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n175_));
AND2X2 AND2X2_5717 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n178_));
AND2X2 AND2X2_5718 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n179_));
AND2X2 AND2X2_5719 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n181_));
AND2X2 AND2X2_572 ( .A(\key_out[1] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3486_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3489_));
AND2X2 AND2X2_5720 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n182_));
AND2X2 AND2X2_5721 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n185_));
AND2X2 AND2X2_5722 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n186_));
AND2X2 AND2X2_5723 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n188_));
AND2X2 AND2X2_5724 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n189_));
AND2X2 AND2X2_5725 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n192_));
AND2X2 AND2X2_5726 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n193_));
AND2X2 AND2X2_5727 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n195_));
AND2X2 AND2X2_5728 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n196_));
AND2X2 AND2X2_5729 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n199_));
AND2X2 AND2X2_573 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3492_));
AND2X2 AND2X2_5730 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n200_));
AND2X2 AND2X2_5731 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n202_));
AND2X2 AND2X2_5732 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n203_));
AND2X2 AND2X2_5733 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n206_));
AND2X2 AND2X2_5734 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n207_));
AND2X2 AND2X2_5735 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n209_));
AND2X2 AND2X2_5736 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n210_));
AND2X2 AND2X2_5737 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n213_));
AND2X2 AND2X2_5738 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n214_));
AND2X2 AND2X2_5739 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n216_));
AND2X2 AND2X2_574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3493_));
AND2X2 AND2X2_5740 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n217_));
AND2X2 AND2X2_5741 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n220_));
AND2X2 AND2X2_5742 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n221_));
AND2X2 AND2X2_5743 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n223_));
AND2X2 AND2X2_5744 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n224_));
AND2X2 AND2X2_5745 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n227_));
AND2X2 AND2X2_5746 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n228_));
AND2X2 AND2X2_5747 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n230_));
AND2X2 AND2X2_5748 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n231_));
AND2X2 AND2X2_5749 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n234_));
AND2X2 AND2X2_575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3491_), .B(AES_CORE_DATAPATH__abc_16009_new_n3495_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3496_));
AND2X2 AND2X2_5750 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n235_));
AND2X2 AND2X2_5751 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n237_));
AND2X2 AND2X2_5752 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n238_));
AND2X2 AND2X2_5753 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n241_));
AND2X2 AND2X2_5754 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n242_));
AND2X2 AND2X2_5755 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n244_));
AND2X2 AND2X2_5756 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n245_));
AND2X2 AND2X2_5757 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n248_));
AND2X2 AND2X2_5758 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n249_));
AND2X2 AND2X2_5759 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n251_));
AND2X2 AND2X2_576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3496_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3497_));
AND2X2 AND2X2_5760 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n252_));
AND2X2 AND2X2_5761 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n255_));
AND2X2 AND2X2_5762 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n256_));
AND2X2 AND2X2_5763 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n258_));
AND2X2 AND2X2_5764 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n259_));
AND2X2 AND2X2_5765 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n262_));
AND2X2 AND2X2_5766 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n263_));
AND2X2 AND2X2_5767 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n265_));
AND2X2 AND2X2_5768 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n266_));
AND2X2 AND2X2_5769 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n269_));
AND2X2 AND2X2_577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3498_));
AND2X2 AND2X2_5770 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n270_));
AND2X2 AND2X2_5771 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n272_));
AND2X2 AND2X2_5772 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n273_));
AND2X2 AND2X2_5773 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n276_));
AND2X2 AND2X2_5774 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n277_));
AND2X2 AND2X2_5775 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n279_));
AND2X2 AND2X2_5776 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n280_));
AND2X2 AND2X2_5777 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n283_));
AND2X2 AND2X2_5778 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n284_));
AND2X2 AND2X2_5779 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n286_));
AND2X2 AND2X2_578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3503_), .B(AES_CORE_DATAPATH__abc_16009_new_n3501_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3504_));
AND2X2 AND2X2_5780 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n287_));
AND2X2 AND2X2_5781 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n68_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n290_));
AND2X2 AND2X2_5782 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n71_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n291_));
AND2X2 AND2X2_5783 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n74_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n293_));
AND2X2 AND2X2_5784 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n76_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n294_));
AND2X2 AND2X2_5785 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n67_), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_));
AND2X2 AND2X2_5786 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n69_));
AND2X2 AND2X2_5787 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n70_), .B(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_));
AND2X2 AND2X2_5788 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n72_));
AND2X2 AND2X2_5789 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n67_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n70_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_));
AND2X2 AND2X2_579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3505_));
AND2X2 AND2X2_5790 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n75_));
AND2X2 AND2X2_5791 ( .A(\data_type[1] ), .B(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_));
AND2X2 AND2X2_5792 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n77_));
AND2X2 AND2X2_5793 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n80_));
AND2X2 AND2X2_5794 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n81_));
AND2X2 AND2X2_5795 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n83_));
AND2X2 AND2X2_5796 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n84_));
AND2X2 AND2X2_5797 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n87_));
AND2X2 AND2X2_5798 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n88_));
AND2X2 AND2X2_5799 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n90_));
AND2X2 AND2X2_58 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_), .B(\aes_mode[0] ), .Y(AES_CORE_CONTROL_UNIT_mode_cbc));
AND2X2 AND2X2_580 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3506_));
AND2X2 AND2X2_5800 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n91_));
AND2X2 AND2X2_5801 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n94_));
AND2X2 AND2X2_5802 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n95_));
AND2X2 AND2X2_5803 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n97_));
AND2X2 AND2X2_5804 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n98_));
AND2X2 AND2X2_5805 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n101_));
AND2X2 AND2X2_5806 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n102_));
AND2X2 AND2X2_5807 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n104_));
AND2X2 AND2X2_5808 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n105_));
AND2X2 AND2X2_5809 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n108_));
AND2X2 AND2X2_581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3507_));
AND2X2 AND2X2_5810 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n109_));
AND2X2 AND2X2_5811 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n111_));
AND2X2 AND2X2_5812 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n112_));
AND2X2 AND2X2_5813 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n115_));
AND2X2 AND2X2_5814 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n116_));
AND2X2 AND2X2_5815 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n118_));
AND2X2 AND2X2_5816 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n119_));
AND2X2 AND2X2_5817 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n122_));
AND2X2 AND2X2_5818 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n123_));
AND2X2 AND2X2_5819 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n125_));
AND2X2 AND2X2_582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3510_), .B(AES_CORE_DATAPATH__abc_16009_new_n3504_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3511_));
AND2X2 AND2X2_5820 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n126_));
AND2X2 AND2X2_5821 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n129_));
AND2X2 AND2X2_5822 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n130_));
AND2X2 AND2X2_5823 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n132_));
AND2X2 AND2X2_5824 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n133_));
AND2X2 AND2X2_5825 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n136_));
AND2X2 AND2X2_5826 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n137_));
AND2X2 AND2X2_5827 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n139_));
AND2X2 AND2X2_5828 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n140_));
AND2X2 AND2X2_5829 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n143_));
AND2X2 AND2X2_583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3514_));
AND2X2 AND2X2_5830 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n144_));
AND2X2 AND2X2_5831 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n146_));
AND2X2 AND2X2_5832 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n147_));
AND2X2 AND2X2_5833 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n150_));
AND2X2 AND2X2_5834 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n151_));
AND2X2 AND2X2_5835 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n153_));
AND2X2 AND2X2_5836 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n154_));
AND2X2 AND2X2_5837 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n157_));
AND2X2 AND2X2_5838 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n158_));
AND2X2 AND2X2_5839 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n160_));
AND2X2 AND2X2_584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3515_));
AND2X2 AND2X2_5840 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n161_));
AND2X2 AND2X2_5841 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n164_));
AND2X2 AND2X2_5842 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n165_));
AND2X2 AND2X2_5843 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n167_));
AND2X2 AND2X2_5844 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n168_));
AND2X2 AND2X2_5845 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n171_));
AND2X2 AND2X2_5846 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n172_));
AND2X2 AND2X2_5847 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n174_));
AND2X2 AND2X2_5848 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n175_));
AND2X2 AND2X2_5849 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n178_));
AND2X2 AND2X2_585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3513_), .B(AES_CORE_DATAPATH__abc_16009_new_n3517_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3518_));
AND2X2 AND2X2_5850 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n179_));
AND2X2 AND2X2_5851 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n181_));
AND2X2 AND2X2_5852 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n182_));
AND2X2 AND2X2_5853 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n185_));
AND2X2 AND2X2_5854 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n186_));
AND2X2 AND2X2_5855 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n188_));
AND2X2 AND2X2_5856 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n189_));
AND2X2 AND2X2_5857 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n192_));
AND2X2 AND2X2_5858 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n193_));
AND2X2 AND2X2_5859 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n195_));
AND2X2 AND2X2_586 ( .A(\key_out[2] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3518_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3521_));
AND2X2 AND2X2_5860 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n196_));
AND2X2 AND2X2_5861 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n199_));
AND2X2 AND2X2_5862 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n200_));
AND2X2 AND2X2_5863 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n202_));
AND2X2 AND2X2_5864 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n203_));
AND2X2 AND2X2_5865 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n206_));
AND2X2 AND2X2_5866 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n207_));
AND2X2 AND2X2_5867 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n209_));
AND2X2 AND2X2_5868 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n210_));
AND2X2 AND2X2_5869 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n213_));
AND2X2 AND2X2_587 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3524_));
AND2X2 AND2X2_5870 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n214_));
AND2X2 AND2X2_5871 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n216_));
AND2X2 AND2X2_5872 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n217_));
AND2X2 AND2X2_5873 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n220_));
AND2X2 AND2X2_5874 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n221_));
AND2X2 AND2X2_5875 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n223_));
AND2X2 AND2X2_5876 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n224_));
AND2X2 AND2X2_5877 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n227_));
AND2X2 AND2X2_5878 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n228_));
AND2X2 AND2X2_5879 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n230_));
AND2X2 AND2X2_588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3525_));
AND2X2 AND2X2_5880 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n231_));
AND2X2 AND2X2_5881 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n234_));
AND2X2 AND2X2_5882 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n235_));
AND2X2 AND2X2_5883 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n237_));
AND2X2 AND2X2_5884 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n238_));
AND2X2 AND2X2_5885 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n241_));
AND2X2 AND2X2_5886 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n242_));
AND2X2 AND2X2_5887 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n244_));
AND2X2 AND2X2_5888 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n245_));
AND2X2 AND2X2_5889 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n248_));
AND2X2 AND2X2_589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3523_), .B(AES_CORE_DATAPATH__abc_16009_new_n3527_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3528_));
AND2X2 AND2X2_5890 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n249_));
AND2X2 AND2X2_5891 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n251_));
AND2X2 AND2X2_5892 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n252_));
AND2X2 AND2X2_5893 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n255_));
AND2X2 AND2X2_5894 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n256_));
AND2X2 AND2X2_5895 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n258_));
AND2X2 AND2X2_5896 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n259_));
AND2X2 AND2X2_5897 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n262_));
AND2X2 AND2X2_5898 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n263_));
AND2X2 AND2X2_5899 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n265_));
AND2X2 AND2X2_59 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n168_));
AND2X2 AND2X2_590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3528_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3529_));
AND2X2 AND2X2_5900 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n266_));
AND2X2 AND2X2_5901 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n269_));
AND2X2 AND2X2_5902 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n270_));
AND2X2 AND2X2_5903 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n272_));
AND2X2 AND2X2_5904 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n273_));
AND2X2 AND2X2_5905 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n276_));
AND2X2 AND2X2_5906 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n277_));
AND2X2 AND2X2_5907 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n279_));
AND2X2 AND2X2_5908 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n280_));
AND2X2 AND2X2_5909 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n283_));
AND2X2 AND2X2_591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3530_));
AND2X2 AND2X2_5910 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n284_));
AND2X2 AND2X2_5911 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n286_));
AND2X2 AND2X2_5912 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n287_));
AND2X2 AND2X2_5913 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n290_));
AND2X2 AND2X2_5914 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n71_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n291_));
AND2X2 AND2X2_5915 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n293_));
AND2X2 AND2X2_5916 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n294_));
AND2X2 AND2X2_592 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3535_), .B(AES_CORE_DATAPATH__abc_16009_new_n3533_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3536_));
AND2X2 AND2X2_593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3537_));
AND2X2 AND2X2_594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3538_));
AND2X2 AND2X2_595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3539_));
AND2X2 AND2X2_596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3542_), .B(AES_CORE_DATAPATH__abc_16009_new_n3536_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3543_));
AND2X2 AND2X2_597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3546_));
AND2X2 AND2X2_598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3547_));
AND2X2 AND2X2_599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3545_), .B(AES_CORE_DATAPATH__abc_16009_new_n3549_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3550_));
AND2X2 AND2X2_6 ( .A(_abc_15574_new_n15_), .B(\addr[1] ), .Y(AES_CORE_DATAPATH_col_en_host_3_));
AND2X2 AND2X2_60 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n169_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n167_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n170_));
AND2X2 AND2X2_600 ( .A(\key_out[3] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3553_));
AND2X2 AND2X2_601 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3556_));
AND2X2 AND2X2_602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3557_));
AND2X2 AND2X2_603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3555_), .B(AES_CORE_DATAPATH__abc_16009_new_n3559_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3560_));
AND2X2 AND2X2_604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3560_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3561_));
AND2X2 AND2X2_605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3562_));
AND2X2 AND2X2_606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3567_), .B(AES_CORE_DATAPATH__abc_16009_new_n3565_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3568_));
AND2X2 AND2X2_607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3569_));
AND2X2 AND2X2_608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3570_));
AND2X2 AND2X2_609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3571_));
AND2X2 AND2X2_61 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .B(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_));
AND2X2 AND2X2_610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3574_), .B(AES_CORE_DATAPATH__abc_16009_new_n3568_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3575_));
AND2X2 AND2X2_611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3578_));
AND2X2 AND2X2_612 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3579_));
AND2X2 AND2X2_613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3577_), .B(AES_CORE_DATAPATH__abc_16009_new_n3581_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3582_));
AND2X2 AND2X2_614 ( .A(\key_out[4] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3582_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3585_));
AND2X2 AND2X2_615 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3588_));
AND2X2 AND2X2_616 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3589_));
AND2X2 AND2X2_617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3587_), .B(AES_CORE_DATAPATH__abc_16009_new_n3591_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3592_));
AND2X2 AND2X2_618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3592_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3593_));
AND2X2 AND2X2_619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3594_));
AND2X2 AND2X2_62 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n172_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n175_));
AND2X2 AND2X2_620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3599_), .B(AES_CORE_DATAPATH__abc_16009_new_n3597_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3600_));
AND2X2 AND2X2_621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3601_));
AND2X2 AND2X2_622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3602_));
AND2X2 AND2X2_623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3603_));
AND2X2 AND2X2_624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3606_), .B(AES_CORE_DATAPATH__abc_16009_new_n3600_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3607_));
AND2X2 AND2X2_625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3610_));
AND2X2 AND2X2_626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3611_));
AND2X2 AND2X2_627 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3609_), .B(AES_CORE_DATAPATH__abc_16009_new_n3613_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3614_));
AND2X2 AND2X2_628 ( .A(\key_out[5] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3614_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3617_));
AND2X2 AND2X2_629 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3620_));
AND2X2 AND2X2_63 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n170_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n175_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__0_));
AND2X2 AND2X2_630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3621_));
AND2X2 AND2X2_631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3619_), .B(AES_CORE_DATAPATH__abc_16009_new_n3623_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3624_));
AND2X2 AND2X2_632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3624_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3625_));
AND2X2 AND2X2_633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3626_));
AND2X2 AND2X2_634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3631_), .B(AES_CORE_DATAPATH__abc_16009_new_n3629_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3632_));
AND2X2 AND2X2_635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3633_));
AND2X2 AND2X2_636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3634_));
AND2X2 AND2X2_637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3635_));
AND2X2 AND2X2_638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3638_), .B(AES_CORE_DATAPATH__abc_16009_new_n3632_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3639_));
AND2X2 AND2X2_639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3642_));
AND2X2 AND2X2_64 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_), .B(AES_CORE_CONTROL_UNIT_rd_count_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_));
AND2X2 AND2X2_640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3643_));
AND2X2 AND2X2_641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3641_), .B(AES_CORE_DATAPATH__abc_16009_new_n3645_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3646_));
AND2X2 AND2X2_642 ( .A(\key_out[6] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3646_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3649_));
AND2X2 AND2X2_643 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3652_));
AND2X2 AND2X2_644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3653_));
AND2X2 AND2X2_645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3651_), .B(AES_CORE_DATAPATH__abc_16009_new_n3655_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3656_));
AND2X2 AND2X2_646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3656_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3657_));
AND2X2 AND2X2_647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3658_));
AND2X2 AND2X2_648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3663_), .B(AES_CORE_DATAPATH__abc_16009_new_n3661_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3664_));
AND2X2 AND2X2_649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3665_));
AND2X2 AND2X2_65 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n179_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n177_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n180_));
AND2X2 AND2X2_650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3666_));
AND2X2 AND2X2_651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3667_));
AND2X2 AND2X2_652 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3670_), .B(AES_CORE_DATAPATH__abc_16009_new_n3664_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3671_));
AND2X2 AND2X2_653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3674_));
AND2X2 AND2X2_654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3675_));
AND2X2 AND2X2_655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3673_), .B(AES_CORE_DATAPATH__abc_16009_new_n3677_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3678_));
AND2X2 AND2X2_656 ( .A(\key_out[7] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3678_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3681_));
AND2X2 AND2X2_657 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3684_));
AND2X2 AND2X2_658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3685_));
AND2X2 AND2X2_659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3683_), .B(AES_CORE_DATAPATH__abc_16009_new_n3687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3688_));
AND2X2 AND2X2_66 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n180_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n170_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__1_));
AND2X2 AND2X2_660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3688_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3689_));
AND2X2 AND2X2_661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3690_));
AND2X2 AND2X2_662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3695_), .B(AES_CORE_DATAPATH__abc_16009_new_n3693_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3696_));
AND2X2 AND2X2_663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3697_));
AND2X2 AND2X2_664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3698_));
AND2X2 AND2X2_665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3699_));
AND2X2 AND2X2_666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3702_), .B(AES_CORE_DATAPATH__abc_16009_new_n3696_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3703_));
AND2X2 AND2X2_667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3706_));
AND2X2 AND2X2_668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3707_));
AND2X2 AND2X2_669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3705_), .B(AES_CORE_DATAPATH__abc_16009_new_n3709_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3710_));
AND2X2 AND2X2_67 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .B(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n182_));
AND2X2 AND2X2_670 ( .A(\key_out[8] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3710_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3713_));
AND2X2 AND2X2_671 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3716_));
AND2X2 AND2X2_672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3717_));
AND2X2 AND2X2_673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3715_), .B(AES_CORE_DATAPATH__abc_16009_new_n3719_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3720_));
AND2X2 AND2X2_674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3720_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3721_));
AND2X2 AND2X2_675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3722_));
AND2X2 AND2X2_676 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3727_), .B(AES_CORE_DATAPATH__abc_16009_new_n3725_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3728_));
AND2X2 AND2X2_677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3729_));
AND2X2 AND2X2_678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3730_));
AND2X2 AND2X2_679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3731_));
AND2X2 AND2X2_68 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n170_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n184_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n185_));
AND2X2 AND2X2_680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3734_), .B(AES_CORE_DATAPATH__abc_16009_new_n3728_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3735_));
AND2X2 AND2X2_681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3738_));
AND2X2 AND2X2_682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3739_));
AND2X2 AND2X2_683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3737_), .B(AES_CORE_DATAPATH__abc_16009_new_n3741_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3742_));
AND2X2 AND2X2_684 ( .A(\key_out[9] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3742_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3745_));
AND2X2 AND2X2_685 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3748_));
AND2X2 AND2X2_686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3749_));
AND2X2 AND2X2_687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3747_), .B(AES_CORE_DATAPATH__abc_16009_new_n3751_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3752_));
AND2X2 AND2X2_688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3752_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3753_));
AND2X2 AND2X2_689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3754_));
AND2X2 AND2X2_69 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n185_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n183_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__2_));
AND2X2 AND2X2_690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3759_), .B(AES_CORE_DATAPATH__abc_16009_new_n3757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3760_));
AND2X2 AND2X2_691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3761_));
AND2X2 AND2X2_692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3762_));
AND2X2 AND2X2_693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3763_));
AND2X2 AND2X2_694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3766_), .B(AES_CORE_DATAPATH__abc_16009_new_n3760_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3767_));
AND2X2 AND2X2_695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3770_));
AND2X2 AND2X2_696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3771_));
AND2X2 AND2X2_697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3769_), .B(AES_CORE_DATAPATH__abc_16009_new_n3773_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3774_));
AND2X2 AND2X2_698 ( .A(\key_out[10] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3774_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3777_));
AND2X2 AND2X2_699 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3780_));
AND2X2 AND2X2_7 ( .A(\addr[0] ), .B(read_en), .Y(AES_CORE_DATAPATH_col_sel_host_0_));
AND2X2 AND2X2_70 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n183_), .B(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n187_));
AND2X2 AND2X2_700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3781_));
AND2X2 AND2X2_701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3779_), .B(AES_CORE_DATAPATH__abc_16009_new_n3783_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3784_));
AND2X2 AND2X2_702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3784_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3785_));
AND2X2 AND2X2_703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3786_));
AND2X2 AND2X2_704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3791_), .B(AES_CORE_DATAPATH__abc_16009_new_n3789_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3792_));
AND2X2 AND2X2_705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3793_));
AND2X2 AND2X2_706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3794_));
AND2X2 AND2X2_707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3795_));
AND2X2 AND2X2_708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3798_), .B(AES_CORE_DATAPATH__abc_16009_new_n3792_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3799_));
AND2X2 AND2X2_709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3802_));
AND2X2 AND2X2_71 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n182_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n188_));
AND2X2 AND2X2_710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3803_));
AND2X2 AND2X2_711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3801_), .B(AES_CORE_DATAPATH__abc_16009_new_n3805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3806_));
AND2X2 AND2X2_712 ( .A(\key_out[11] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3806_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3809_));
AND2X2 AND2X2_713 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3812_));
AND2X2 AND2X2_714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3813_));
AND2X2 AND2X2_715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3811_), .B(AES_CORE_DATAPATH__abc_16009_new_n3815_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3816_));
AND2X2 AND2X2_716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3816_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3817_));
AND2X2 AND2X2_717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3818_));
AND2X2 AND2X2_718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3823_), .B(AES_CORE_DATAPATH__abc_16009_new_n3821_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3824_));
AND2X2 AND2X2_719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3825_));
AND2X2 AND2X2_72 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n189_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n170_), .Y(AES_CORE_CONTROL_UNIT__0rd_count_3_0__3_));
AND2X2 AND2X2_720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3826_));
AND2X2 AND2X2_721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3827_));
AND2X2 AND2X2_722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3830_), .B(AES_CORE_DATAPATH__abc_16009_new_n3824_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3831_));
AND2X2 AND2X2_723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3834_));
AND2X2 AND2X2_724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3835_));
AND2X2 AND2X2_725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3833_), .B(AES_CORE_DATAPATH__abc_16009_new_n3837_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3838_));
AND2X2 AND2X2_726 ( .A(\key_out[12] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3838_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3841_));
AND2X2 AND2X2_727 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3844_));
AND2X2 AND2X2_728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3845_));
AND2X2 AND2X2_729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3843_), .B(AES_CORE_DATAPATH__abc_16009_new_n3847_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3848_));
AND2X2 AND2X2_73 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n193_), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT_rk_sel_0_));
AND2X2 AND2X2_730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3848_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3849_));
AND2X2 AND2X2_731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3850_));
AND2X2 AND2X2_732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3855_), .B(AES_CORE_DATAPATH__abc_16009_new_n3853_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3856_));
AND2X2 AND2X2_733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3857_));
AND2X2 AND2X2_734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3858_));
AND2X2 AND2X2_735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3859_));
AND2X2 AND2X2_736 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3862_), .B(AES_CORE_DATAPATH__abc_16009_new_n3856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3863_));
AND2X2 AND2X2_737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3866_));
AND2X2 AND2X2_738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3867_));
AND2X2 AND2X2_739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3865_), .B(AES_CORE_DATAPATH__abc_16009_new_n3869_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3870_));
AND2X2 AND2X2_74 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n142_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n193_), .Y(AES_CORE_CONTROL_UNIT_rk_sel_1_));
AND2X2 AND2X2_740 ( .A(\key_out[13] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3870_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3873_));
AND2X2 AND2X2_741 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3876_));
AND2X2 AND2X2_742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3877_));
AND2X2 AND2X2_743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3875_), .B(AES_CORE_DATAPATH__abc_16009_new_n3879_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3880_));
AND2X2 AND2X2_744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3880_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3881_));
AND2X2 AND2X2_745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3882_));
AND2X2 AND2X2_746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3887_), .B(AES_CORE_DATAPATH__abc_16009_new_n3885_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3888_));
AND2X2 AND2X2_747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3889_));
AND2X2 AND2X2_748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3890_));
AND2X2 AND2X2_749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3891_));
AND2X2 AND2X2_75 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n197_));
AND2X2 AND2X2_750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3894_), .B(AES_CORE_DATAPATH__abc_16009_new_n3888_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3895_));
AND2X2 AND2X2_751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3898_));
AND2X2 AND2X2_752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3899_));
AND2X2 AND2X2_753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3897_), .B(AES_CORE_DATAPATH__abc_16009_new_n3901_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3902_));
AND2X2 AND2X2_754 ( .A(\key_out[14] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3902_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3905_));
AND2X2 AND2X2_755 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3908_));
AND2X2 AND2X2_756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3909_));
AND2X2 AND2X2_757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3907_), .B(AES_CORE_DATAPATH__abc_16009_new_n3911_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3912_));
AND2X2 AND2X2_758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3912_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3913_));
AND2X2 AND2X2_759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3914_));
AND2X2 AND2X2_76 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n142_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n199_));
AND2X2 AND2X2_760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3919_), .B(AES_CORE_DATAPATH__abc_16009_new_n3917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3920_));
AND2X2 AND2X2_761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3921_));
AND2X2 AND2X2_762 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3922_));
AND2X2 AND2X2_763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3923_));
AND2X2 AND2X2_764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3926_), .B(AES_CORE_DATAPATH__abc_16009_new_n3920_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3927_));
AND2X2 AND2X2_765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3930_));
AND2X2 AND2X2_766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3931_));
AND2X2 AND2X2_767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3929_), .B(AES_CORE_DATAPATH__abc_16009_new_n3933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3934_));
AND2X2 AND2X2_768 ( .A(\key_out[15] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3934_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3937_));
AND2X2 AND2X2_769 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3940_));
AND2X2 AND2X2_77 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n199_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n200_));
AND2X2 AND2X2_770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3941_));
AND2X2 AND2X2_771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3939_), .B(AES_CORE_DATAPATH__abc_16009_new_n3943_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3944_));
AND2X2 AND2X2_772 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3944_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3945_));
AND2X2 AND2X2_773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3946_));
AND2X2 AND2X2_774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3951_), .B(AES_CORE_DATAPATH__abc_16009_new_n3949_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3952_));
AND2X2 AND2X2_775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3953_));
AND2X2 AND2X2_776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3954_));
AND2X2 AND2X2_777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3955_));
AND2X2 AND2X2_778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3958_), .B(AES_CORE_DATAPATH__abc_16009_new_n3952_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3959_));
AND2X2 AND2X2_779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3962_));
AND2X2 AND2X2_78 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n211_));
AND2X2 AND2X2_780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3963_));
AND2X2 AND2X2_781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3961_), .B(AES_CORE_DATAPATH__abc_16009_new_n3965_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3966_));
AND2X2 AND2X2_782 ( .A(\key_out[16] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3966_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3969_));
AND2X2 AND2X2_783 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3972_));
AND2X2 AND2X2_784 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3973_));
AND2X2 AND2X2_785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3971_), .B(AES_CORE_DATAPATH__abc_16009_new_n3975_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3976_));
AND2X2 AND2X2_786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3976_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n3977_));
AND2X2 AND2X2_787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3978_));
AND2X2 AND2X2_788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3983_), .B(AES_CORE_DATAPATH__abc_16009_new_n3981_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3984_));
AND2X2 AND2X2_789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3985_));
AND2X2 AND2X2_79 ( .A(AES_CORE_CONTROL_UNIT_last_round), .B(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n212_));
AND2X2 AND2X2_790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3986_));
AND2X2 AND2X2_791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3987_));
AND2X2 AND2X2_792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3990_), .B(AES_CORE_DATAPATH__abc_16009_new_n3984_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3991_));
AND2X2 AND2X2_793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3994_));
AND2X2 AND2X2_794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3995_));
AND2X2 AND2X2_795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3993_), .B(AES_CORE_DATAPATH__abc_16009_new_n3997_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3998_));
AND2X2 AND2X2_796 ( .A(\key_out[17] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3998_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4001_));
AND2X2 AND2X2_797 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4004_));
AND2X2 AND2X2_798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4005_));
AND2X2 AND2X2_799 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4003_), .B(AES_CORE_DATAPATH__abc_16009_new_n4007_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4008_));
AND2X2 AND2X2_8 ( .A(\addr[1] ), .B(read_en), .Y(AES_CORE_DATAPATH_col_sel_host_1_));
AND2X2 AND2X2_80 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n212_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n213_));
AND2X2 AND2X2_800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4008_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4009_));
AND2X2 AND2X2_801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4010_));
AND2X2 AND2X2_802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4015_), .B(AES_CORE_DATAPATH__abc_16009_new_n4013_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4016_));
AND2X2 AND2X2_803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4017_));
AND2X2 AND2X2_804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4018_));
AND2X2 AND2X2_805 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4019_));
AND2X2 AND2X2_806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4022_), .B(AES_CORE_DATAPATH__abc_16009_new_n4016_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4023_));
AND2X2 AND2X2_807 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4026_));
AND2X2 AND2X2_808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4027_));
AND2X2 AND2X2_809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4025_), .B(AES_CORE_DATAPATH__abc_16009_new_n4029_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4030_));
AND2X2 AND2X2_81 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n216_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n217_));
AND2X2 AND2X2_810 ( .A(\key_out[18] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4033_));
AND2X2 AND2X2_811 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4036_));
AND2X2 AND2X2_812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4037_));
AND2X2 AND2X2_813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4035_), .B(AES_CORE_DATAPATH__abc_16009_new_n4039_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4040_));
AND2X2 AND2X2_814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4040_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4041_));
AND2X2 AND2X2_815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4042_));
AND2X2 AND2X2_816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4047_), .B(AES_CORE_DATAPATH__abc_16009_new_n4045_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4048_));
AND2X2 AND2X2_817 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4049_));
AND2X2 AND2X2_818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4050_));
AND2X2 AND2X2_819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4051_));
AND2X2 AND2X2_82 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n218_), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n219_));
AND2X2 AND2X2_820 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4054_), .B(AES_CORE_DATAPATH__abc_16009_new_n4048_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4055_));
AND2X2 AND2X2_821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4058_));
AND2X2 AND2X2_822 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4059_));
AND2X2 AND2X2_823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4057_), .B(AES_CORE_DATAPATH__abc_16009_new_n4061_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4062_));
AND2X2 AND2X2_824 ( .A(\key_out[19] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4062_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4065_));
AND2X2 AND2X2_825 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4068_));
AND2X2 AND2X2_826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4069_));
AND2X2 AND2X2_827 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4067_), .B(AES_CORE_DATAPATH__abc_16009_new_n4071_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4072_));
AND2X2 AND2X2_828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4072_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4073_));
AND2X2 AND2X2_829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4074_));
AND2X2 AND2X2_83 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n221_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n215_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n222_));
AND2X2 AND2X2_830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4079_), .B(AES_CORE_DATAPATH__abc_16009_new_n4077_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4080_));
AND2X2 AND2X2_831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4081_));
AND2X2 AND2X2_832 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4082_));
AND2X2 AND2X2_833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4083_));
AND2X2 AND2X2_834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4086_), .B(AES_CORE_DATAPATH__abc_16009_new_n4080_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4087_));
AND2X2 AND2X2_835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4090_));
AND2X2 AND2X2_836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4091_));
AND2X2 AND2X2_837 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4089_), .B(AES_CORE_DATAPATH__abc_16009_new_n4093_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4094_));
AND2X2 AND2X2_838 ( .A(\key_out[20] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4094_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4097_));
AND2X2 AND2X2_839 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4100_));
AND2X2 AND2X2_84 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n223_));
AND2X2 AND2X2_840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4101_));
AND2X2 AND2X2_841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4099_), .B(AES_CORE_DATAPATH__abc_16009_new_n4103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4104_));
AND2X2 AND2X2_842 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4104_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4105_));
AND2X2 AND2X2_843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4106_));
AND2X2 AND2X2_844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4111_), .B(AES_CORE_DATAPATH__abc_16009_new_n4109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4112_));
AND2X2 AND2X2_845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4113_));
AND2X2 AND2X2_846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4114_));
AND2X2 AND2X2_847 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4115_));
AND2X2 AND2X2_848 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4118_), .B(AES_CORE_DATAPATH__abc_16009_new_n4112_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4119_));
AND2X2 AND2X2_849 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4122_));
AND2X2 AND2X2_85 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n214_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n193_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n227_));
AND2X2 AND2X2_850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4123_));
AND2X2 AND2X2_851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4121_), .B(AES_CORE_DATAPATH__abc_16009_new_n4125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4126_));
AND2X2 AND2X2_852 ( .A(\key_out[21] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4129_));
AND2X2 AND2X2_853 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4132_));
AND2X2 AND2X2_854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4133_));
AND2X2 AND2X2_855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4131_), .B(AES_CORE_DATAPATH__abc_16009_new_n4135_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4136_));
AND2X2 AND2X2_856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4136_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4137_));
AND2X2 AND2X2_857 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4138_));
AND2X2 AND2X2_858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4143_), .B(AES_CORE_DATAPATH__abc_16009_new_n4141_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4144_));
AND2X2 AND2X2_859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4145_));
AND2X2 AND2X2_86 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n228_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n229_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n230_));
AND2X2 AND2X2_860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4146_));
AND2X2 AND2X2_861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4147_));
AND2X2 AND2X2_862 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4150_), .B(AES_CORE_DATAPATH__abc_16009_new_n4144_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4151_));
AND2X2 AND2X2_863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4154_));
AND2X2 AND2X2_864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4155_));
AND2X2 AND2X2_865 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4153_), .B(AES_CORE_DATAPATH__abc_16009_new_n4157_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4158_));
AND2X2 AND2X2_866 ( .A(\key_out[22] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4158_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4161_));
AND2X2 AND2X2_867 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4164_));
AND2X2 AND2X2_868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4165_));
AND2X2 AND2X2_869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4163_), .B(AES_CORE_DATAPATH__abc_16009_new_n4167_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4168_));
AND2X2 AND2X2_87 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n231_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n232_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n233_));
AND2X2 AND2X2_870 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4168_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4169_));
AND2X2 AND2X2_871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4170_));
AND2X2 AND2X2_872 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4175_), .B(AES_CORE_DATAPATH__abc_16009_new_n4173_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4176_));
AND2X2 AND2X2_873 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4177_));
AND2X2 AND2X2_874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4178_));
AND2X2 AND2X2_875 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4179_));
AND2X2 AND2X2_876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4182_), .B(AES_CORE_DATAPATH__abc_16009_new_n4176_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4183_));
AND2X2 AND2X2_877 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4186_));
AND2X2 AND2X2_878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4187_));
AND2X2 AND2X2_879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4185_), .B(AES_CORE_DATAPATH__abc_16009_new_n4189_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4190_));
AND2X2 AND2X2_88 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n230_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n233_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n234_));
AND2X2 AND2X2_880 ( .A(\key_out[23] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4190_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4193_));
AND2X2 AND2X2_881 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4196_));
AND2X2 AND2X2_882 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4197_));
AND2X2 AND2X2_883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4195_), .B(AES_CORE_DATAPATH__abc_16009_new_n4199_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4200_));
AND2X2 AND2X2_884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4200_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4201_));
AND2X2 AND2X2_885 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4202_));
AND2X2 AND2X2_886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4207_), .B(AES_CORE_DATAPATH__abc_16009_new_n4205_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4208_));
AND2X2 AND2X2_887 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4209_));
AND2X2 AND2X2_888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4210_));
AND2X2 AND2X2_889 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4211_));
AND2X2 AND2X2_89 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n139_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n238_));
AND2X2 AND2X2_890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4214_), .B(AES_CORE_DATAPATH__abc_16009_new_n4208_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4215_));
AND2X2 AND2X2_891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4218_));
AND2X2 AND2X2_892 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4219_));
AND2X2 AND2X2_893 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4217_), .B(AES_CORE_DATAPATH__abc_16009_new_n4221_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4222_));
AND2X2 AND2X2_894 ( .A(\key_out[24] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4222_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4225_));
AND2X2 AND2X2_895 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4228_));
AND2X2 AND2X2_896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4229_));
AND2X2 AND2X2_897 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4227_), .B(AES_CORE_DATAPATH__abc_16009_new_n4231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4232_));
AND2X2 AND2X2_898 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4232_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4233_));
AND2X2 AND2X2_899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4234_));
AND2X2 AND2X2_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n74_), .B(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_));
AND2X2 AND2X2_90 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n243_));
AND2X2 AND2X2_900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4239_), .B(AES_CORE_DATAPATH__abc_16009_new_n4237_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4240_));
AND2X2 AND2X2_901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4241_));
AND2X2 AND2X2_902 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4242_));
AND2X2 AND2X2_903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4243_));
AND2X2 AND2X2_904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4246_), .B(AES_CORE_DATAPATH__abc_16009_new_n4240_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4247_));
AND2X2 AND2X2_905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4250_));
AND2X2 AND2X2_906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4251_));
AND2X2 AND2X2_907 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4249_), .B(AES_CORE_DATAPATH__abc_16009_new_n4253_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4254_));
AND2X2 AND2X2_908 ( .A(\key_out[25] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4254_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4257_));
AND2X2 AND2X2_909 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4260_));
AND2X2 AND2X2_91 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n244_));
AND2X2 AND2X2_910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4261_));
AND2X2 AND2X2_911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4259_), .B(AES_CORE_DATAPATH__abc_16009_new_n4263_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4264_));
AND2X2 AND2X2_912 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4264_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4265_));
AND2X2 AND2X2_913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4266_));
AND2X2 AND2X2_914 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4271_), .B(AES_CORE_DATAPATH__abc_16009_new_n4269_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4272_));
AND2X2 AND2X2_915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4273_));
AND2X2 AND2X2_916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4274_));
AND2X2 AND2X2_917 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4275_));
AND2X2 AND2X2_918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4278_), .B(AES_CORE_DATAPATH__abc_16009_new_n4272_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4279_));
AND2X2 AND2X2_919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4282_));
AND2X2 AND2X2_92 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n247_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n117_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n248_));
AND2X2 AND2X2_920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4283_));
AND2X2 AND2X2_921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4281_), .B(AES_CORE_DATAPATH__abc_16009_new_n4285_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4286_));
AND2X2 AND2X2_922 ( .A(\key_out[26] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4289_));
AND2X2 AND2X2_923 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4292_));
AND2X2 AND2X2_924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4293_));
AND2X2 AND2X2_925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4291_), .B(AES_CORE_DATAPATH__abc_16009_new_n4295_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4296_));
AND2X2 AND2X2_926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4296_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4297_));
AND2X2 AND2X2_927 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4298_));
AND2X2 AND2X2_928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4303_), .B(AES_CORE_DATAPATH__abc_16009_new_n4301_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4304_));
AND2X2 AND2X2_929 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4305_));
AND2X2 AND2X2_93 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n251_));
AND2X2 AND2X2_930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4306_));
AND2X2 AND2X2_931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4307_));
AND2X2 AND2X2_932 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4310_), .B(AES_CORE_DATAPATH__abc_16009_new_n4304_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4311_));
AND2X2 AND2X2_933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4314_));
AND2X2 AND2X2_934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4315_));
AND2X2 AND2X2_935 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4313_), .B(AES_CORE_DATAPATH__abc_16009_new_n4317_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4318_));
AND2X2 AND2X2_936 ( .A(\key_out[27] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4318_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4321_));
AND2X2 AND2X2_937 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4324_));
AND2X2 AND2X2_938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4325_));
AND2X2 AND2X2_939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4323_), .B(AES_CORE_DATAPATH__abc_16009_new_n4327_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4328_));
AND2X2 AND2X2_94 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n252_));
AND2X2 AND2X2_940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4328_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4329_));
AND2X2 AND2X2_941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4330_));
AND2X2 AND2X2_942 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4335_), .B(AES_CORE_DATAPATH__abc_16009_new_n4333_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4336_));
AND2X2 AND2X2_943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4337_));
AND2X2 AND2X2_944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4338_));
AND2X2 AND2X2_945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4339_));
AND2X2 AND2X2_946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4342_), .B(AES_CORE_DATAPATH__abc_16009_new_n4336_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4343_));
AND2X2 AND2X2_947 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4346_));
AND2X2 AND2X2_948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4347_));
AND2X2 AND2X2_949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4345_), .B(AES_CORE_DATAPATH__abc_16009_new_n4349_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4350_));
AND2X2 AND2X2_95 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1856));
AND2X2 AND2X2_950 ( .A(\key_out[28] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4350_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4353_));
AND2X2 AND2X2_951 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4356_));
AND2X2 AND2X2_952 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4357_));
AND2X2 AND2X2_953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4355_), .B(AES_CORE_DATAPATH__abc_16009_new_n4359_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4360_));
AND2X2 AND2X2_954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4360_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4361_));
AND2X2 AND2X2_955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4362_));
AND2X2 AND2X2_956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4367_), .B(AES_CORE_DATAPATH__abc_16009_new_n4365_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4368_));
AND2X2 AND2X2_957 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4369_));
AND2X2 AND2X2_958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4370_));
AND2X2 AND2X2_959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4371_));
AND2X2 AND2X2_96 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1897));
AND2X2 AND2X2_960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4374_), .B(AES_CORE_DATAPATH__abc_16009_new_n4368_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4375_));
AND2X2 AND2X2_961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4378_));
AND2X2 AND2X2_962 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4379_));
AND2X2 AND2X2_963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4377_), .B(AES_CORE_DATAPATH__abc_16009_new_n4381_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4382_));
AND2X2 AND2X2_964 ( .A(\key_out[29] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4382_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4385_));
AND2X2 AND2X2_965 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4388_));
AND2X2 AND2X2_966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4389_));
AND2X2 AND2X2_967 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4387_), .B(AES_CORE_DATAPATH__abc_16009_new_n4391_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4392_));
AND2X2 AND2X2_968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4392_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4393_));
AND2X2 AND2X2_969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4394_));
AND2X2 AND2X2_97 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n257_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n258_));
AND2X2 AND2X2_970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4399_), .B(AES_CORE_DATAPATH__abc_16009_new_n4397_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4400_));
AND2X2 AND2X2_971 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4401_));
AND2X2 AND2X2_972 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4402_));
AND2X2 AND2X2_973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4403_));
AND2X2 AND2X2_974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4406_), .B(AES_CORE_DATAPATH__abc_16009_new_n4400_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4407_));
AND2X2 AND2X2_975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4410_));
AND2X2 AND2X2_976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4411_));
AND2X2 AND2X2_977 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4409_), .B(AES_CORE_DATAPATH__abc_16009_new_n4413_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4414_));
AND2X2 AND2X2_978 ( .A(\key_out[30] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4414_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4417_));
AND2X2 AND2X2_979 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4420_));
AND2X2 AND2X2_98 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n258_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n160_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1928));
AND2X2 AND2X2_980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4421_));
AND2X2 AND2X2_981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4419_), .B(AES_CORE_DATAPATH__abc_16009_new_n4423_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4424_));
AND2X2 AND2X2_982 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4424_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4425_));
AND2X2 AND2X2_983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4426_));
AND2X2 AND2X2_984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4431_), .B(AES_CORE_DATAPATH__abc_16009_new_n4429_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4432_));
AND2X2 AND2X2_985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3422_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4433_));
AND2X2 AND2X2_986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3430_), .B(AES_CORE_DATAPATH_col_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4434_));
AND2X2 AND2X2_987 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3438_), .B(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4435_));
AND2X2 AND2X2_988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4438_), .B(AES_CORE_DATAPATH__abc_16009_new_n4432_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4439_));
AND2X2 AND2X2_989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3445_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4442_));
AND2X2 AND2X2_99 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n94_), .B(end_aes), .Y(AES_CORE_CONTROL_UNIT_key_derivation_en));
AND2X2 AND2X2_990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3447_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4443_));
AND2X2 AND2X2_991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4441_), .B(AES_CORE_DATAPATH__abc_16009_new_n4445_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4446_));
AND2X2 AND2X2_992 ( .A(\key_out[31] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4446_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4449_));
AND2X2 AND2X2_993 ( .A(AES_CORE_DATAPATH_last_round_pp2), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4452_));
AND2X2 AND2X2_994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3460_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4453_));
AND2X2 AND2X2_995 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4451_), .B(AES_CORE_DATAPATH__abc_16009_new_n4455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4456_));
AND2X2 AND2X2_996 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4456_), .B(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n4457_));
AND2X2 AND2X2_997 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2801_), .B(AES_CORE_DATAPATH_col_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4458_));
AND2X2 AND2X2_998 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4460_));
AND2X2 AND2X2_999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3464_), .B(AES_CORE_DATAPATH__abc_16009_new_n2801_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4461_));
DFFPOSX1 DFFPOSX1_1 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__0_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__0_));
DFFPOSX1 DFFPOSX1_10 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__9_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__1_));
DFFPOSX1 DFFPOSX1_11 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__10_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__2_));
DFFPOSX1 DFFPOSX1_12 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__11_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__3_));
DFFPOSX1 DFFPOSX1_13 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__12_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__4_));
DFFPOSX1 DFFPOSX1_14 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__13_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__5_));
DFFPOSX1 DFFPOSX1_15 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__14_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__6_));
DFFPOSX1 DFFPOSX1_16 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__15_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__7_));
DFFPOSX1 DFFPOSX1_17 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__16_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__0_));
DFFPOSX1 DFFPOSX1_18 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__17_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__1_));
DFFPOSX1 DFFPOSX1_19 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__18_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__2_));
DFFPOSX1 DFFPOSX1_2 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__1_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__1_));
DFFPOSX1 DFFPOSX1_20 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__19_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__3_));
DFFPOSX1 DFFPOSX1_21 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__20_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__4_));
DFFPOSX1 DFFPOSX1_22 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__21_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__5_));
DFFPOSX1 DFFPOSX1_23 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__22_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__6_));
DFFPOSX1 DFFPOSX1_24 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__23_), .Q(AES_CORE_DATAPATH_MIX_COL_col_2__7_));
DFFPOSX1 DFFPOSX1_25 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__24_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__0_));
DFFPOSX1 DFFPOSX1_26 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__25_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__1_));
DFFPOSX1 DFFPOSX1_27 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__26_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__2_));
DFFPOSX1 DFFPOSX1_28 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__27_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__3_));
DFFPOSX1 DFFPOSX1_29 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__28_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__4_));
DFFPOSX1 DFFPOSX1_3 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__2_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__2_));
DFFPOSX1 DFFPOSX1_30 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__29_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__5_));
DFFPOSX1 DFFPOSX1_31 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__30_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__6_));
DFFPOSX1 DFFPOSX1_32 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__31_), .Q(AES_CORE_DATAPATH_MIX_COL_col_3__7_));
DFFPOSX1 DFFPOSX1_33 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_34 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_35 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_36 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_37 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_38 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_39 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_4 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__3_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__3_));
DFFPOSX1 DFFPOSX1_40 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_41 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_42 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_43 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_44 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_45 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_46 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_47 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_48 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_49 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_5 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__4_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__4_));
DFFPOSX1 DFFPOSX1_50 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_51 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_52 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_53 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_54 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_55 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_56 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_57 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_58 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_59 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_6 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__5_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__5_));
DFFPOSX1 DFFPOSX1_60 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_61 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_62 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_63 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_64 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_65 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_66 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_67 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_68 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_69 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_));
DFFPOSX1 DFFPOSX1_7 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__6_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__6_));
DFFPOSX1 DFFPOSX1_70 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_));
DFFPOSX1 DFFPOSX1_71 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_));
DFFPOSX1 DFFPOSX1_72 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_));
DFFPOSX1 DFFPOSX1_73 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_));
DFFPOSX1 DFFPOSX1_74 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_));
DFFPOSX1 DFFPOSX1_75 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_));
DFFPOSX1 DFFPOSX1_76 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_));
DFFPOSX1 DFFPOSX1_77 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_));
DFFPOSX1 DFFPOSX1_78 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_));
DFFPOSX1 DFFPOSX1_79 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_));
DFFPOSX1 DFFPOSX1_8 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__7_), .Q(AES_CORE_DATAPATH_MIX_COL_col_0__7_));
DFFPOSX1 DFFPOSX1_80 ( .CLK(clk), .D(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Q(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_));
DFFPOSX1 DFFPOSX1_9 ( .CLK(clk), .D(AES_CORE_DATAPATH__0sbox_pp2_31_0__8_), .Q(AES_CORE_DATAPATH_MIX_COL_col_1__0_));
DFFSR DFFSR_1 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_0_), .Q(AES_CORE_CONTROL_UNIT_state_0_), .R(1'h1), .S(rst_n));
DFFSR DFFSR_10 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_9_), .Q(AES_CORE_CONTROL_UNIT_state_9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_100 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_101 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_102 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_103 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_104 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_105 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_106 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_107 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_108 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_109 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_11 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_10_), .Q(AES_CORE_CONTROL_UNIT_key_gen), .R(rst_n), .S(1'h1));
DFFSR DFFSR_110 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_111 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_112 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_113 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_114 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_115 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_116 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_117 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_118 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_119 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_12 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1897), .Q(AES_CORE_CONTROL_UNIT_state_11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_120 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_121 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_122 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_123 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_124 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_125 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_126 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_127 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_128 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_129 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_13 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_12_), .Q(AES_CORE_CONTROL_UNIT_state_12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_130 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_131 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_132 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_133 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_134 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_135 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_136 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_137 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_138 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_139 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_14 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_13_), .Q(AES_CORE_CONTROL_UNIT_state_13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_140 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_141 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_142 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_143 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_144 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_145 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_146 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_147 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_148 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_1__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_149 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_15 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_14_), .Q(AES_CORE_CONTROL_UNIT_state_14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_150 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_151 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_152 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_153 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_154 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_155 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_156 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_157 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_158 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_159 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_16 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1928), .Q(AES_CORE_CONTROL_UNIT_state_15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_160 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_161 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_162 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_163 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_164 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_165 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_166 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_167 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_168 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_169 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_17 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__0_), .Q(AES_CORE_CONTROL_UNIT_rd_count_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_170 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_171 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_172 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_173 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_174 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_175 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_176 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_177 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_178 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_179 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_18 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__1_), .Q(AES_CORE_CONTROL_UNIT_rd_count_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_180 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_2__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_181 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_182 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_183 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_184 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_185 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_186 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_187 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_188 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_189 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_19 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__2_), .Q(AES_CORE_CONTROL_UNIT_rd_count_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_190 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_191 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_192 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_193 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_194 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_195 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_196 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_197 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_198 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_199 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_2 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_1_), .Q(AES_CORE_CONTROL_UNIT_state_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_20 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__0rd_count_3_0__3_), .Q(AES_CORE_CONTROL_UNIT_rd_count_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_200 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_201 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_202 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_203 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_204 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_205 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_206 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_207 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_208 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_209 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_21 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_210 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_211 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_212 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_2__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_213 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_214 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_215 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_216 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_217 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_218 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_219 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_22 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_220 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_221 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_222 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_223 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_224 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_225 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_226 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_227 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_228 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_229 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_23 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_230 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_231 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_232 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_233 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_234 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_235 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_236 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_237 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_238 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_239 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_24 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_240 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_241 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_242 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_243 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_244 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_3__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_245 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_246 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_247 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_248 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_249 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_25 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_250 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_251 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_252 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_253 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_254 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_255 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_256 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_257 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_258 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_259 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_26 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_260 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_261 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_262 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_263 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_264 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_265 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_266 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_267 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_268 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_269 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_27 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_270 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_271 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_272 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_273 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_274 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_275 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_276 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_3__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_277 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__0_), .Q(AES_CORE_DATAPATH_col_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_278 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__1_), .Q(AES_CORE_DATAPATH_col_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_279 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__2_), .Q(AES_CORE_DATAPATH_col_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_28 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_280 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__3_), .Q(AES_CORE_DATAPATH_col_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_281 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__4_), .Q(AES_CORE_DATAPATH_col_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_282 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__5_), .Q(AES_CORE_DATAPATH_col_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_283 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__6_), .Q(AES_CORE_DATAPATH_col_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_284 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__7_), .Q(AES_CORE_DATAPATH_col_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_285 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__8_), .Q(AES_CORE_DATAPATH_col_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_286 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__9_), .Q(AES_CORE_DATAPATH_col_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_287 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__10_), .Q(AES_CORE_DATAPATH_col_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_288 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__11_), .Q(AES_CORE_DATAPATH_col_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_289 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__12_), .Q(AES_CORE_DATAPATH_col_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_29 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_290 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__13_), .Q(AES_CORE_DATAPATH_col_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_291 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__14_), .Q(AES_CORE_DATAPATH_col_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_292 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__15_), .Q(AES_CORE_DATAPATH_col_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_293 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__16_), .Q(AES_CORE_DATAPATH_col_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_294 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__17_), .Q(AES_CORE_DATAPATH_col_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_295 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__18_), .Q(AES_CORE_DATAPATH_col_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_296 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__19_), .Q(AES_CORE_DATAPATH_col_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_297 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__20_), .Q(AES_CORE_DATAPATH_col_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_298 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__21_), .Q(AES_CORE_DATAPATH_col_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_299 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__22_), .Q(AES_CORE_DATAPATH_col_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_3 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_2_), .Q(AES_CORE_CONTROL_UNIT_state_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_30 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_300 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__23_), .Q(AES_CORE_DATAPATH_col_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_301 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__24_), .Q(AES_CORE_DATAPATH_col_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_302 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__25_), .Q(AES_CORE_DATAPATH_col_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_303 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__26_), .Q(AES_CORE_DATAPATH_col_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_304 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__27_), .Q(AES_CORE_DATAPATH_col_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_305 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__28_), .Q(AES_CORE_DATAPATH_col_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_306 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__29_), .Q(AES_CORE_DATAPATH_col_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_307 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__30_), .Q(AES_CORE_DATAPATH_col_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_308 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_0__31_0__31_), .Q(AES_CORE_DATAPATH_col_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_309 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__0_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_64_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_31 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_310 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__1_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_65_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_311 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__2_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_66_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_312 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__3_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_67_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_313 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__4_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_68_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_314 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__5_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_69_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_315 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__6_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_70_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_316 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__7_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_71_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_317 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__8_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_72_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_318 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__9_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_73_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_319 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__10_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_74_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_32 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_320 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__11_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_75_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_321 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__12_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_76_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_322 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__13_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_77_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_323 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__14_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_78_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_324 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__15_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_79_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_325 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__16_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_80_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_326 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__17_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_81_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_327 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__18_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_82_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_328 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__19_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_83_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_329 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__20_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_84_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_33 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_330 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__21_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_85_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_331 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__22_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_86_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_332 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__23_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_87_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_333 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__24_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_88_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_334 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__25_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_89_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_335 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__26_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_90_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_336 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__27_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_91_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_337 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__28_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_92_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_338 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__29_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_93_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_339 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__30_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_94_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_34 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_340 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_1__31_0__31_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_95_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_341 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__0_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_32_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_342 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__1_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_33_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_343 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__2_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_34_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_344 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__3_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_35_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_345 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__4_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_36_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_346 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__5_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_37_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_347 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__6_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_38_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_348 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__7_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_39_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_349 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__8_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_40_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_35 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_350 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__9_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_41_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_351 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__10_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_42_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_352 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__11_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_43_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_353 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__12_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_44_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_354 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__13_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_45_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_355 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__14_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_46_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_356 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__15_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_47_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_357 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__16_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_48_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_358 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__17_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_49_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_359 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__18_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_50_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_36 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__15_), .Q(AES_CORE_DATAPATH_key_host_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_360 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__19_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_51_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_361 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__20_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_52_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_362 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__21_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_53_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_363 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__22_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_54_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_364 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__23_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_55_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_365 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__24_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_56_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_366 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__25_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_57_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_367 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__26_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_58_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_368 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__27_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_59_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_369 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__28_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_60_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_37 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__16_), .Q(AES_CORE_DATAPATH_key_host_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_370 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__29_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_61_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_371 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__30_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_62_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_372 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_2__31_0__31_), .Q(AES_CORE_DATAPATH_SHIFT_ROW_data_in_63_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_373 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__0_), .Q(AES_CORE_DATAPATH_col_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_374 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__1_), .Q(AES_CORE_DATAPATH_col_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_375 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__2_), .Q(AES_CORE_DATAPATH_col_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_376 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__3_), .Q(AES_CORE_DATAPATH_col_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_377 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__4_), .Q(AES_CORE_DATAPATH_col_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_378 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__5_), .Q(AES_CORE_DATAPATH_col_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_379 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__6_), .Q(AES_CORE_DATAPATH_col_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_38 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__17_), .Q(AES_CORE_DATAPATH_key_host_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_380 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__7_), .Q(AES_CORE_DATAPATH_col_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_381 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__8_), .Q(AES_CORE_DATAPATH_col_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_382 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__9_), .Q(AES_CORE_DATAPATH_col_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_383 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__10_), .Q(AES_CORE_DATAPATH_col_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_384 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__11_), .Q(AES_CORE_DATAPATH_col_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_385 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__12_), .Q(AES_CORE_DATAPATH_col_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_386 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__13_), .Q(AES_CORE_DATAPATH_col_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_387 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__14_), .Q(AES_CORE_DATAPATH_col_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_388 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__15_), .Q(AES_CORE_DATAPATH_col_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_389 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__16_), .Q(AES_CORE_DATAPATH_col_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_39 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__18_), .Q(AES_CORE_DATAPATH_key_host_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_390 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__17_), .Q(AES_CORE_DATAPATH_col_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_391 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__18_), .Q(AES_CORE_DATAPATH_col_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_392 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__19_), .Q(AES_CORE_DATAPATH_col_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_393 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__20_), .Q(AES_CORE_DATAPATH_col_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_394 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__21_), .Q(AES_CORE_DATAPATH_col_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_395 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__22_), .Q(AES_CORE_DATAPATH_col_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_396 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__23_), .Q(AES_CORE_DATAPATH_col_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_397 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__24_), .Q(AES_CORE_DATAPATH_col_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_398 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__25_), .Q(AES_CORE_DATAPATH_col_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_399 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__26_), .Q(AES_CORE_DATAPATH_col_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_4 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1817), .Q(AES_CORE_CONTROL_UNIT_state_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_40 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__19_), .Q(AES_CORE_DATAPATH_key_host_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_400 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__27_), .Q(AES_CORE_DATAPATH_col_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_401 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__28_), .Q(AES_CORE_DATAPATH_col_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_402 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__29_), .Q(AES_CORE_DATAPATH_col_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_403 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__30_), .Q(AES_CORE_DATAPATH_col_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_404 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_3__31_0__31_), .Q(AES_CORE_DATAPATH_col_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_405 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__0_), .Q(AES_CORE_DATAPATH_iv_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_406 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__1_), .Q(AES_CORE_DATAPATH_iv_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_407 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__2_), .Q(AES_CORE_DATAPATH_iv_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_408 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__3_), .Q(AES_CORE_DATAPATH_iv_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_409 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__4_), .Q(AES_CORE_DATAPATH_iv_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_41 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__20_), .Q(AES_CORE_DATAPATH_key_host_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_410 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__5_), .Q(AES_CORE_DATAPATH_iv_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_411 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__6_), .Q(AES_CORE_DATAPATH_iv_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_412 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__7_), .Q(AES_CORE_DATAPATH_iv_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_413 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__8_), .Q(AES_CORE_DATAPATH_iv_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_414 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__9_), .Q(AES_CORE_DATAPATH_iv_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_415 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__10_), .Q(AES_CORE_DATAPATH_iv_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_416 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__11_), .Q(AES_CORE_DATAPATH_iv_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_417 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__12_), .Q(AES_CORE_DATAPATH_iv_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_418 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__13_), .Q(AES_CORE_DATAPATH_iv_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_419 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__14_), .Q(AES_CORE_DATAPATH_iv_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_42 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__21_), .Q(AES_CORE_DATAPATH_key_host_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_420 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__15_), .Q(AES_CORE_DATAPATH_iv_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_421 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__16_), .Q(AES_CORE_DATAPATH_iv_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_422 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__17_), .Q(AES_CORE_DATAPATH_iv_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_423 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__18_), .Q(AES_CORE_DATAPATH_iv_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_424 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__19_), .Q(AES_CORE_DATAPATH_iv_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_425 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__20_), .Q(AES_CORE_DATAPATH_iv_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_426 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__21_), .Q(AES_CORE_DATAPATH_iv_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_427 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__22_), .Q(AES_CORE_DATAPATH_iv_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_428 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__23_), .Q(AES_CORE_DATAPATH_iv_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_429 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__24_), .Q(AES_CORE_DATAPATH_iv_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_43 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__22_), .Q(AES_CORE_DATAPATH_key_host_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_430 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__25_), .Q(AES_CORE_DATAPATH_iv_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_431 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__26_), .Q(AES_CORE_DATAPATH_iv_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_432 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__27_), .Q(AES_CORE_DATAPATH_iv_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_433 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__28_), .Q(AES_CORE_DATAPATH_iv_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_434 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__29_), .Q(AES_CORE_DATAPATH_iv_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_435 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__30_), .Q(AES_CORE_DATAPATH_iv_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_436 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_3__31_0__31_), .Q(AES_CORE_DATAPATH_iv_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_437 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_438 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_439 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_44 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__23_), .Q(AES_CORE_DATAPATH_key_host_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_440 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_441 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_442 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_443 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_444 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_445 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_446 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_447 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_448 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_449 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_45 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__24_), .Q(AES_CORE_DATAPATH_key_host_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_450 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_451 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_452 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_453 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_454 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_455 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_456 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_457 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_458 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_459 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_46 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__25_), .Q(AES_CORE_DATAPATH_key_host_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_460 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_461 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_462 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_463 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_464 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_465 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_466 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_467 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_468 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_3__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_469 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_3__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_47 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__26_), .Q(AES_CORE_DATAPATH_key_host_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_470 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_3__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_471 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_3__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_472 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_3__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_473 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_3__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_474 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_3__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_475 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_3__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_476 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_3__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_477 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_3__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_478 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_3__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_479 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_3__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_48 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__27_), .Q(AES_CORE_DATAPATH_key_host_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_480 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_3__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_481 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_3__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_482 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_3__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_483 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_3__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_484 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_3__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_485 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_3__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_486 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_3__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_487 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_3__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_488 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_3__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_489 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_3__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_49 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__28_), .Q(AES_CORE_DATAPATH_key_host_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_490 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_3__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_491 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_3__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_492 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_3__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_493 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_3__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_494 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_3__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_495 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_3__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_496 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_3__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_497 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_3__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_498 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_3__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_499 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_3__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_5 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_4_), .Q(AES_CORE_CONTROL_UNIT_state_4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_50 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__29_), .Q(AES_CORE_DATAPATH_key_host_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_500 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_3__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_3__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_501 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__0_), .Q(AES_CORE_DATAPATH_iv_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_502 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__1_), .Q(AES_CORE_DATAPATH_iv_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_503 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__2_), .Q(AES_CORE_DATAPATH_iv_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_504 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__3_), .Q(AES_CORE_DATAPATH_iv_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_505 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__4_), .Q(AES_CORE_DATAPATH_iv_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_506 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__5_), .Q(AES_CORE_DATAPATH_iv_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_507 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__6_), .Q(AES_CORE_DATAPATH_iv_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_508 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__7_), .Q(AES_CORE_DATAPATH_iv_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_509 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__8_), .Q(AES_CORE_DATAPATH_iv_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_51 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__30_), .Q(AES_CORE_DATAPATH_key_host_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_510 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__9_), .Q(AES_CORE_DATAPATH_iv_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_511 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__10_), .Q(AES_CORE_DATAPATH_iv_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_512 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__11_), .Q(AES_CORE_DATAPATH_iv_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_513 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__12_), .Q(AES_CORE_DATAPATH_iv_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_514 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__13_), .Q(AES_CORE_DATAPATH_iv_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_515 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__14_), .Q(AES_CORE_DATAPATH_iv_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_516 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__15_), .Q(AES_CORE_DATAPATH_iv_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_517 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__16_), .Q(AES_CORE_DATAPATH_iv_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_518 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__17_), .Q(AES_CORE_DATAPATH_iv_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_519 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__18_), .Q(AES_CORE_DATAPATH_iv_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_52 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_0__31_0__31_), .Q(AES_CORE_DATAPATH_key_host_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_520 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__19_), .Q(AES_CORE_DATAPATH_iv_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_521 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__20_), .Q(AES_CORE_DATAPATH_iv_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_522 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__21_), .Q(AES_CORE_DATAPATH_iv_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_523 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__22_), .Q(AES_CORE_DATAPATH_iv_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_524 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__23_), .Q(AES_CORE_DATAPATH_iv_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_525 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__24_), .Q(AES_CORE_DATAPATH_iv_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_526 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__25_), .Q(AES_CORE_DATAPATH_iv_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_527 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__26_), .Q(AES_CORE_DATAPATH_iv_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_528 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__27_), .Q(AES_CORE_DATAPATH_iv_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_529 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__28_), .Q(AES_CORE_DATAPATH_iv_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_53 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_530 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__29_), .Q(AES_CORE_DATAPATH_iv_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_531 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__30_), .Q(AES_CORE_DATAPATH_iv_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_532 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_2__31_0__31_), .Q(AES_CORE_DATAPATH_iv_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_533 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_534 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_535 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_536 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_537 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_538 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_539 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_54 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_540 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_541 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_542 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_543 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_544 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_545 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_546 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_547 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_548 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_549 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_55 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_550 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_551 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_552 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_553 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_554 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_555 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_556 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_557 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_558 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_559 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_56 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_560 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_561 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_562 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_563 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_564 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_2__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_565 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_2__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_566 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_2__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_567 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_2__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_568 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_2__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_569 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_2__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_57 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__4_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_570 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_2__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_571 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_2__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_572 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_2__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_573 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_2__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_574 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_2__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_575 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_2__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_576 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_2__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_577 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_2__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_578 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_2__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_579 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_2__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_58 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__5_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_580 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_2__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_581 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_2__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_582 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_2__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_583 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_2__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_584 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_2__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_585 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_2__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_586 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_2__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_587 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_2__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_588 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_2__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_589 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_2__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_59 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__6_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_590 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_2__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_591 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_2__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_592 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_2__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_593 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_2__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_594 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_2__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_595 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_2__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_596 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_2__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_2__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_597 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__0_), .Q(AES_CORE_DATAPATH_iv_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_598 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__1_), .Q(AES_CORE_DATAPATH_iv_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_599 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__2_), .Q(AES_CORE_DATAPATH_iv_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_6 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_5_), .Q(end_aes), .R(rst_n), .S(1'h1));
DFFSR DFFSR_60 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__7_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_600 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__3_), .Q(AES_CORE_DATAPATH_iv_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_601 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__4_), .Q(AES_CORE_DATAPATH_iv_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_602 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__5_), .Q(AES_CORE_DATAPATH_iv_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_603 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__6_), .Q(AES_CORE_DATAPATH_iv_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_604 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__7_), .Q(AES_CORE_DATAPATH_iv_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_605 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__8_), .Q(AES_CORE_DATAPATH_iv_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_606 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__9_), .Q(AES_CORE_DATAPATH_iv_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_607 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__10_), .Q(AES_CORE_DATAPATH_iv_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_608 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__11_), .Q(AES_CORE_DATAPATH_iv_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_609 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__12_), .Q(AES_CORE_DATAPATH_iv_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_61 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__8_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_610 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__13_), .Q(AES_CORE_DATAPATH_iv_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_611 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__14_), .Q(AES_CORE_DATAPATH_iv_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_612 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__15_), .Q(AES_CORE_DATAPATH_iv_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_613 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__16_), .Q(AES_CORE_DATAPATH_iv_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_614 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__17_), .Q(AES_CORE_DATAPATH_iv_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_615 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__18_), .Q(AES_CORE_DATAPATH_iv_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_616 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__19_), .Q(AES_CORE_DATAPATH_iv_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_617 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__20_), .Q(AES_CORE_DATAPATH_iv_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_618 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__21_), .Q(AES_CORE_DATAPATH_iv_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_619 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__22_), .Q(AES_CORE_DATAPATH_iv_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_62 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__9_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_620 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__23_), .Q(AES_CORE_DATAPATH_iv_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_621 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__24_), .Q(AES_CORE_DATAPATH_iv_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_622 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__25_), .Q(AES_CORE_DATAPATH_iv_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_623 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__26_), .Q(AES_CORE_DATAPATH_iv_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_624 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__27_), .Q(AES_CORE_DATAPATH_iv_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_625 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__28_), .Q(AES_CORE_DATAPATH_iv_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_626 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__29_), .Q(AES_CORE_DATAPATH_iv_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_627 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__30_), .Q(AES_CORE_DATAPATH_iv_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_628 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_1__31_0__31_), .Q(AES_CORE_DATAPATH_iv_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_629 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_63 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__10_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_630 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_631 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_632 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_633 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_634 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_635 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_636 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_637 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_638 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_639 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_64 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__11_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_640 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_641 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_642 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_643 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_644 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_645 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_646 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_647 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_648 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_649 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_65 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__12_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_650 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_651 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_652 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_653 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_654 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_655 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_656 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_657 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_658 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_659 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_66 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__13_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_660 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_661 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_662 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_663 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_664 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_665 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_666 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_667 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_668 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_669 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_67 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__14_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_670 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_671 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_672 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_673 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_674 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_675 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_1__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_676 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_1__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_677 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_1__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_678 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_1__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_679 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_1__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_68 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__15_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_680 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_1__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_681 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_1__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_682 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_1__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_683 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_1__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_684 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_1__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_685 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_1__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_686 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_1__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_687 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_1__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_688 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_1__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_689 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_1__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_69 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__16_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_690 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_1__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_691 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_1__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_692 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_1__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_1__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_693 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__0_), .Q(AES_CORE_DATAPATH_iv_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_694 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__1_), .Q(AES_CORE_DATAPATH_iv_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_695 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__2_), .Q(AES_CORE_DATAPATH_iv_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_696 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__3_), .Q(AES_CORE_DATAPATH_iv_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_697 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__4_), .Q(AES_CORE_DATAPATH_iv_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_698 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__5_), .Q(AES_CORE_DATAPATH_iv_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_699 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__6_), .Q(AES_CORE_DATAPATH_iv_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_7 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_6_), .Q(AES_CORE_CONTROL_UNIT_state_6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_70 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__17_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_700 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__7_), .Q(AES_CORE_DATAPATH_iv_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_701 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__8_), .Q(AES_CORE_DATAPATH_iv_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_702 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__9_), .Q(AES_CORE_DATAPATH_iv_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_703 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__10_), .Q(AES_CORE_DATAPATH_iv_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_704 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__11_), .Q(AES_CORE_DATAPATH_iv_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_705 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__12_), .Q(AES_CORE_DATAPATH_iv_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_706 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__13_), .Q(AES_CORE_DATAPATH_iv_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_707 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__14_), .Q(AES_CORE_DATAPATH_iv_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_708 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__15_), .Q(AES_CORE_DATAPATH_iv_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_709 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__16_), .Q(AES_CORE_DATAPATH_iv_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_71 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__18_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_710 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__17_), .Q(AES_CORE_DATAPATH_iv_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_711 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__18_), .Q(AES_CORE_DATAPATH_iv_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_712 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__19_), .Q(AES_CORE_DATAPATH_iv_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_713 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__20_), .Q(AES_CORE_DATAPATH_iv_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_714 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__21_), .Q(AES_CORE_DATAPATH_iv_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_715 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__22_), .Q(AES_CORE_DATAPATH_iv_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_716 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__23_), .Q(AES_CORE_DATAPATH_iv_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_717 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__24_), .Q(AES_CORE_DATAPATH_iv_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_718 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__25_), .Q(AES_CORE_DATAPATH_iv_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_719 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__26_), .Q(AES_CORE_DATAPATH_iv_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_72 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__19_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_720 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__27_), .Q(AES_CORE_DATAPATH_iv_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_721 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__28_), .Q(AES_CORE_DATAPATH_iv_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_722 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__29_), .Q(AES_CORE_DATAPATH_iv_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_723 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__30_), .Q(AES_CORE_DATAPATH_iv_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_724 ( .CLK(clk), .D(AES_CORE_DATAPATH__0iv_0__31_0__31_), .Q(AES_CORE_DATAPATH_iv_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_725 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_726 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_727 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_728 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_729 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_73 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__20_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_730 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_731 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_732 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_733 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_734 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_735 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_736 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_737 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_738 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_739 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_74 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__21_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_740 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_741 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_742 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_743 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_744 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_745 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_746 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_747 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_748 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_749 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_75 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__22_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_750 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_751 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_752 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_753 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_754 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_755 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_756 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_0__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_757 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__0_), .Q(AES_CORE_DATAPATH_bkp_1_0__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_758 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__1_), .Q(AES_CORE_DATAPATH_bkp_1_0__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_759 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__2_), .Q(AES_CORE_DATAPATH_bkp_1_0__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_76 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__23_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_760 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__3_), .Q(AES_CORE_DATAPATH_bkp_1_0__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_761 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__4_), .Q(AES_CORE_DATAPATH_bkp_1_0__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_762 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__5_), .Q(AES_CORE_DATAPATH_bkp_1_0__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_763 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__6_), .Q(AES_CORE_DATAPATH_bkp_1_0__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_764 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__7_), .Q(AES_CORE_DATAPATH_bkp_1_0__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_765 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__8_), .Q(AES_CORE_DATAPATH_bkp_1_0__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_766 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__9_), .Q(AES_CORE_DATAPATH_bkp_1_0__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_767 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__10_), .Q(AES_CORE_DATAPATH_bkp_1_0__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_768 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__11_), .Q(AES_CORE_DATAPATH_bkp_1_0__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_769 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__12_), .Q(AES_CORE_DATAPATH_bkp_1_0__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_77 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__24_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_770 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__13_), .Q(AES_CORE_DATAPATH_bkp_1_0__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_771 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__14_), .Q(AES_CORE_DATAPATH_bkp_1_0__14_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_772 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__15_), .Q(AES_CORE_DATAPATH_bkp_1_0__15_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_773 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__16_), .Q(AES_CORE_DATAPATH_bkp_1_0__16_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_774 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__17_), .Q(AES_CORE_DATAPATH_bkp_1_0__17_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_775 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__18_), .Q(AES_CORE_DATAPATH_bkp_1_0__18_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_776 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__19_), .Q(AES_CORE_DATAPATH_bkp_1_0__19_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_777 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__20_), .Q(AES_CORE_DATAPATH_bkp_1_0__20_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_778 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__21_), .Q(AES_CORE_DATAPATH_bkp_1_0__21_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_779 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__22_), .Q(AES_CORE_DATAPATH_bkp_1_0__22_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_78 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__25_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_780 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__23_), .Q(AES_CORE_DATAPATH_bkp_1_0__23_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_781 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__24_), .Q(AES_CORE_DATAPATH_bkp_1_0__24_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_782 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__25_), .Q(AES_CORE_DATAPATH_bkp_1_0__25_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_783 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__26_), .Q(AES_CORE_DATAPATH_bkp_1_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_784 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__27_), .Q(AES_CORE_DATAPATH_bkp_1_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_785 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__28_), .Q(AES_CORE_DATAPATH_bkp_1_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_786 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__29_), .Q(AES_CORE_DATAPATH_bkp_1_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_787 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__30_), .Q(AES_CORE_DATAPATH_bkp_1_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_788 ( .CLK(clk), .D(AES_CORE_DATAPATH__0bkp_1_0__31_0__31_), .Q(AES_CORE_DATAPATH_bkp_1_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_789 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__0_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_79 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__26_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_790 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__1_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_791 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__2_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_792 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp1_3_0__3_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_793 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__0_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_794 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__1_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_795 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__2_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_796 ( .CLK(clk), .D(AES_CORE_DATAPATH__0col_en_cnt_unit_pp2_3_0__3_), .Q(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_797 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__0_), .Q(AES_CORE_DATAPATH_key_en_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_798 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__1_), .Q(AES_CORE_DATAPATH_key_en_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_799 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__2_), .Q(AES_CORE_DATAPATH_key_en_pp1_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_8 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_118_implement_pattern_cache_1856), .Q(AES_CORE_CONTROL_UNIT_state_7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_80 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__27_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_800 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_en_pp1_3_0__3_), .Q(AES_CORE_DATAPATH_key_en_pp1_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_801 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_0_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_802 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_1_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_803 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_2_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_804 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rd_count_3_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_805 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_col_sel_0_), .Q(AES_CORE_DATAPATH_col_sel_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_806 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_col_sel_1_), .Q(AES_CORE_DATAPATH_col_sel_pp1_1_), .R(1'h1), .S(rst_n));
DFFSR DFFSR_807 ( .CLK(clk), .D(AES_CORE_DATAPATH_col_sel_pp1_0_), .Q(AES_CORE_DATAPATH_col_sel_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_808 ( .CLK(clk), .D(AES_CORE_DATAPATH_col_sel_pp1_1_), .Q(AES_CORE_DATAPATH_col_sel_pp2_1_), .R(1'h1), .S(rst_n));
DFFSR DFFSR_809 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_key_out_sel_0_), .Q(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_81 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__28_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_810 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_key_out_sel_1_), .Q(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_811 ( .CLK(clk), .D(AES_CORE_DATAPATH_key_out_sel_pp1_0_), .Q(AES_CORE_DATAPATH_key_out_sel_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_812 ( .CLK(clk), .D(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Q(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_813 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rk_sel_0_), .Q(AES_CORE_DATAPATH_rk_sel_pp1_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_814 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_rk_sel_1_), .Q(AES_CORE_DATAPATH_rk_sel_pp1_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_815 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_sel_pp1_0_), .Q(AES_CORE_DATAPATH_rk_sel_pp2_0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_816 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_sel_pp1_1_), .Q(AES_CORE_DATAPATH_rk_sel_pp2_1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_817 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_key_sel), .Q(AES_CORE_DATAPATH_key_sel_pp1), .R(rst_n), .S(1'h1));
DFFSR DFFSR_818 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_out_sel), .Q(AES_CORE_DATAPATH_rk_out_sel_pp1), .R(1'h1), .S(rst_n));
DFFSR DFFSR_819 ( .CLK(clk), .D(AES_CORE_DATAPATH_rk_out_sel_pp1), .Q(AES_CORE_DATAPATH_rk_out_sel_pp2), .R(1'h1), .S(rst_n));
DFFSR DFFSR_82 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__29_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_820 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT_last_round), .Q(AES_CORE_DATAPATH_last_round_pp1), .R(1'h1), .S(rst_n));
DFFSR DFFSR_821 ( .CLK(clk), .D(AES_CORE_DATAPATH_last_round_pp1), .Q(AES_CORE_DATAPATH_last_round_pp2), .R(rst_n), .S(1'h1));
DFFSR DFFSR_83 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__30_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_84 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_0__31_0__31_), .Q(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_85 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__0_), .Q(AES_CORE_DATAPATH_key_host_1__0_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_86 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__1_), .Q(AES_CORE_DATAPATH_key_host_1__1_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_87 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__2_), .Q(AES_CORE_DATAPATH_key_host_1__2_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_88 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__3_), .Q(AES_CORE_DATAPATH_key_host_1__3_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_89 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__4_), .Q(AES_CORE_DATAPATH_key_host_1__4_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_9 ( .CLK(clk), .D(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_8_), .Q(AES_CORE_CONTROL_UNIT_state_8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_90 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__5_), .Q(AES_CORE_DATAPATH_key_host_1__5_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_91 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__6_), .Q(AES_CORE_DATAPATH_key_host_1__6_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_92 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__7_), .Q(AES_CORE_DATAPATH_key_host_1__7_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_93 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__8_), .Q(AES_CORE_DATAPATH_key_host_1__8_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_94 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__9_), .Q(AES_CORE_DATAPATH_key_host_1__9_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_95 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__10_), .Q(AES_CORE_DATAPATH_key_host_1__10_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_96 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__11_), .Q(AES_CORE_DATAPATH_key_host_1__11_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_97 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__12_), .Q(AES_CORE_DATAPATH_key_host_1__12_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_98 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__13_), .Q(AES_CORE_DATAPATH_key_host_1__13_), .R(rst_n), .S(1'h1));
DFFSR DFFSR_99 ( .CLK(clk), .D(AES_CORE_DATAPATH__0key_host_1__31_0__14_), .Q(AES_CORE_DATAPATH_key_host_1__14_), .R(rst_n), .S(1'h1));
INVX1 INVX1_1 ( .A(\addr[1] ), .Y(_abc_15574_new_n11_));
INVX1 INVX1_10 ( .A(disable_core), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n86_));
INVX1 INVX1_100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3085_));
INVX1 INVX1_1000 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n118_));
INVX1 INVX1_1001 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n123_));
INVX1 INVX1_1002 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n131_));
INVX1 INVX1_1003 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_));
INVX1 INVX1_1004 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_));
INVX1 INVX1_1005 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n150_));
INVX1 INVX1_1006 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_));
INVX1 INVX1_1007 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n159_));
INVX1 INVX1_1008 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n160_));
INVX1 INVX1_1009 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n163_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n164_));
INVX1 INVX1_101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3087_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3088_));
INVX1 INVX1_1010 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n166_));
INVX1 INVX1_1011 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n169_));
INVX1 INVX1_1012 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n170_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n171_));
INVX1 INVX1_1013 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n178_));
INVX1 INVX1_1014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n181_));
INVX1 INVX1_1015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n183_));
INVX1 INVX1_1016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n186_));
INVX1 INVX1_1017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n188_));
INVX1 INVX1_1018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n190_));
INVX1 INVX1_1019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n193_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n194_));
INVX1 INVX1_102 ( .A(\key_out[14] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3096_));
INVX1 INVX1_1020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n197_));
INVX1 INVX1_1021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n198_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n199_));
INVX1 INVX1_1022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_));
INVX1 INVX1_1023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n214_));
INVX1 INVX1_1024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n215_));
INVX1 INVX1_1025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n216_));
INVX1 INVX1_1026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n221_));
INVX1 INVX1_1027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n233_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n234_));
INVX1 INVX1_1028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n237_));
INVX1 INVX1_1029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n239_));
INVX1 INVX1_103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3102_));
INVX1 INVX1_1030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_));
INVX1 INVX1_1031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n248_));
INVX1 INVX1_1032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n249_));
INVX1 INVX1_1033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n255_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n256_));
INVX1 INVX1_1034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n259_));
INVX1 INVX1_1035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n263_));
INVX1 INVX1_1036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n265_));
INVX1 INVX1_1037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n269_));
INVX1 INVX1_1038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n272_));
INVX1 INVX1_1039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n275_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n276_));
INVX1 INVX1_104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3104_));
INVX1 INVX1_1040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n279_));
INVX1 INVX1_1041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n285_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n286_));
INVX1 INVX1_1042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n289_));
INVX1 INVX1_1043 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n290_));
INVX1 INVX1_1044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n294_));
INVX1 INVX1_1045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n299_));
INVX1 INVX1_1046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n304_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n305_));
INVX1 INVX1_1047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n308_));
INVX1 INVX1_1048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n310_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n311_));
INVX1 INVX1_1049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n314_));
INVX1 INVX1_105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3106_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3107_));
INVX1 INVX1_1050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n316_));
INVX1 INVX1_1051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n320_));
INVX1 INVX1_1052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n329_));
INVX1 INVX1_1053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n332_));
INVX1 INVX1_1054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_));
INVX1 INVX1_1055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n338_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n339_));
INVX1 INVX1_1056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n343_));
INVX1 INVX1_1057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n349_));
INVX1 INVX1_1058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n356_));
INVX1 INVX1_1059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n360_));
INVX1 INVX1_106 ( .A(\key_out[15] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3114_));
INVX1 INVX1_1060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n366_));
INVX1 INVX1_1061 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n378_));
INVX1 INVX1_1062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n385_));
INVX1 INVX1_1063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n390_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n391_));
INVX1 INVX1_1064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n394_));
INVX1 INVX1_1065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n416_));
INVX1 INVX1_1066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n438_));
INVX1 INVX1_1067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n443_));
INVX1 INVX1_1068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n446_));
INVX1 INVX1_1069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n447_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n448_));
INVX1 INVX1_107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3120_));
INVX1 INVX1_1070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n450_));
INVX1 INVX1_1071 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n453_));
INVX1 INVX1_1072 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n457_));
INVX1 INVX1_1073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n460_));
INVX1 INVX1_1074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n468_));
INVX1 INVX1_1075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n475_));
INVX1 INVX1_1076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n478_));
INVX1 INVX1_1077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n480_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n481_));
INVX1 INVX1_1078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n485_));
INVX1 INVX1_1079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n488_));
INVX1 INVX1_108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3122_));
INVX1 INVX1_1080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n491_));
INVX1 INVX1_1081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n498_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n499_));
INVX1 INVX1_1082 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n503_));
INVX1 INVX1_1083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n507_));
INVX1 INVX1_1084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n509_));
INVX1 INVX1_1085 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n508_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n513_));
INVX1 INVX1_1086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n514_));
INVX1 INVX1_1087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n519_));
INVX1 INVX1_1088 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n520_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n521_));
INVX1 INVX1_1089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n523_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n524_));
INVX1 INVX1_109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3125_));
INVX1 INVX1_1090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n526_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n527_));
INVX1 INVX1_1091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n530_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n532_));
INVX1 INVX1_1092 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n536_));
INVX1 INVX1_1093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n538_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n539_));
INVX1 INVX1_1094 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n541_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n542_));
INVX1 INVX1_1095 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n545_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n546_));
INVX1 INVX1_1096 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n551_));
INVX1 INVX1_1097 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n50_));
INVX1 INVX1_1098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n52_));
INVX1 INVX1_1099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n55_));
INVX1 INVX1_11 ( .A(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n87_));
INVX1 INVX1_110 ( .A(\key_out[16] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3131_));
INVX1 INVX1_1100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n57_));
INVX1 INVX1_1101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n60_));
INVX1 INVX1_1102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n62_));
INVX1 INVX1_1103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_));
INVX1 INVX1_1104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n67_));
INVX1 INVX1_1105 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n72_));
INVX1 INVX1_1106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n73_));
INVX1 INVX1_1107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_));
INVX1 INVX1_1108 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n81_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n82_));
INVX1 INVX1_1109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_));
INVX1 INVX1_111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3138_));
INVX1 INVX1_1110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n94_));
INVX1 INVX1_1111 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n98_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n99_));
INVX1 INVX1_1112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n100_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_));
INVX1 INVX1_1113 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n102_));
INVX1 INVX1_1114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n107_));
INVX1 INVX1_1115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n113_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n114_));
INVX1 INVX1_1116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n118_));
INVX1 INVX1_1117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n123_));
INVX1 INVX1_1118 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n131_));
INVX1 INVX1_1119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_));
INVX1 INVX1_112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3140_));
INVX1 INVX1_1120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_));
INVX1 INVX1_1121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n150_));
INVX1 INVX1_1122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_));
INVX1 INVX1_1123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n159_));
INVX1 INVX1_1124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n160_));
INVX1 INVX1_1125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n163_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n164_));
INVX1 INVX1_1126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n166_));
INVX1 INVX1_1127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n169_));
INVX1 INVX1_1128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n170_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n171_));
INVX1 INVX1_1129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n178_));
INVX1 INVX1_113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3143_));
INVX1 INVX1_1130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n181_));
INVX1 INVX1_1131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n183_));
INVX1 INVX1_1132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n186_));
INVX1 INVX1_1133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n188_));
INVX1 INVX1_1134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n190_));
INVX1 INVX1_1135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n193_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n194_));
INVX1 INVX1_1136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n197_));
INVX1 INVX1_1137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n198_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n199_));
INVX1 INVX1_1138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_));
INVX1 INVX1_1139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n214_));
INVX1 INVX1_114 ( .A(\key_out[17] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3150_));
INVX1 INVX1_1140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n215_));
INVX1 INVX1_1141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n216_));
INVX1 INVX1_1142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n221_));
INVX1 INVX1_1143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n233_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n234_));
INVX1 INVX1_1144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n237_));
INVX1 INVX1_1145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n239_));
INVX1 INVX1_1146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_));
INVX1 INVX1_1147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n248_));
INVX1 INVX1_1148 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n249_));
INVX1 INVX1_1149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n255_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n256_));
INVX1 INVX1_115 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3156_));
INVX1 INVX1_1150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n259_));
INVX1 INVX1_1151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n263_));
INVX1 INVX1_1152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n265_));
INVX1 INVX1_1153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n269_));
INVX1 INVX1_1154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n272_));
INVX1 INVX1_1155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n275_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n276_));
INVX1 INVX1_1156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n279_));
INVX1 INVX1_1157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n285_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n286_));
INVX1 INVX1_1158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n289_));
INVX1 INVX1_1159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n290_));
INVX1 INVX1_116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3158_));
INVX1 INVX1_1160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n294_));
INVX1 INVX1_1161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n299_));
INVX1 INVX1_1162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n304_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n305_));
INVX1 INVX1_1163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n308_));
INVX1 INVX1_1164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n310_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n311_));
INVX1 INVX1_1165 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n314_));
INVX1 INVX1_1166 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n316_));
INVX1 INVX1_1167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n320_));
INVX1 INVX1_1168 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n329_));
INVX1 INVX1_1169 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n332_));
INVX1 INVX1_117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3160_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3161_));
INVX1 INVX1_1170 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_));
INVX1 INVX1_1171 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n338_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n339_));
INVX1 INVX1_1172 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n343_));
INVX1 INVX1_1173 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n349_));
INVX1 INVX1_1174 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n356_));
INVX1 INVX1_1175 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n360_));
INVX1 INVX1_1176 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n366_));
INVX1 INVX1_1177 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n378_));
INVX1 INVX1_1178 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n385_));
INVX1 INVX1_1179 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n390_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n391_));
INVX1 INVX1_118 ( .A(\key_out[18] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3168_));
INVX1 INVX1_1180 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n394_));
INVX1 INVX1_1181 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n416_));
INVX1 INVX1_1182 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n438_));
INVX1 INVX1_1183 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n443_));
INVX1 INVX1_1184 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n446_));
INVX1 INVX1_1185 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n447_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n448_));
INVX1 INVX1_1186 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n450_));
INVX1 INVX1_1187 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n453_));
INVX1 INVX1_1188 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n457_));
INVX1 INVX1_1189 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n460_));
INVX1 INVX1_119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3174_));
INVX1 INVX1_1190 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n468_));
INVX1 INVX1_1191 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n475_));
INVX1 INVX1_1192 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n478_));
INVX1 INVX1_1193 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n480_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n481_));
INVX1 INVX1_1194 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n485_));
INVX1 INVX1_1195 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n488_));
INVX1 INVX1_1196 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n491_));
INVX1 INVX1_1197 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n498_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n499_));
INVX1 INVX1_1198 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n503_));
INVX1 INVX1_1199 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n507_));
INVX1 INVX1_12 ( .A(\op_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n92_));
INVX1 INVX1_120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3176_));
INVX1 INVX1_1200 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n509_));
INVX1 INVX1_1201 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n508_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n513_));
INVX1 INVX1_1202 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n514_));
INVX1 INVX1_1203 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n519_));
INVX1 INVX1_1204 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n520_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n521_));
INVX1 INVX1_1205 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n523_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n524_));
INVX1 INVX1_1206 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n526_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n527_));
INVX1 INVX1_1207 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n530_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n532_));
INVX1 INVX1_1208 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n536_));
INVX1 INVX1_1209 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n538_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n539_));
INVX1 INVX1_121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3178_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3179_));
INVX1 INVX1_1210 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n541_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n542_));
INVX1 INVX1_1211 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n545_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n546_));
INVX1 INVX1_1212 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n551_));
INVX1 INVX1_1213 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n50_));
INVX1 INVX1_1214 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n52_));
INVX1 INVX1_1215 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n55_));
INVX1 INVX1_1216 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n57_));
INVX1 INVX1_1217 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n60_));
INVX1 INVX1_1218 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n62_));
INVX1 INVX1_1219 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_));
INVX1 INVX1_122 ( .A(\key_out[19] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3186_));
INVX1 INVX1_1220 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n67_));
INVX1 INVX1_1221 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n72_));
INVX1 INVX1_1222 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n73_));
INVX1 INVX1_1223 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_));
INVX1 INVX1_1224 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n81_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n82_));
INVX1 INVX1_1225 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_));
INVX1 INVX1_1226 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n94_));
INVX1 INVX1_1227 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n98_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n99_));
INVX1 INVX1_1228 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n100_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_));
INVX1 INVX1_1229 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n102_));
INVX1 INVX1_123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3192_));
INVX1 INVX1_1230 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n107_));
INVX1 INVX1_1231 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n113_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n114_));
INVX1 INVX1_1232 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n118_));
INVX1 INVX1_1233 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n123_));
INVX1 INVX1_1234 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n131_));
INVX1 INVX1_1235 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_));
INVX1 INVX1_1236 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_));
INVX1 INVX1_1237 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n150_));
INVX1 INVX1_1238 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_));
INVX1 INVX1_1239 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n159_));
INVX1 INVX1_124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3194_));
INVX1 INVX1_1240 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n160_));
INVX1 INVX1_1241 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n163_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n164_));
INVX1 INVX1_1242 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n166_));
INVX1 INVX1_1243 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n169_));
INVX1 INVX1_1244 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n170_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n171_));
INVX1 INVX1_1245 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n178_));
INVX1 INVX1_1246 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n181_));
INVX1 INVX1_1247 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n183_));
INVX1 INVX1_1248 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n186_));
INVX1 INVX1_1249 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n188_));
INVX1 INVX1_125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3196_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3197_));
INVX1 INVX1_1250 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n190_));
INVX1 INVX1_1251 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n193_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n194_));
INVX1 INVX1_1252 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n197_));
INVX1 INVX1_1253 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n198_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n199_));
INVX1 INVX1_1254 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_));
INVX1 INVX1_1255 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n214_));
INVX1 INVX1_1256 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n215_));
INVX1 INVX1_1257 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n216_));
INVX1 INVX1_1258 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n221_));
INVX1 INVX1_1259 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n233_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n234_));
INVX1 INVX1_126 ( .A(\key_out[20] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3204_));
INVX1 INVX1_1260 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n237_));
INVX1 INVX1_1261 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n239_));
INVX1 INVX1_1262 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_));
INVX1 INVX1_1263 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n248_));
INVX1 INVX1_1264 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n249_));
INVX1 INVX1_1265 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n255_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n256_));
INVX1 INVX1_1266 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n259_));
INVX1 INVX1_1267 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n263_));
INVX1 INVX1_1268 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n265_));
INVX1 INVX1_1269 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n269_));
INVX1 INVX1_127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3210_));
INVX1 INVX1_1270 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n272_));
INVX1 INVX1_1271 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n275_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n276_));
INVX1 INVX1_1272 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n279_));
INVX1 INVX1_1273 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n285_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n286_));
INVX1 INVX1_1274 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n289_));
INVX1 INVX1_1275 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n290_));
INVX1 INVX1_1276 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n294_));
INVX1 INVX1_1277 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n299_));
INVX1 INVX1_1278 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n304_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n305_));
INVX1 INVX1_1279 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n308_));
INVX1 INVX1_128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3212_));
INVX1 INVX1_1280 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n310_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n311_));
INVX1 INVX1_1281 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n314_));
INVX1 INVX1_1282 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n316_));
INVX1 INVX1_1283 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n320_));
INVX1 INVX1_1284 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n329_));
INVX1 INVX1_1285 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n332_));
INVX1 INVX1_1286 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_));
INVX1 INVX1_1287 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n338_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n339_));
INVX1 INVX1_1288 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n343_));
INVX1 INVX1_1289 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n349_));
INVX1 INVX1_129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3214_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3215_));
INVX1 INVX1_1290 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n356_));
INVX1 INVX1_1291 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n360_));
INVX1 INVX1_1292 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n366_));
INVX1 INVX1_1293 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n378_));
INVX1 INVX1_1294 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n385_));
INVX1 INVX1_1295 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n390_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n391_));
INVX1 INVX1_1296 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n394_));
INVX1 INVX1_1297 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n416_));
INVX1 INVX1_1298 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n438_));
INVX1 INVX1_1299 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n443_));
INVX1 INVX1_13 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n94_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n99_));
INVX1 INVX1_130 ( .A(\key_out[21] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3222_));
INVX1 INVX1_1300 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n446_));
INVX1 INVX1_1301 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n447_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n448_));
INVX1 INVX1_1302 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n450_));
INVX1 INVX1_1303 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n453_));
INVX1 INVX1_1304 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n457_));
INVX1 INVX1_1305 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n460_));
INVX1 INVX1_1306 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n468_));
INVX1 INVX1_1307 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n475_));
INVX1 INVX1_1308 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n478_));
INVX1 INVX1_1309 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n480_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n481_));
INVX1 INVX1_131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3228_));
INVX1 INVX1_1310 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n485_));
INVX1 INVX1_1311 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n488_));
INVX1 INVX1_1312 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n491_));
INVX1 INVX1_1313 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n498_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n499_));
INVX1 INVX1_1314 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n503_));
INVX1 INVX1_1315 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n507_));
INVX1 INVX1_1316 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n509_));
INVX1 INVX1_1317 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n508_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n513_));
INVX1 INVX1_1318 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n514_));
INVX1 INVX1_1319 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n519_));
INVX1 INVX1_132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3230_));
INVX1 INVX1_1320 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n520_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n521_));
INVX1 INVX1_1321 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n523_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n524_));
INVX1 INVX1_1322 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n526_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n527_));
INVX1 INVX1_1323 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n530_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n532_));
INVX1 INVX1_1324 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n536_));
INVX1 INVX1_1325 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n538_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n539_));
INVX1 INVX1_1326 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n541_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n542_));
INVX1 INVX1_1327 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n545_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n546_));
INVX1 INVX1_1328 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n551_));
INVX1 INVX1_1329 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n50_));
INVX1 INVX1_133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3232_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3233_));
INVX1 INVX1_1330 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n52_));
INVX1 INVX1_1331 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n55_));
INVX1 INVX1_1332 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n57_));
INVX1 INVX1_1333 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n60_));
INVX1 INVX1_1334 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n62_));
INVX1 INVX1_1335 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_));
INVX1 INVX1_1336 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n67_));
INVX1 INVX1_1337 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n72_));
INVX1 INVX1_1338 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n73_));
INVX1 INVX1_1339 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_));
INVX1 INVX1_134 ( .A(\key_out[22] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3240_));
INVX1 INVX1_1340 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n81_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n82_));
INVX1 INVX1_1341 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_));
INVX1 INVX1_1342 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n94_));
INVX1 INVX1_1343 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n98_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n99_));
INVX1 INVX1_1344 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n100_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_));
INVX1 INVX1_1345 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n102_));
INVX1 INVX1_1346 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n107_));
INVX1 INVX1_1347 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n113_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n114_));
INVX1 INVX1_1348 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n117_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n118_));
INVX1 INVX1_1349 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n122_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n123_));
INVX1 INVX1_135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3246_));
INVX1 INVX1_1350 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n130_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n131_));
INVX1 INVX1_1351 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_));
INVX1 INVX1_1352 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_));
INVX1 INVX1_1353 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n148_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n150_));
INVX1 INVX1_1354 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n154_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_));
INVX1 INVX1_1355 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n159_));
INVX1 INVX1_1356 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n160_));
INVX1 INVX1_1357 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n163_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n164_));
INVX1 INVX1_1358 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n165_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n166_));
INVX1 INVX1_1359 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n168_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n169_));
INVX1 INVX1_136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3248_));
INVX1 INVX1_1360 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n170_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n171_));
INVX1 INVX1_1361 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n178_));
INVX1 INVX1_1362 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n181_));
INVX1 INVX1_1363 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n183_));
INVX1 INVX1_1364 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n186_));
INVX1 INVX1_1365 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n188_));
INVX1 INVX1_1366 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n190_));
INVX1 INVX1_1367 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n193_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n194_));
INVX1 INVX1_1368 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n172_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n197_));
INVX1 INVX1_1369 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n198_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n199_));
INVX1 INVX1_137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3250_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3251_));
INVX1 INVX1_1370 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_));
INVX1 INVX1_1371 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n214_));
INVX1 INVX1_1372 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n215_));
INVX1 INVX1_1373 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n175_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n216_));
INVX1 INVX1_1374 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n192_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n221_));
INVX1 INVX1_1375 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n233_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n234_));
INVX1 INVX1_1376 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n237_));
INVX1 INVX1_1377 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n239_));
INVX1 INVX1_1378 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_));
INVX1 INVX1_1379 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n248_));
INVX1 INVX1_138 ( .A(\key_out[23] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3258_));
INVX1 INVX1_1380 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n249_));
INVX1 INVX1_1381 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n255_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n256_));
INVX1 INVX1_1382 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n259_));
INVX1 INVX1_1383 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n263_));
INVX1 INVX1_1384 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n265_));
INVX1 INVX1_1385 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n268_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n269_));
INVX1 INVX1_1386 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n271_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n272_));
INVX1 INVX1_1387 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n275_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n276_));
INVX1 INVX1_1388 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n279_));
INVX1 INVX1_1389 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n285_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n286_));
INVX1 INVX1_139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3264_));
INVX1 INVX1_1390 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n288_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n289_));
INVX1 INVX1_1391 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n274_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n290_));
INVX1 INVX1_1392 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n294_));
INVX1 INVX1_1393 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n299_));
INVX1 INVX1_1394 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n304_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n305_));
INVX1 INVX1_1395 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n231_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n308_));
INVX1 INVX1_1396 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n310_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n311_));
INVX1 INVX1_1397 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n313_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n314_));
INVX1 INVX1_1398 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n307_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n316_));
INVX1 INVX1_1399 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n319_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n320_));
INVX1 INVX1_14 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n93_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n102_));
INVX1 INVX1_140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3265_));
INVX1 INVX1_1400 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n328_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n329_));
INVX1 INVX1_1401 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n332_));
INVX1 INVX1_1402 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_));
INVX1 INVX1_1403 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n338_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n339_));
INVX1 INVX1_1404 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n343_));
INVX1 INVX1_1405 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n349_));
INVX1 INVX1_1406 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n355_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n356_));
INVX1 INVX1_1407 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n360_));
INVX1 INVX1_1408 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n366_));
INVX1 INVX1_1409 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n378_));
INVX1 INVX1_141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3267_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3268_));
INVX1 INVX1_1410 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n385_));
INVX1 INVX1_1411 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n390_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n391_));
INVX1 INVX1_1412 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n394_));
INVX1 INVX1_1413 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n416_));
INVX1 INVX1_1414 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n438_));
INVX1 INVX1_1415 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n443_));
INVX1 INVX1_1416 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n446_));
INVX1 INVX1_1417 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n447_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n448_));
INVX1 INVX1_1418 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n449_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n450_));
INVX1 INVX1_1419 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n452_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n453_));
INVX1 INVX1_142 ( .A(\key_out[24] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3275_));
INVX1 INVX1_1420 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n456_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n457_));
INVX1 INVX1_1421 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n459_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n460_));
INVX1 INVX1_1422 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n468_));
INVX1 INVX1_1423 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n474_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n475_));
INVX1 INVX1_1424 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n477_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n478_));
INVX1 INVX1_1425 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n480_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n481_));
INVX1 INVX1_1426 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n445_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n485_));
INVX1 INVX1_1427 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n487_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n488_));
INVX1 INVX1_1428 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n491_));
INVX1 INVX1_1429 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n498_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n499_));
INVX1 INVX1_143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3282_));
INVX1 INVX1_1430 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n494_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n503_));
INVX1 INVX1_1431 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n507_));
INVX1 INVX1_1432 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n509_));
INVX1 INVX1_1433 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n508_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n513_));
INVX1 INVX1_1434 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n514_));
INVX1 INVX1_1435 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n519_));
INVX1 INVX1_1436 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n520_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n521_));
INVX1 INVX1_1437 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n523_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n524_));
INVX1 INVX1_1438 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n526_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n527_));
INVX1 INVX1_1439 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n530_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n532_));
INVX1 INVX1_144 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3283_));
INVX1 INVX1_1440 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n536_));
INVX1 INVX1_1441 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n538_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n539_));
INVX1 INVX1_1442 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n541_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n542_));
INVX1 INVX1_1443 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n545_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n546_));
INVX1 INVX1_1444 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n551_));
INVX1 INVX1_1445 ( .A(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n67_));
INVX1 INVX1_1446 ( .A(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n70_));
INVX1 INVX1_1447 ( .A(\data_type[1] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n67_));
INVX1 INVX1_1448 ( .A(\data_type[0] ), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n70_));
INVX1 INVX1_145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3285_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3286_));
INVX1 INVX1_146 ( .A(\key_out[25] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3294_));
INVX1 INVX1_147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3300_));
INVX1 INVX1_148 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3301_));
INVX1 INVX1_149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3303_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3304_));
INVX1 INVX1_15 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n76_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n113_));
INVX1 INVX1_150 ( .A(\key_out[26] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3312_));
INVX1 INVX1_151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3318_));
INVX1 INVX1_152 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3319_));
INVX1 INVX1_153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3321_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3322_));
INVX1 INVX1_154 ( .A(\key_out[27] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3330_));
INVX1 INVX1_155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3336_));
INVX1 INVX1_156 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3337_));
INVX1 INVX1_157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3339_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3340_));
INVX1 INVX1_158 ( .A(\key_out[28] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3347_));
INVX1 INVX1_159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3354_));
INVX1 INVX1_16 ( .A(start), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n121_));
INVX1 INVX1_160 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3355_));
INVX1 INVX1_161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3357_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3358_));
INVX1 INVX1_162 ( .A(\key_out[29] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3365_));
INVX1 INVX1_163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3372_));
INVX1 INVX1_164 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3373_));
INVX1 INVX1_165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3376_));
INVX1 INVX1_166 ( .A(\key_out[30] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3383_));
INVX1 INVX1_167 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3390_));
INVX1 INVX1_168 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3392_));
INVX1 INVX1_169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3394_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3395_));
INVX1 INVX1_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n126_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n127_));
INVX1 INVX1_170 ( .A(\key_out[31] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3402_));
INVX1 INVX1_171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3409_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3410_));
INVX1 INVX1_172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3413_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3414_));
INVX1 INVX1_173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3415_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3416_));
INVX1 INVX1_174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3418_));
INVX1 INVX1_175 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3419_));
INVX1 INVX1_176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3423_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3424_));
INVX1 INVX1_177 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3425_));
INVX1 INVX1_178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3431_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3432_));
INVX1 INVX1_179 ( .A(AES_CORE_DATAPATH_col_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3433_));
INVX1 INVX1_18 ( .A(AES_CORE_CONTROL_UNIT_rd_count_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n128_));
INVX1 INVX1_180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3437_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3438_));
INVX1 INVX1_181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3439_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3440_));
INVX1 INVX1_182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3449_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3450_));
INVX1 INVX1_183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3452_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3453_));
INVX1 INVX1_184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3456_));
INVX1 INVX1_185 ( .A(AES_CORE_DATAPATH_last_round_pp2), .Y(AES_CORE_DATAPATH__abc_16009_new_n3460_));
INVX1 INVX1_186 ( .A(AES_CORE_DATAPATH_col_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3468_));
INVX1 INVX1_187 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3470_));
INVX1 INVX1_188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3477_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3478_));
INVX1 INVX1_189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3479_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_));
INVX1 INVX1_19 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n142_));
INVX1 INVX1_190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3484_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3485_));
INVX1 INVX1_191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3487_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3488_));
INVX1 INVX1_192 ( .A(AES_CORE_DATAPATH_col_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3500_));
INVX1 INVX1_193 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3502_));
INVX1 INVX1_194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3509_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3510_));
INVX1 INVX1_195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3511_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_));
INVX1 INVX1_196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3516_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3517_));
INVX1 INVX1_197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3519_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3520_));
INVX1 INVX1_198 ( .A(AES_CORE_DATAPATH_col_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3532_));
INVX1 INVX1_199 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3534_));
INVX1 INVX1_2 ( .A(\addr[0] ), .Y(_abc_15574_new_n12_));
INVX1 INVX1_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n79_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n149_));
INVX1 INVX1_200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3541_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3542_));
INVX1 INVX1_201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3543_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_));
INVX1 INVX1_202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3548_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3549_));
INVX1 INVX1_203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3551_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3552_));
INVX1 INVX1_204 ( .A(AES_CORE_DATAPATH_col_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3564_));
INVX1 INVX1_205 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3566_));
INVX1 INVX1_206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3573_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3574_));
INVX1 INVX1_207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3575_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_));
INVX1 INVX1_208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3580_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3581_));
INVX1 INVX1_209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3583_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3584_));
INVX1 INVX1_21 ( .A(AES_CORE_CONTROL_UNIT_state_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n167_));
INVX1 INVX1_210 ( .A(AES_CORE_DATAPATH_col_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3596_));
INVX1 INVX1_211 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3598_));
INVX1 INVX1_212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3605_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3606_));
INVX1 INVX1_213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3607_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_));
INVX1 INVX1_214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3612_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3613_));
INVX1 INVX1_215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3615_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3616_));
INVX1 INVX1_216 ( .A(AES_CORE_DATAPATH_col_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3628_));
INVX1 INVX1_217 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3630_));
INVX1 INVX1_218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3637_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3638_));
INVX1 INVX1_219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3639_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_));
INVX1 INVX1_22 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n168_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n169_));
INVX1 INVX1_220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3644_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3645_));
INVX1 INVX1_221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3647_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3648_));
INVX1 INVX1_222 ( .A(AES_CORE_DATAPATH_col_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3660_));
INVX1 INVX1_223 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3662_));
INVX1 INVX1_224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3669_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3670_));
INVX1 INVX1_225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3671_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_));
INVX1 INVX1_226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3676_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3677_));
INVX1 INVX1_227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3679_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3680_));
INVX1 INVX1_228 ( .A(AES_CORE_DATAPATH_col_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3692_));
INVX1 INVX1_229 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3694_));
INVX1 INVX1_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n174_));
INVX1 INVX1_230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3701_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3702_));
INVX1 INVX1_231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3703_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_));
INVX1 INVX1_232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3708_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3709_));
INVX1 INVX1_233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3711_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3712_));
INVX1 INVX1_234 ( .A(AES_CORE_DATAPATH_col_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3724_));
INVX1 INVX1_235 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3726_));
INVX1 INVX1_236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3733_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3734_));
INVX1 INVX1_237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3735_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_1_));
INVX1 INVX1_238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3740_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3741_));
INVX1 INVX1_239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3743_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3744_));
INVX1 INVX1_24 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n179_));
INVX1 INVX1_240 ( .A(AES_CORE_DATAPATH_col_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3756_));
INVX1 INVX1_241 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3758_));
INVX1 INVX1_242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3765_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3766_));
INVX1 INVX1_243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3767_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_2_));
INVX1 INVX1_244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3772_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3773_));
INVX1 INVX1_245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3775_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3776_));
INVX1 INVX1_246 ( .A(AES_CORE_DATAPATH_col_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3788_));
INVX1 INVX1_247 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3790_));
INVX1 INVX1_248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3797_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3798_));
INVX1 INVX1_249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3799_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_));
INVX1 INVX1_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n182_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n183_));
INVX1 INVX1_250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3804_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3805_));
INVX1 INVX1_251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3807_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3808_));
INVX1 INVX1_252 ( .A(AES_CORE_DATAPATH_col_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3820_));
INVX1 INVX1_253 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3822_));
INVX1 INVX1_254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3829_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3830_));
INVX1 INVX1_255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3831_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_));
INVX1 INVX1_256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3836_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3837_));
INVX1 INVX1_257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3839_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3840_));
INVX1 INVX1_258 ( .A(AES_CORE_DATAPATH_col_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3852_));
INVX1 INVX1_259 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3854_));
INVX1 INVX1_26 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n214_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n215_));
INVX1 INVX1_260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3861_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3862_));
INVX1 INVX1_261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3863_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_));
INVX1 INVX1_262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3868_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3869_));
INVX1 INVX1_263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3871_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3872_));
INVX1 INVX1_264 ( .A(AES_CORE_DATAPATH_col_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3884_));
INVX1 INVX1_265 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3886_));
INVX1 INVX1_266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3893_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3894_));
INVX1 INVX1_267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3895_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_));
INVX1 INVX1_268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3900_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3901_));
INVX1 INVX1_269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3903_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3904_));
INVX1 INVX1_27 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n199_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n216_));
INVX1 INVX1_270 ( .A(AES_CORE_DATAPATH_col_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3916_));
INVX1 INVX1_271 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3918_));
INVX1 INVX1_272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3925_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3926_));
INVX1 INVX1_273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3927_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_));
INVX1 INVX1_274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3932_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3933_));
INVX1 INVX1_275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3935_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3936_));
INVX1 INVX1_276 ( .A(AES_CORE_DATAPATH_col_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3948_));
INVX1 INVX1_277 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3950_));
INVX1 INVX1_278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3957_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3958_));
INVX1 INVX1_279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3959_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_));
INVX1 INVX1_28 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n228_));
INVX1 INVX1_280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3964_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3965_));
INVX1 INVX1_281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3967_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3968_));
INVX1 INVX1_282 ( .A(AES_CORE_DATAPATH_col_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3980_));
INVX1 INVX1_283 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3982_));
INVX1 INVX1_284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3989_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3990_));
INVX1 INVX1_285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3991_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_1_));
INVX1 INVX1_286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3997_));
INVX1 INVX1_287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3999_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4000_));
INVX1 INVX1_288 ( .A(AES_CORE_DATAPATH_col_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4012_));
INVX1 INVX1_289 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4014_));
INVX1 INVX1_29 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n191_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n229_));
INVX1 INVX1_290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4021_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4022_));
INVX1 INVX1_291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4023_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_2_));
INVX1 INVX1_292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4028_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4029_));
INVX1 INVX1_293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4032_));
INVX1 INVX1_294 ( .A(AES_CORE_DATAPATH_col_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4044_));
INVX1 INVX1_295 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4046_));
INVX1 INVX1_296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4053_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4054_));
INVX1 INVX1_297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4055_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_));
INVX1 INVX1_298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4060_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4061_));
INVX1 INVX1_299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4063_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4064_));
INVX1 INVX1_3 ( .A(\aes_mode[1] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_));
INVX1 INVX1_30 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n138_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n231_));
INVX1 INVX1_300 ( .A(AES_CORE_DATAPATH_col_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4076_));
INVX1 INVX1_301 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4078_));
INVX1 INVX1_302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4085_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4086_));
INVX1 INVX1_303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4087_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_));
INVX1 INVX1_304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4092_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4093_));
INVX1 INVX1_305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4095_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4096_));
INVX1 INVX1_306 ( .A(AES_CORE_DATAPATH_col_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4108_));
INVX1 INVX1_307 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4110_));
INVX1 INVX1_308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4118_));
INVX1 INVX1_309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4119_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_));
INVX1 INVX1_31 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n232_));
INVX1 INVX1_310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4125_));
INVX1 INVX1_311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4128_));
INVX1 INVX1_312 ( .A(AES_CORE_DATAPATH_col_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4140_));
INVX1 INVX1_313 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4142_));
INVX1 INVX1_314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4149_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4150_));
INVX1 INVX1_315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4151_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_));
INVX1 INVX1_316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4156_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4157_));
INVX1 INVX1_317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4159_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4160_));
INVX1 INVX1_318 ( .A(AES_CORE_DATAPATH_col_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4172_));
INVX1 INVX1_319 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4174_));
INVX1 INVX1_32 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n130_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n257_));
INVX1 INVX1_320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4181_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4182_));
INVX1 INVX1_321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4183_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_));
INVX1 INVX1_322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4188_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4189_));
INVX1 INVX1_323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4191_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4192_));
INVX1 INVX1_324 ( .A(AES_CORE_DATAPATH_col_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4204_));
INVX1 INVX1_325 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4206_));
INVX1 INVX1_326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4213_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4214_));
INVX1 INVX1_327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4215_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_));
INVX1 INVX1_328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4220_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4221_));
INVX1 INVX1_329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4223_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4224_));
INVX1 INVX1_33 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_DATAPATH__abc_16009_new_n2457_));
INVX1 INVX1_330 ( .A(AES_CORE_DATAPATH_col_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4236_));
INVX1 INVX1_331 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4238_));
INVX1 INVX1_332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4245_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4246_));
INVX1 INVX1_333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4247_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_1_));
INVX1 INVX1_334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4252_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4253_));
INVX1 INVX1_335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4255_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4256_));
INVX1 INVX1_336 ( .A(AES_CORE_DATAPATH_col_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4268_));
INVX1 INVX1_337 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4270_));
INVX1 INVX1_338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4277_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4278_));
INVX1 INVX1_339 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4279_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_2_));
INVX1 INVX1_34 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2467_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2475_));
INVX1 INVX1_340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4284_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4285_));
INVX1 INVX1_341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4287_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4288_));
INVX1 INVX1_342 ( .A(AES_CORE_DATAPATH_col_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4300_));
INVX1 INVX1_343 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4302_));
INVX1 INVX1_344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4310_));
INVX1 INVX1_345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4311_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_));
INVX1 INVX1_346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4316_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4317_));
INVX1 INVX1_347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4319_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4320_));
INVX1 INVX1_348 ( .A(AES_CORE_DATAPATH_col_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4332_));
INVX1 INVX1_349 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4334_));
INVX1 INVX1_35 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2483_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2484_));
INVX1 INVX1_350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4341_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4342_));
INVX1 INVX1_351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_));
INVX1 INVX1_352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4348_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4349_));
INVX1 INVX1_353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4351_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4352_));
INVX1 INVX1_354 ( .A(AES_CORE_DATAPATH_col_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4364_));
INVX1 INVX1_355 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4366_));
INVX1 INVX1_356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4373_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4374_));
INVX1 INVX1_357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_));
INVX1 INVX1_358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4380_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4381_));
INVX1 INVX1_359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4383_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4384_));
INVX1 INVX1_36 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2485_));
INVX1 INVX1_360 ( .A(AES_CORE_DATAPATH_col_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4396_));
INVX1 INVX1_361 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4398_));
INVX1 INVX1_362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4405_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4406_));
INVX1 INVX1_363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4407_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_));
INVX1 INVX1_364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4412_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4413_));
INVX1 INVX1_365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4415_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4416_));
INVX1 INVX1_366 ( .A(AES_CORE_DATAPATH_col_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4428_));
INVX1 INVX1_367 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_in_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4430_));
INVX1 INVX1_368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4437_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4438_));
INVX1 INVX1_369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4439_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_));
INVX1 INVX1_37 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .Y(AES_CORE_DATAPATH__abc_16009_new_n2801_));
INVX1 INVX1_370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4444_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4445_));
INVX1 INVX1_371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4447_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4448_));
INVX1 INVX1_372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4559_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4560_));
INVX1 INVX1_373 ( .A(start), .Y(AES_CORE_DATAPATH__abc_16009_new_n4561_));
INVX1 INVX1_374 ( .A(\key_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4562_));
INVX1 INVX1_375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4572_));
INVX1 INVX1_376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4576_));
INVX1 INVX1_377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4860_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4861_));
INVX1 INVX1_378 ( .A(\key_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n4862_));
INVX1 INVX1_379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4865_));
INVX1 INVX1_38 ( .A(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_16009_new_n2802_));
INVX1 INVX1_380 ( .A(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5155_));
INVX1 INVX1_381 ( .A(\key_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5253_));
INVX1 INVX1_382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5542_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5543_));
INVX1 INVX1_383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5550_));
INVX1 INVX1_384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5739_));
INVX1 INVX1_385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5743_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5744_));
INVX1 INVX1_386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5747_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5748_));
INVX1 INVX1_387 ( .A(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n5757_));
INVX1 INVX1_388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5759_));
INVX1 INVX1_389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5764_));
INVX1 INVX1_39 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2806_));
INVX1 INVX1_390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3454_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5779_));
INVX1 INVX1_391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3463_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5782_));
INVX1 INVX1_392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5761_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5785_));
INVX1 INVX1_393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5787_));
INVX1 INVX1_394 ( .A(AES_CORE_CONTROL_UNIT_mode_cbc), .Y(AES_CORE_DATAPATH__abc_16009_new_n5792_));
INVX1 INVX1_395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5798_));
INVX1 INVX1_396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3489_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5816_));
INVX1 INVX1_397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3495_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5819_));
INVX1 INVX1_398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5823_));
INVX1 INVX1_399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5837_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5838_));
INVX1 INVX1_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n74_), .Y(AES_CORE_CONTROL_UNIT_mode_ctr));
INVX1 INVX1_40 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n2807_));
INVX1 INVX1_400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3521_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5883_));
INVX1 INVX1_401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3527_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5886_));
INVX1 INVX1_402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5889_));
INVX1 INVX1_403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5881_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5891_));
INVX1 INVX1_404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3553_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5916_));
INVX1 INVX1_405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3559_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5919_));
INVX1 INVX1_406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5923_));
INVX1 INVX1_407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5938_));
INVX1 INVX1_408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3585_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5983_));
INVX1 INVX1_409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3591_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5986_));
INVX1 INVX1_41 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2824_));
INVX1 INVX1_410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5967_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5989_));
INVX1 INVX1_411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5981_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5991_));
INVX1 INVX1_412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3617_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6033_));
INVX1 INVX1_413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3623_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6036_));
INVX1 INVX1_414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6017_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6039_));
INVX1 INVX1_415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6041_));
INVX1 INVX1_416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3649_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6083_));
INVX1 INVX1_417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3655_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6086_));
INVX1 INVX1_418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6067_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6089_));
INVX1 INVX1_419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6081_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6091_));
INVX1 INVX1_42 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2826_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2827_));
INVX1 INVX1_420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3681_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6116_));
INVX1 INVX1_421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6119_));
INVX1 INVX1_422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6123_));
INVX1 INVX1_423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6137_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6138_));
INVX1 INVX1_424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3713_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6183_));
INVX1 INVX1_425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3719_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6186_));
INVX1 INVX1_426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6167_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6189_));
INVX1 INVX1_427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6181_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6191_));
INVX1 INVX1_428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3745_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6216_));
INVX1 INVX1_429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3751_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6219_));
INVX1 INVX1_43 ( .A(AES_CORE_DATAPATH_key_out_sel_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2830_));
INVX1 INVX1_430 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6222_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6223_));
INVX1 INVX1_431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6237_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6238_));
INVX1 INVX1_432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6283_));
INVX1 INVX1_433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3783_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6286_));
INVX1 INVX1_434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6267_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6289_));
INVX1 INVX1_435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6281_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6291_));
INVX1 INVX1_436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3809_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6316_));
INVX1 INVX1_437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3815_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6319_));
INVX1 INVX1_438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6322_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6323_));
INVX1 INVX1_439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6337_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6338_));
INVX1 INVX1_44 ( .A(AES_CORE_DATAPATH_key_out_sel_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2832_));
INVX1 INVX1_440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3841_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6383_));
INVX1 INVX1_441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3847_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6386_));
INVX1 INVX1_442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6389_));
INVX1 INVX1_443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6381_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6391_));
INVX1 INVX1_444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3873_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6416_));
INVX1 INVX1_445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3879_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6419_));
INVX1 INVX1_446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6422_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6423_));
INVX1 INVX1_447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6437_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6438_));
INVX1 INVX1_448 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3905_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6483_));
INVX1 INVX1_449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3911_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6486_));
INVX1 INVX1_45 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2836_));
INVX1 INVX1_450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6467_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6489_));
INVX1 INVX1_451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6481_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6491_));
INVX1 INVX1_452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6516_));
INVX1 INVX1_453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3943_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6519_));
INVX1 INVX1_454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6522_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6523_));
INVX1 INVX1_455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6537_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6538_));
INVX1 INVX1_456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3969_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6583_));
INVX1 INVX1_457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3975_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6586_));
INVX1 INVX1_458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6567_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6589_));
INVX1 INVX1_459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6581_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6591_));
INVX1 INVX1_46 ( .A(\key_out[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2844_));
INVX1 INVX1_460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4001_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6616_));
INVX1 INVX1_461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4007_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6619_));
INVX1 INVX1_462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6622_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6623_));
INVX1 INVX1_463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6637_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6638_));
INVX1 INVX1_464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4033_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6666_));
INVX1 INVX1_465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4039_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6669_));
INVX1 INVX1_466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6672_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6673_));
INVX1 INVX1_467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6688_));
INVX1 INVX1_468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4065_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6716_));
INVX1 INVX1_469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4071_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6719_));
INVX1 INVX1_47 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2850_));
INVX1 INVX1_470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6722_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6723_));
INVX1 INVX1_471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6737_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6738_));
INVX1 INVX1_472 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4097_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6783_));
INVX1 INVX1_473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6786_));
INVX1 INVX1_474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6767_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6789_));
INVX1 INVX1_475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6781_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6791_));
INVX1 INVX1_476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4129_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6816_));
INVX1 INVX1_477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4135_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6819_));
INVX1 INVX1_478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6823_));
INVX1 INVX1_479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6837_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6838_));
INVX1 INVX1_48 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2851_));
INVX1 INVX1_480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4161_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6883_));
INVX1 INVX1_481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4167_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6886_));
INVX1 INVX1_482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6889_));
INVX1 INVX1_483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6881_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6891_));
INVX1 INVX1_484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4193_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6916_));
INVX1 INVX1_485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4199_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6919_));
INVX1 INVX1_486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6923_));
INVX1 INVX1_487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6938_));
INVX1 INVX1_488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4225_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6983_));
INVX1 INVX1_489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6986_));
INVX1 INVX1_49 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2853_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2854_));
INVX1 INVX1_490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6967_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6989_));
INVX1 INVX1_491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6981_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6991_));
INVX1 INVX1_492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4257_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7016_));
INVX1 INVX1_493 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4263_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7019_));
INVX1 INVX1_494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7022_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7023_));
INVX1 INVX1_495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7037_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7038_));
INVX1 INVX1_496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4289_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7066_));
INVX1 INVX1_497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4295_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7069_));
INVX1 INVX1_498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7072_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7073_));
INVX1 INVX1_499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7087_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7088_));
INVX1 INVX1_5 ( .A(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n77_));
INVX1 INVX1_50 ( .A(\key_out[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2862_));
INVX1 INVX1_500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4321_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7133_));
INVX1 INVX1_501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4327_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7136_));
INVX1 INVX1_502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7139_));
INVX1 INVX1_503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7131_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7141_));
INVX1 INVX1_504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4353_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7166_));
INVX1 INVX1_505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4359_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7169_));
INVX1 INVX1_506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7172_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7173_));
INVX1 INVX1_507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7187_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7188_));
INVX1 INVX1_508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4385_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7233_));
INVX1 INVX1_509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4391_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7236_));
INVX1 INVX1_51 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2868_));
INVX1 INVX1_510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7217_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7239_));
INVX1 INVX1_511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7241_));
INVX1 INVX1_512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7283_));
INVX1 INVX1_513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4423_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7286_));
INVX1 INVX1_514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7267_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7289_));
INVX1 INVX1_515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7281_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7291_));
INVX1 INVX1_516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4449_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7316_));
INVX1 INVX1_517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7319_));
INVX1 INVX1_518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7322_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7323_));
INVX1 INVX1_519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7337_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7338_));
INVX1 INVX1_52 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2869_));
INVX1 INVX1_520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7363_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7364_));
INVX1 INVX1_521 ( .A(\key_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n7365_));
INVX1 INVX1_522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7375_));
INVX1 INVX1_523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2482_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7753_));
INVX1 INVX1_524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2466_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8010_));
INVX1 INVX1_525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8267_));
INVX1 INVX1_526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8524_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8525_));
INVX1 INVX1_527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8531_));
INVX1 INVX1_528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8628_));
INVX1 INVX1_529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8918_));
INVX1 INVX1_53 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2871_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2872_));
INVX1 INVX1_530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8920_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8921_));
INVX1 INVX1_531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8925_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8926_));
INVX1 INVX1_532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8934_));
INVX1 INVX1_533 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8937_));
INVX1 INVX1_534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8948_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8949_));
INVX1 INVX1_535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8960_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8961_));
INVX1 INVX1_536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8970_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8971_));
INVX1 INVX1_537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8978_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8979_));
INVX1 INVX1_538 ( .A(AES_CORE_DATAPATH_iv_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8990_));
INVX1 INVX1_539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8999_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9000_));
INVX1 INVX1_54 ( .A(\key_out[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2880_));
INVX1 INVX1_540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9009_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9010_));
INVX1 INVX1_541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9022_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9023_));
INVX1 INVX1_542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9033_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9034_));
INVX1 INVX1_543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9046_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9047_));
INVX1 INVX1_544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9056_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9057_));
INVX1 INVX1_545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9068_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9069_));
INVX1 INVX1_546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9080_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9081_));
INVX1 INVX1_547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9092_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9093_));
INVX1 INVX1_548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9104_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9105_));
INVX1 INVX1_549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9116_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9117_));
INVX1 INVX1_55 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2886_));
INVX1 INVX1_550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9130_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9131_));
INVX1 INVX1_551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9141_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9142_));
INVX1 INVX1_552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9156_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9157_));
INVX1 INVX1_553 ( .A(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9168_));
INVX1 INVX1_554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9183_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9184_));
INVX1 INVX1_555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9194_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9195_));
INVX1 INVX1_556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9209_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9210_));
INVX1 INVX1_557 ( .A(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9221_));
INVX1 INVX1_558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9234_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9235_));
INVX1 INVX1_559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9246_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9247_));
INVX1 INVX1_56 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2888_));
INVX1 INVX1_560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9258_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9259_));
INVX1 INVX1_561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9270_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9271_));
INVX1 INVX1_562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9281_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9282_));
INVX1 INVX1_563 ( .A(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9294_));
INVX1 INVX1_564 ( .A(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9305_));
INVX1 INVX1_565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9404_));
INVX1 INVX1_566 ( .A(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9758_));
INVX1 INVX1_567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9857_));
INVX1 INVX1_568 ( .A(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10211_));
INVX1 INVX1_569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10310_));
INVX1 INVX1_57 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2890_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2891_));
INVX1 INVX1_570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3443_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_));
INVX1 INVX1_571 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n327_));
INVX1 INVX1_572 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n329_));
INVX1 INVX1_573 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n331_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n332_));
INVX1 INVX1_574 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n333_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n335_));
INVX1 INVX1_575 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n338_));
INVX1 INVX1_576 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n340_));
INVX1 INVX1_577 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n342_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n343_));
INVX1 INVX1_578 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n344_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n346_));
INVX1 INVX1_579 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n349_));
INVX1 INVX1_58 ( .A(\key_out[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2898_));
INVX1 INVX1_580 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n351_));
INVX1 INVX1_581 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n353_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n354_));
INVX1 INVX1_582 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n355_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n357_));
INVX1 INVX1_583 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n360_));
INVX1 INVX1_584 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n362_));
INVX1 INVX1_585 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n364_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n365_));
INVX1 INVX1_586 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n366_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n368_));
INVX1 INVX1_587 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n371_));
INVX1 INVX1_588 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n373_));
INVX1 INVX1_589 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n375_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n376_));
INVX1 INVX1_59 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2904_));
INVX1 INVX1_590 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n377_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n379_));
INVX1 INVX1_591 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n382_));
INVX1 INVX1_592 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n384_));
INVX1 INVX1_593 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n386_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n387_));
INVX1 INVX1_594 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n388_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n390_));
INVX1 INVX1_595 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n393_));
INVX1 INVX1_596 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n395_));
INVX1 INVX1_597 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n397_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n398_));
INVX1 INVX1_598 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n399_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n401_));
INVX1 INVX1_599 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n404_));
INVX1 INVX1_6 ( .A(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n78_));
INVX1 INVX1_60 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2906_));
INVX1 INVX1_600 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n406_));
INVX1 INVX1_601 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n408_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n409_));
INVX1 INVX1_602 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n410_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n412_));
INVX1 INVX1_603 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n415_));
INVX1 INVX1_604 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n417_));
INVX1 INVX1_605 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n419_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n420_));
INVX1 INVX1_606 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n421_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n423_));
INVX1 INVX1_607 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n426_));
INVX1 INVX1_608 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n428_));
INVX1 INVX1_609 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n430_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n431_));
INVX1 INVX1_61 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2908_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2909_));
INVX1 INVX1_610 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n432_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n434_));
INVX1 INVX1_611 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n437_));
INVX1 INVX1_612 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n439_));
INVX1 INVX1_613 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n441_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n442_));
INVX1 INVX1_614 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n443_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n445_));
INVX1 INVX1_615 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n448_));
INVX1 INVX1_616 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n450_));
INVX1 INVX1_617 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n452_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n453_));
INVX1 INVX1_618 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n454_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n456_));
INVX1 INVX1_619 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n459_));
INVX1 INVX1_62 ( .A(\key_out[4] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2916_));
INVX1 INVX1_620 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n461_));
INVX1 INVX1_621 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n463_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n464_));
INVX1 INVX1_622 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n465_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n467_));
INVX1 INVX1_623 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n470_));
INVX1 INVX1_624 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n472_));
INVX1 INVX1_625 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n474_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n475_));
INVX1 INVX1_626 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n476_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n478_));
INVX1 INVX1_627 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n481_));
INVX1 INVX1_628 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n483_));
INVX1 INVX1_629 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n485_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n486_));
INVX1 INVX1_63 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2922_));
INVX1 INVX1_630 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n487_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n489_));
INVX1 INVX1_631 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n492_));
INVX1 INVX1_632 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n494_));
INVX1 INVX1_633 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n496_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n497_));
INVX1 INVX1_634 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n498_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n500_));
INVX1 INVX1_635 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n503_));
INVX1 INVX1_636 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n505_));
INVX1 INVX1_637 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n507_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n508_));
INVX1 INVX1_638 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n509_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n511_));
INVX1 INVX1_639 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n514_));
INVX1 INVX1_64 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2923_));
INVX1 INVX1_640 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n516_));
INVX1 INVX1_641 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n518_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n519_));
INVX1 INVX1_642 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n520_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n522_));
INVX1 INVX1_643 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n525_));
INVX1 INVX1_644 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n527_));
INVX1 INVX1_645 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n529_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n530_));
INVX1 INVX1_646 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n531_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n533_));
INVX1 INVX1_647 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n536_));
INVX1 INVX1_648 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n538_));
INVX1 INVX1_649 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n540_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n541_));
INVX1 INVX1_65 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2925_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2926_));
INVX1 INVX1_650 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n542_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n544_));
INVX1 INVX1_651 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n547_));
INVX1 INVX1_652 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n549_));
INVX1 INVX1_653 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n551_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n552_));
INVX1 INVX1_654 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n553_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n555_));
INVX1 INVX1_655 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n558_));
INVX1 INVX1_656 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n560_));
INVX1 INVX1_657 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n562_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n563_));
INVX1 INVX1_658 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n564_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n566_));
INVX1 INVX1_659 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n569_));
INVX1 INVX1_66 ( .A(\key_out[5] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2934_));
INVX1 INVX1_660 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n571_));
INVX1 INVX1_661 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n573_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n574_));
INVX1 INVX1_662 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n575_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n577_));
INVX1 INVX1_663 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n580_));
INVX1 INVX1_664 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n582_));
INVX1 INVX1_665 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n584_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n585_));
INVX1 INVX1_666 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n586_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n588_));
INVX1 INVX1_667 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n592_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n593_));
INVX1 INVX1_668 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n595_));
INVX1 INVX1_669 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n596_));
INVX1 INVX1_67 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2940_));
INVX1 INVX1_670 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_));
INVX1 INVX1_671 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n600_));
INVX1 INVX1_672 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n603_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n604_));
INVX1 INVX1_673 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n606_));
INVX1 INVX1_674 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n608_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n609_));
INVX1 INVX1_675 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n610_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n611_));
INVX1 INVX1_676 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n594_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n613_));
INVX1 INVX1_677 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n617_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n618_));
INVX1 INVX1_678 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n619_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n620_));
INVX1 INVX1_679 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n621_));
INVX1 INVX1_68 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2942_));
INVX1 INVX1_680 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n624_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n625_));
INVX1 INVX1_681 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n637_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n638_));
INVX1 INVX1_682 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_add_w_out), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_));
INVX1 INVX1_683 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n636_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n643_));
INVX1 INVX1_684 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n649_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n650_));
INVX1 INVX1_685 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n651_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n652_));
INVX1 INVX1_686 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n653_));
INVX1 INVX1_687 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n655_));
INVX1 INVX1_688 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n657_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n658_));
INVX1 INVX1_689 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n664_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n665_));
INVX1 INVX1_69 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2944_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2945_));
INVX1 INVX1_690 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n601_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n676_));
INVX1 INVX1_691 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n693_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n694_));
INVX1 INVX1_692 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n695_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n696_));
INVX1 INVX1_693 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n702_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n703_));
INVX1 INVX1_694 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n704_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n708_));
INVX1 INVX1_695 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n714_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n715_));
INVX1 INVX1_696 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n717_));
INVX1 INVX1_697 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n718_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n719_));
INVX1 INVX1_698 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n721_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n722_));
INVX1 INVX1_699 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n724_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n725_));
INVX1 INVX1_7 ( .A(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n80_));
INVX1 INVX1_70 ( .A(\key_out[6] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2952_));
INVX1 INVX1_700 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n729_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n730_));
INVX1 INVX1_701 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n716_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n732_));
INVX1 INVX1_702 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n736_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n737_));
INVX1 INVX1_703 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n738_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n739_));
INVX1 INVX1_704 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n740_));
INVX1 INVX1_705 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n760_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n761_));
INVX1 INVX1_706 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n762_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n763_));
INVX1 INVX1_707 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n767_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n768_));
INVX1 INVX1_708 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n771_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n773_));
INVX1 INVX1_709 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n777_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n778_));
INVX1 INVX1_71 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2958_));
INVX1 INVX1_710 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n779_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n780_));
INVX1 INVX1_711 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n783_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n784_));
INVX1 INVX1_712 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n785_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n786_));
INVX1 INVX1_713 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n787_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n791_));
INVX1 INVX1_714 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n797_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n798_));
INVX1 INVX1_715 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n804_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n805_));
INVX1 INVX1_716 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n811_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n812_));
INVX1 INVX1_717 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n818_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n819_));
INVX1 INVX1_718 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n825_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n826_));
INVX1 INVX1_719 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n832_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n833_));
INVX1 INVX1_72 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2959_));
INVX1 INVX1_720 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n839_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n840_));
INVX1 INVX1_721 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n846_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n847_));
INVX1 INVX1_722 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n853_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n854_));
INVX1 INVX1_723 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n860_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n861_));
INVX1 INVX1_724 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n867_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n868_));
INVX1 INVX1_725 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n874_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n875_));
INVX1 INVX1_726 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n881_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n882_));
INVX1 INVX1_727 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n888_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n889_));
INVX1 INVX1_728 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n895_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n896_));
INVX1 INVX1_729 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n902_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n903_));
INVX1 INVX1_73 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2961_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2962_));
INVX1 INVX1_730 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n909_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n910_));
INVX1 INVX1_731 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n916_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n917_));
INVX1 INVX1_732 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n923_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n924_));
INVX1 INVX1_733 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n930_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n931_));
INVX1 INVX1_734 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n937_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n938_));
INVX1 INVX1_735 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n944_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n945_));
INVX1 INVX1_736 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n951_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n952_));
INVX1 INVX1_737 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n958_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n959_));
INVX1 INVX1_738 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n965_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n966_));
INVX1 INVX1_739 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n972_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n973_));
INVX1 INVX1_74 ( .A(\key_out[7] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2970_));
INVX1 INVX1_740 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n979_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n980_));
INVX1 INVX1_741 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n986_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n987_));
INVX1 INVX1_742 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n993_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n994_));
INVX1 INVX1_743 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1000_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1001_));
INVX1 INVX1_744 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1007_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1008_));
INVX1 INVX1_745 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1014_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1015_));
INVX1 INVX1_746 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1021_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1022_));
INVX1 INVX1_747 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1025_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1026_));
INVX1 INVX1_748 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1029_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1030_));
INVX1 INVX1_749 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1033_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1034_));
INVX1 INVX1_75 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2976_));
INVX1 INVX1_750 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1037_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1038_));
INVX1 INVX1_751 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1041_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1042_));
INVX1 INVX1_752 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1045_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1046_));
INVX1 INVX1_753 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1049_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1050_));
INVX1 INVX1_754 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1053_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1054_));
INVX1 INVX1_755 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1057_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1058_));
INVX1 INVX1_756 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1061_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1062_));
INVX1 INVX1_757 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1065_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1066_));
INVX1 INVX1_758 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1069_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1070_));
INVX1 INVX1_759 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1073_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1074_));
INVX1 INVX1_76 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2977_));
INVX1 INVX1_760 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1077_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1078_));
INVX1 INVX1_761 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1081_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1082_));
INVX1 INVX1_762 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1085_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1086_));
INVX1 INVX1_763 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1089_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1090_));
INVX1 INVX1_764 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1093_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1094_));
INVX1 INVX1_765 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1097_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1098_));
INVX1 INVX1_766 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1101_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1102_));
INVX1 INVX1_767 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1105_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1106_));
INVX1 INVX1_768 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1109_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1110_));
INVX1 INVX1_769 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1113_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1114_));
INVX1 INVX1_77 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2979_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2980_));
INVX1 INVX1_770 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1116_));
INVX1 INVX1_771 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1120_));
INVX1 INVX1_772 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1124_));
INVX1 INVX1_773 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1128_));
INVX1 INVX1_774 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1132_));
INVX1 INVX1_775 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n728_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1134_));
INVX1 INVX1_776 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1137_));
INVX1 INVX1_777 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1142_));
INVX1 INVX1_778 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n770_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1143_));
INVX1 INVX1_779 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1147_));
INVX1 INVX1_78 ( .A(\key_out[8] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2987_));
INVX1 INVX1_780 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1151_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1152_));
INVX1 INVX1_781 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1155_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1156_));
INVX1 INVX1_782 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1159_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1160_));
INVX1 INVX1_783 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1163_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1164_));
INVX1 INVX1_784 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1167_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1168_));
INVX1 INVX1_785 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1171_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1172_));
INVX1 INVX1_786 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1175_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1176_));
INVX1 INVX1_787 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1179_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1180_));
INVX1 INVX1_788 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1183_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1184_));
INVX1 INVX1_789 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1187_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1188_));
INVX1 INVX1_79 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2994_));
INVX1 INVX1_790 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1191_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1192_));
INVX1 INVX1_791 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1195_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1196_));
INVX1 INVX1_792 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1199_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1200_));
INVX1 INVX1_793 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1203_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1204_));
INVX1 INVX1_794 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1207_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1208_));
INVX1 INVX1_795 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1211_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1212_));
INVX1 INVX1_796 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1215_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1216_));
INVX1 INVX1_797 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1219_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1220_));
INVX1 INVX1_798 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1223_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1224_));
INVX1 INVX1_799 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1227_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1228_));
INVX1 INVX1_8 ( .A(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n81_));
INVX1 INVX1_80 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2995_));
INVX1 INVX1_800 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1231_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1232_));
INVX1 INVX1_801 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1235_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1236_));
INVX1 INVX1_802 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1239_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1240_));
INVX1 INVX1_803 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1243_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1244_));
INVX1 INVX1_804 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1247_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1248_));
INVX1 INVX1_805 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1251_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1252_));
INVX1 INVX1_806 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1255_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1256_));
INVX1 INVX1_807 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1259_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1260_));
INVX1 INVX1_808 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1263_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1264_));
INVX1 INVX1_809 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1267_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1268_));
INVX1 INVX1_81 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2997_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2998_));
INVX1 INVX1_810 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1271_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1272_));
INVX1 INVX1_811 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1275_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1276_));
INVX1 INVX1_812 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n97_));
INVX1 INVX1_813 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n98_));
INVX1 INVX1_814 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n102_));
INVX1 INVX1_815 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n104_));
INVX1 INVX1_816 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n106_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_));
INVX1 INVX1_817 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n109_));
INVX1 INVX1_818 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n100_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n114_));
INVX1 INVX1_819 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n111_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n116_));
INVX1 INVX1_82 ( .A(\key_out[9] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3006_));
INVX1 INVX1_820 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n119_));
INVX1 INVX1_821 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n120_));
INVX1 INVX1_822 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n121_));
INVX1 INVX1_823 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n126_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n127_));
INVX1 INVX1_824 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n130_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n131_));
INVX1 INVX1_825 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n134_));
INVX1 INVX1_826 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_));
INVX1 INVX1_827 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n138_));
INVX1 INVX1_828 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n139_));
INVX1 INVX1_829 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n123_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n146_));
INVX1 INVX1_83 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3012_));
INVX1 INVX1_830 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_));
INVX1 INVX1_831 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n163_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n164_));
INVX1 INVX1_832 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n166_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n167_));
INVX1 INVX1_833 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n169_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n170_));
INVX1 INVX1_834 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n173_));
INVX1 INVX1_835 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n174_));
INVX1 INVX1_836 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_));
INVX1 INVX1_837 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n179_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n180_));
INVX1 INVX1_838 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n183_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_));
INVX1 INVX1_839 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n186_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n187_));
INVX1 INVX1_84 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3013_));
INVX1 INVX1_840 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_));
INVX1 INVX1_841 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_));
INVX1 INVX1_842 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n196_));
INVX1 INVX1_843 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n198_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n202_));
INVX1 INVX1_844 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n222_));
INVX1 INVX1_845 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n225_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n226_));
INVX1 INVX1_846 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n228_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n229_));
INVX1 INVX1_847 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_));
INVX1 INVX1_848 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n232_));
INVX1 INVX1_849 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n234_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n235_));
INVX1 INVX1_85 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3015_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3016_));
INVX1 INVX1_850 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n240_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n241_));
INVX1 INVX1_851 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n248_));
INVX1 INVX1_852 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n250_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n254_));
INVX1 INVX1_853 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n263_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n264_));
INVX1 INVX1_854 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n270_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n271_));
INVX1 INVX1_855 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n273_));
INVX1 INVX1_856 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n277_));
INVX1 INVX1_857 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n280_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n281_));
INVX1 INVX1_858 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n283_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n284_));
INVX1 INVX1_859 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_));
INVX1 INVX1_86 ( .A(\key_out[10] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3023_));
INVX1 INVX1_860 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n287_));
INVX1 INVX1_861 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n291_));
INVX1 INVX1_862 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n289_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n292_));
INVX1 INVX1_863 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n294_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n295_));
INVX1 INVX1_864 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n298_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_));
INVX1 INVX1_865 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n316_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n317_));
INVX1 INVX1_866 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n340_));
INVX1 INVX1_867 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n343_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n344_));
INVX1 INVX1_868 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n346_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n347_));
INVX1 INVX1_869 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n348_));
INVX1 INVX1_87 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3030_));
INVX1 INVX1_870 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n350_));
INVX1 INVX1_871 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n353_));
INVX1 INVX1_872 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n355_));
INVX1 INVX1_873 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n357_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n358_));
INVX1 INVX1_874 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n361_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_));
INVX1 INVX1_875 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n364_));
INVX1 INVX1_876 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n366_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n368_));
INVX1 INVX1_877 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n403_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n404_));
INVX1 INVX1_878 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n405_));
INVX1 INVX1_879 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n408_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n409_));
INVX1 INVX1_88 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3031_));
INVX1 INVX1_880 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n412_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_));
INVX1 INVX1_881 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n415_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n416_));
INVX1 INVX1_882 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n417_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n418_));
INVX1 INVX1_883 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n421_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n432_));
INVX1 INVX1_884 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n447_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n448_));
INVX1 INVX1_885 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n450_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n455_));
INVX1 INVX1_886 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n453_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n456_));
INVX1 INVX1_887 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n459_));
INVX1 INVX1_888 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n465_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n466_));
INVX1 INVX1_889 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n471_));
INVX1 INVX1_89 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3033_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3034_));
INVX1 INVX1_890 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n469_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n472_));
INVX1 INVX1_891 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n474_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n475_));
INVX1 INVX1_892 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n481_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n482_));
INVX1 INVX1_893 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n485_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n487_));
INVX1 INVX1_894 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n490_));
INVX1 INVX1_895 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n493_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n494_));
INVX1 INVX1_896 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n497_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n499_));
INVX1 INVX1_897 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n507_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n508_));
INVX1 INVX1_898 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_));
INVX1 INVX1_899 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_8_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n513_));
INVX1 INVX1_9 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .Y(AES_CORE_CONTROL_UNIT_encrypt_decrypt));
INVX1 INVX1_90 ( .A(\key_out[11] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3042_));
INVX1 INVX1_900 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n516_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n517_));
INVX1 INVX1_901 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n523_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n524_));
INVX1 INVX1_902 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n530_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n531_));
INVX1 INVX1_903 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n532_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n533_));
INVX1 INVX1_904 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n535_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_9_));
INVX1 INVX1_905 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n539_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n541_));
INVX1 INVX1_906 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n549_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n550_));
INVX1 INVX1_907 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n546_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n552_));
INVX1 INVX1_908 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n555_));
INVX1 INVX1_909 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n558_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n560_));
INVX1 INVX1_91 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3048_));
INVX1 INVX1_910 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n565_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n566_));
INVX1 INVX1_911 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n569_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n570_));
INVX1 INVX1_912 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n573_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n574_));
INVX1 INVX1_913 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n582_));
INVX1 INVX1_914 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n590_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n591_));
INVX1 INVX1_915 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n594_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n595_));
INVX1 INVX1_916 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n598_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n599_));
INVX1 INVX1_917 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n607_));
INVX1 INVX1_918 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n618_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n619_));
INVX1 INVX1_919 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n615_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n621_));
INVX1 INVX1_92 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3049_));
INVX1 INVX1_920 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n624_));
INVX1 INVX1_921 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n636_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n637_));
INVX1 INVX1_922 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n640_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n641_));
INVX1 INVX1_923 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n644_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_));
INVX1 INVX1_924 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n648_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n650_));
INVX1 INVX1_925 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n658_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_));
INVX1 INVX1_926 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n662_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n663_));
INVX1 INVX1_927 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n655_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n665_));
INVX1 INVX1_928 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n667_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_));
INVX1 INVX1_929 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n671_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n673_));
INVX1 INVX1_93 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3051_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3052_));
INVX1 INVX1_930 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n681_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n682_));
INVX1 INVX1_931 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n678_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_));
INVX1 INVX1_932 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n687_));
INVX1 INVX1_933 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n693_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n694_));
INVX1 INVX1_934 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n697_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n698_));
INVX1 INVX1_935 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n701_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n702_));
INVX1 INVX1_936 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n705_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_));
INVX1 INVX1_937 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n712_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n717_));
INVX1 INVX1_938 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n715_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n718_));
INVX1 INVX1_939 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n721_));
INVX1 INVX1_94 ( .A(\key_out[12] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3060_));
INVX1 INVX1_940 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n727_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n729_));
INVX1 INVX1_941 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n735_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n736_));
INVX1 INVX1_942 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n740_));
INVX1 INVX1_943 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n746_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n747_));
INVX1 INVX1_944 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n749_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n750_));
INVX1 INVX1_945 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n753_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n754_));
INVX1 INVX1_946 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n757_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_));
INVX1 INVX1_947 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n765_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n766_));
INVX1 INVX1_948 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n768_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n770_));
INVX1 INVX1_949 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n772_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_));
INVX1 INVX1_95 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3066_));
INVX1 INVX1_950 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n779_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n780_));
INVX1 INVX1_951 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n783_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n784_));
INVX1 INVX1_952 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n788_));
INVX1 INVX1_953 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n797_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n798_));
INVX1 INVX1_954 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n799_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n800_));
INVX1 INVX1_955 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n802_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_));
INVX1 INVX1_956 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n809_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n810_));
INVX1 INVX1_957 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n814_));
INVX1 INVX1_958 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n821_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n822_));
INVX1 INVX1_959 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n824_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n825_));
INVX1 INVX1_96 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3068_));
INVX1 INVX1_960 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n829_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n830_));
INVX1 INVX1_961 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n832_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_));
INVX1 INVX1_962 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n841_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n842_));
INVX1 INVX1_963 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n843_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n844_));
INVX1 INVX1_964 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n847_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_26_));
INVX1 INVX1_965 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n855_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n856_));
INVX1 INVX1_966 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n858_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n859_));
INVX1 INVX1_967 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n862_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n863_));
INVX1 INVX1_968 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n868_));
INVX1 INVX1_969 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n873_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n874_));
INVX1 INVX1_97 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3070_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3071_));
INVX1 INVX1_970 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n878_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n879_));
INVX1 INVX1_971 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n881_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n882_));
INVX1 INVX1_972 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n885_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_));
INVX1 INVX1_973 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n892_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n893_));
INVX1 INVX1_974 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n896_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n898_));
INVX1 INVX1_975 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n900_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_));
INVX1 INVX1_976 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n907_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n909_));
INVX1 INVX1_977 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n911_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n912_));
INVX1 INVX1_978 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n916_));
INVX1 INVX1_979 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n922_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n923_));
INVX1 INVX1_98 ( .A(\key_out[13] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n3078_));
INVX1 INVX1_980 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n926_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_31_));
INVX1 INVX1_981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n50_));
INVX1 INVX1_982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n52_));
INVX1 INVX1_983 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n55_));
INVX1 INVX1_984 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n57_));
INVX1 INVX1_985 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n59_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n60_));
INVX1 INVX1_986 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n54_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n62_));
INVX1 INVX1_987 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_));
INVX1 INVX1_988 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n67_));
INVX1 INVX1_989 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n72_));
INVX1 INVX1_99 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3084_));
INVX1 INVX1_990 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n70_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n73_));
INVX1 INVX1_991 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_));
INVX1 INVX1_992 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n81_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n82_));
INVX1 INVX1_993 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_));
INVX1 INVX1_994 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n93_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n94_));
INVX1 INVX1_995 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n98_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n99_));
INVX1 INVX1_996 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n100_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_));
INVX1 INVX1_997 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n102_));
INVX1 INVX1_998 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n105_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n107_));
INVX1 INVX1_999 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n113_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n114_));
OR2X2 OR2X2_1 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n73_), .B(\aes_mode[0] ), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n74_));
OR2X2 OR2X2_10 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n122_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n123_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_0_));
OR2X2 OR2X2_100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2524_), .B(AES_CORE_DATAPATH__abc_16009_new_n2522_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2525_));
OR2X2 OR2X2_1000 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4827_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4828_));
OR2X2 OR2X2_1001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4829_));
OR2X2 OR2X2_1002 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4831_));
OR2X2 OR2X2_1003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4832_), .B(AES_CORE_DATAPATH__abc_16009_new_n4833_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4834_));
OR2X2 OR2X2_1004 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4834_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4835_));
OR2X2 OR2X2_1005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4837_), .B(AES_CORE_DATAPATH__abc_16009_new_n4838_), .Y(AES_CORE_DATAPATH__0key_1__31_0__29_));
OR2X2 OR2X2_1006 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4840_));
OR2X2 OR2X2_1007 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4841_), .B(AES_CORE_DATAPATH__abc_16009_new_n4842_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4843_));
OR2X2 OR2X2_1008 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4843_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4844_));
OR2X2 OR2X2_1009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4845_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4846_));
OR2X2 OR2X2_101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2526_));
OR2X2 OR2X2_1010 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4847_));
OR2X2 OR2X2_1011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4849_), .B(AES_CORE_DATAPATH__abc_16009_new_n4850_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4851_));
OR2X2 OR2X2_1012 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4851_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4852_));
OR2X2 OR2X2_1013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4853_));
OR2X2 OR2X2_1014 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4855_), .B(AES_CORE_DATAPATH__abc_16009_new_n4856_), .Y(AES_CORE_DATAPATH__0key_1__31_0__31_));
OR2X2 OR2X2_1015 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4858_), .B(AES_CORE_DATAPATH__abc_16009_new_n4859_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4860_));
OR2X2 OR2X2_1016 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4868_), .B(AES_CORE_DATAPATH__abc_16009_new_n4867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4869_));
OR2X2 OR2X2_1017 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4870_), .B(AES_CORE_DATAPATH__abc_16009_new_n4866_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4871_));
OR2X2 OR2X2_1018 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4872_), .B(AES_CORE_DATAPATH__abc_16009_new_n4873_), .Y(AES_CORE_DATAPATH__0key_0__31_0__0_));
OR2X2 OR2X2_1019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_97_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4875_));
OR2X2 OR2X2_102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2528_), .B(AES_CORE_DATAPATH__abc_16009_new_n2529_), .Y(\iv_out[4] ));
OR2X2 OR2X2_1020 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4876_), .B(AES_CORE_DATAPATH__abc_16009_new_n4877_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4878_));
OR2X2 OR2X2_1021 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4878_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4879_));
OR2X2 OR2X2_1022 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4881_), .B(AES_CORE_DATAPATH__abc_16009_new_n4882_), .Y(AES_CORE_DATAPATH__0key_0__31_0__1_));
OR2X2 OR2X2_1023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_98_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4884_));
OR2X2 OR2X2_1024 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4885_), .B(AES_CORE_DATAPATH__abc_16009_new_n4886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4887_));
OR2X2 OR2X2_1025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4887_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4888_));
OR2X2 OR2X2_1026 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4890_), .B(AES_CORE_DATAPATH__abc_16009_new_n4891_), .Y(AES_CORE_DATAPATH__0key_0__31_0__2_));
OR2X2 OR2X2_1027 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_99_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4893_));
OR2X2 OR2X2_1028 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4894_), .B(AES_CORE_DATAPATH__abc_16009_new_n4895_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4896_));
OR2X2 OR2X2_1029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4896_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4897_));
OR2X2 OR2X2_103 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2533_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2534_));
OR2X2 OR2X2_1030 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4899_), .B(AES_CORE_DATAPATH__abc_16009_new_n4900_), .Y(AES_CORE_DATAPATH__0key_0__31_0__3_));
OR2X2 OR2X2_1031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4902_));
OR2X2 OR2X2_1032 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4903_), .B(AES_CORE_DATAPATH__abc_16009_new_n4904_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4905_));
OR2X2 OR2X2_1033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4905_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4906_));
OR2X2 OR2X2_1034 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4907_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4908_));
OR2X2 OR2X2_1035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4909_));
OR2X2 OR2X2_1036 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_101_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4911_));
OR2X2 OR2X2_1037 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4912_), .B(AES_CORE_DATAPATH__abc_16009_new_n4913_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4914_));
OR2X2 OR2X2_1038 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4914_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4915_));
OR2X2 OR2X2_1039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4917_), .B(AES_CORE_DATAPATH__abc_16009_new_n4918_), .Y(AES_CORE_DATAPATH__0key_0__31_0__5_));
OR2X2 OR2X2_104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2534_), .B(AES_CORE_DATAPATH__abc_16009_new_n2532_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2535_));
OR2X2 OR2X2_1040 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4920_));
OR2X2 OR2X2_1041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4921_), .B(AES_CORE_DATAPATH__abc_16009_new_n4922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4923_));
OR2X2 OR2X2_1042 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4923_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4924_));
OR2X2 OR2X2_1043 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4925_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4926_));
OR2X2 OR2X2_1044 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4927_));
OR2X2 OR2X2_1045 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4929_));
OR2X2 OR2X2_1046 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4930_), .B(AES_CORE_DATAPATH__abc_16009_new_n4931_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4932_));
OR2X2 OR2X2_1047 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4932_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4933_));
OR2X2 OR2X2_1048 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4935_), .B(AES_CORE_DATAPATH__abc_16009_new_n4936_), .Y(AES_CORE_DATAPATH__0key_0__31_0__7_));
OR2X2 OR2X2_1049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_104_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4938_));
OR2X2 OR2X2_105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2536_));
OR2X2 OR2X2_1050 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4939_), .B(AES_CORE_DATAPATH__abc_16009_new_n4940_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4941_));
OR2X2 OR2X2_1051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4941_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4942_));
OR2X2 OR2X2_1052 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4944_), .B(AES_CORE_DATAPATH__abc_16009_new_n4945_), .Y(AES_CORE_DATAPATH__0key_0__31_0__8_));
OR2X2 OR2X2_1053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_105_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4947_));
OR2X2 OR2X2_1054 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4948_), .B(AES_CORE_DATAPATH__abc_16009_new_n4949_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4950_));
OR2X2 OR2X2_1055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4950_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4951_));
OR2X2 OR2X2_1056 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4952_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4953_));
OR2X2 OR2X2_1057 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4954_));
OR2X2 OR2X2_1058 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_106_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4956_));
OR2X2 OR2X2_1059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4957_), .B(AES_CORE_DATAPATH__abc_16009_new_n4958_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4959_));
OR2X2 OR2X2_106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2538_), .B(AES_CORE_DATAPATH__abc_16009_new_n2539_), .Y(\iv_out[5] ));
OR2X2 OR2X2_1060 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4959_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4960_));
OR2X2 OR2X2_1061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4962_), .B(AES_CORE_DATAPATH__abc_16009_new_n4963_), .Y(AES_CORE_DATAPATH__0key_0__31_0__10_));
OR2X2 OR2X2_1062 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_107_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4965_));
OR2X2 OR2X2_1063 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4966_), .B(AES_CORE_DATAPATH__abc_16009_new_n4967_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4968_));
OR2X2 OR2X2_1064 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4968_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4969_));
OR2X2 OR2X2_1065 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4971_), .B(AES_CORE_DATAPATH__abc_16009_new_n4972_), .Y(AES_CORE_DATAPATH__0key_0__31_0__11_));
OR2X2 OR2X2_1066 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_108_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4974_));
OR2X2 OR2X2_1067 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4975_), .B(AES_CORE_DATAPATH__abc_16009_new_n4976_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4977_));
OR2X2 OR2X2_1068 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4977_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4978_));
OR2X2 OR2X2_1069 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4980_), .B(AES_CORE_DATAPATH__abc_16009_new_n4981_), .Y(AES_CORE_DATAPATH__0key_0__31_0__12_));
OR2X2 OR2X2_107 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2543_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2544_));
OR2X2 OR2X2_1070 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4983_));
OR2X2 OR2X2_1071 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4984_), .B(AES_CORE_DATAPATH__abc_16009_new_n4985_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4986_));
OR2X2 OR2X2_1072 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4986_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4987_));
OR2X2 OR2X2_1073 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4988_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4989_));
OR2X2 OR2X2_1074 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4990_));
OR2X2 OR2X2_1075 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4992_));
OR2X2 OR2X2_1076 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4993_), .B(AES_CORE_DATAPATH__abc_16009_new_n4994_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4995_));
OR2X2 OR2X2_1077 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4995_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4996_));
OR2X2 OR2X2_1078 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4998_), .B(AES_CORE_DATAPATH__abc_16009_new_n4999_), .Y(AES_CORE_DATAPATH__0key_0__31_0__14_));
OR2X2 OR2X2_1079 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_111_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5001_));
OR2X2 OR2X2_108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2544_), .B(AES_CORE_DATAPATH__abc_16009_new_n2542_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2545_));
OR2X2 OR2X2_1080 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5002_), .B(AES_CORE_DATAPATH__abc_16009_new_n5003_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5004_));
OR2X2 OR2X2_1081 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5004_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5005_));
OR2X2 OR2X2_1082 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5007_), .B(AES_CORE_DATAPATH__abc_16009_new_n5008_), .Y(AES_CORE_DATAPATH__0key_0__31_0__15_));
OR2X2 OR2X2_1083 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_112_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5010_));
OR2X2 OR2X2_1084 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5011_), .B(AES_CORE_DATAPATH__abc_16009_new_n5012_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5013_));
OR2X2 OR2X2_1085 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5013_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5014_));
OR2X2 OR2X2_1086 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5016_), .B(AES_CORE_DATAPATH__abc_16009_new_n5017_), .Y(AES_CORE_DATAPATH__0key_0__31_0__16_));
OR2X2 OR2X2_1087 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5019_));
OR2X2 OR2X2_1088 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5020_), .B(AES_CORE_DATAPATH__abc_16009_new_n5021_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5022_));
OR2X2 OR2X2_1089 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5022_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5023_));
OR2X2 OR2X2_109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2546_));
OR2X2 OR2X2_1090 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5025_), .B(AES_CORE_DATAPATH__abc_16009_new_n5026_), .Y(AES_CORE_DATAPATH__0key_0__31_0__17_));
OR2X2 OR2X2_1091 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_114_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5028_));
OR2X2 OR2X2_1092 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5029_), .B(AES_CORE_DATAPATH__abc_16009_new_n5030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5031_));
OR2X2 OR2X2_1093 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5032_));
OR2X2 OR2X2_1094 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5034_), .B(AES_CORE_DATAPATH__abc_16009_new_n5035_), .Y(AES_CORE_DATAPATH__0key_0__31_0__18_));
OR2X2 OR2X2_1095 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_115_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5037_));
OR2X2 OR2X2_1096 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5038_), .B(AES_CORE_DATAPATH__abc_16009_new_n5039_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5040_));
OR2X2 OR2X2_1097 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5040_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5041_));
OR2X2 OR2X2_1098 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5043_), .B(AES_CORE_DATAPATH__abc_16009_new_n5044_), .Y(AES_CORE_DATAPATH__0key_0__31_0__19_));
OR2X2 OR2X2_1099 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_116_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5046_));
OR2X2 OR2X2_11 ( .A(AES_CORE_CONTROL_UNIT_rd_count_1_), .B(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n126_));
OR2X2 OR2X2_110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2548_), .B(AES_CORE_DATAPATH__abc_16009_new_n2549_), .Y(\iv_out[6] ));
OR2X2 OR2X2_1100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5047_), .B(AES_CORE_DATAPATH__abc_16009_new_n5048_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5049_));
OR2X2 OR2X2_1101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5049_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5050_));
OR2X2 OR2X2_1102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5051_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5052_));
OR2X2 OR2X2_1103 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5053_));
OR2X2 OR2X2_1104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5055_));
OR2X2 OR2X2_1105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5056_), .B(AES_CORE_DATAPATH__abc_16009_new_n5057_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5058_));
OR2X2 OR2X2_1106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5058_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5059_));
OR2X2 OR2X2_1107 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5061_), .B(AES_CORE_DATAPATH__abc_16009_new_n5062_), .Y(AES_CORE_DATAPATH__0key_0__31_0__21_));
OR2X2 OR2X2_1108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_118_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5064_));
OR2X2 OR2X2_1109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5065_), .B(AES_CORE_DATAPATH__abc_16009_new_n5066_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5067_));
OR2X2 OR2X2_111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2553_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2554_));
OR2X2 OR2X2_1110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5067_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5068_));
OR2X2 OR2X2_1111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5070_), .B(AES_CORE_DATAPATH__abc_16009_new_n5071_), .Y(AES_CORE_DATAPATH__0key_0__31_0__22_));
OR2X2 OR2X2_1112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_119_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5073_));
OR2X2 OR2X2_1113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5074_), .B(AES_CORE_DATAPATH__abc_16009_new_n5075_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5076_));
OR2X2 OR2X2_1114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5076_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5077_));
OR2X2 OR2X2_1115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5078_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5079_));
OR2X2 OR2X2_1116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5080_));
OR2X2 OR2X2_1117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5082_));
OR2X2 OR2X2_1118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5083_), .B(AES_CORE_DATAPATH__abc_16009_new_n5084_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5085_));
OR2X2 OR2X2_1119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5085_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5086_));
OR2X2 OR2X2_112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2554_), .B(AES_CORE_DATAPATH__abc_16009_new_n2552_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2555_));
OR2X2 OR2X2_1120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5087_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5088_));
OR2X2 OR2X2_1121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5089_));
OR2X2 OR2X2_1122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_121_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5091_));
OR2X2 OR2X2_1123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5092_), .B(AES_CORE_DATAPATH__abc_16009_new_n5093_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5094_));
OR2X2 OR2X2_1124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5094_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5095_));
OR2X2 OR2X2_1125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5097_), .B(AES_CORE_DATAPATH__abc_16009_new_n5098_), .Y(AES_CORE_DATAPATH__0key_0__31_0__25_));
OR2X2 OR2X2_1126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5100_));
OR2X2 OR2X2_1127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5101_), .B(AES_CORE_DATAPATH__abc_16009_new_n5102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5103_));
OR2X2 OR2X2_1128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5104_));
OR2X2 OR2X2_1129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5105_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5106_));
OR2X2 OR2X2_113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2556_));
OR2X2 OR2X2_1130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5107_));
OR2X2 OR2X2_1131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_123_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5109_));
OR2X2 OR2X2_1132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5110_), .B(AES_CORE_DATAPATH__abc_16009_new_n5111_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5112_));
OR2X2 OR2X2_1133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5112_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5113_));
OR2X2 OR2X2_1134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5115_), .B(AES_CORE_DATAPATH__abc_16009_new_n5116_), .Y(AES_CORE_DATAPATH__0key_0__31_0__27_));
OR2X2 OR2X2_1135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5118_));
OR2X2 OR2X2_1136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5119_), .B(AES_CORE_DATAPATH__abc_16009_new_n5120_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5121_));
OR2X2 OR2X2_1137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5121_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5122_));
OR2X2 OR2X2_1138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5123_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5124_));
OR2X2 OR2X2_1139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5125_));
OR2X2 OR2X2_114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2558_), .B(AES_CORE_DATAPATH__abc_16009_new_n2559_), .Y(\iv_out[7] ));
OR2X2 OR2X2_1140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5127_));
OR2X2 OR2X2_1141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5128_), .B(AES_CORE_DATAPATH__abc_16009_new_n5129_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5130_));
OR2X2 OR2X2_1142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5130_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5131_));
OR2X2 OR2X2_1143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5133_), .B(AES_CORE_DATAPATH__abc_16009_new_n5134_), .Y(AES_CORE_DATAPATH__0key_0__31_0__29_));
OR2X2 OR2X2_1144 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5136_));
OR2X2 OR2X2_1145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5137_), .B(AES_CORE_DATAPATH__abc_16009_new_n5138_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5139_));
OR2X2 OR2X2_1146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5139_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5140_));
OR2X2 OR2X2_1147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5141_), .B(AES_CORE_DATAPATH__abc_16009_new_n4864_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5142_));
OR2X2 OR2X2_1148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4865_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5143_));
OR2X2 OR2X2_1149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5145_), .B(AES_CORE_DATAPATH__abc_16009_new_n5146_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5147_));
OR2X2 OR2X2_115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2563_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2564_));
OR2X2 OR2X2_1150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5147_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5148_));
OR2X2 OR2X2_1151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5149_));
OR2X2 OR2X2_1152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5151_), .B(AES_CORE_DATAPATH__abc_16009_new_n5152_), .Y(AES_CORE_DATAPATH__0key_0__31_0__31_));
OR2X2 OR2X2_1153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5156_), .B(AES_CORE_DATAPATH__abc_16009_new_n5154_), .Y(AES_CORE_DATAPATH__0key_host_0__31_0__0_));
OR2X2 OR2X2_1154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5158_));
OR2X2 OR2X2_1155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4878_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5159_));
OR2X2 OR2X2_1156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5161_));
OR2X2 OR2X2_1157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4887_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5162_));
OR2X2 OR2X2_1158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5164_));
OR2X2 OR2X2_1159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4896_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5165_));
OR2X2 OR2X2_116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2564_), .B(AES_CORE_DATAPATH__abc_16009_new_n2562_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2565_));
OR2X2 OR2X2_1160 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5167_));
OR2X2 OR2X2_1161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4905_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5168_));
OR2X2 OR2X2_1162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5170_));
OR2X2 OR2X2_1163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4914_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5171_));
OR2X2 OR2X2_1164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5173_));
OR2X2 OR2X2_1165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4923_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5174_));
OR2X2 OR2X2_1166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5176_));
OR2X2 OR2X2_1167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4932_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5177_));
OR2X2 OR2X2_1168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5179_));
OR2X2 OR2X2_1169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4941_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5180_));
OR2X2 OR2X2_117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2566_));
OR2X2 OR2X2_1170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5182_));
OR2X2 OR2X2_1171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4950_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5183_));
OR2X2 OR2X2_1172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5185_));
OR2X2 OR2X2_1173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4959_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5186_));
OR2X2 OR2X2_1174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5188_));
OR2X2 OR2X2_1175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4968_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5189_));
OR2X2 OR2X2_1176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5191_));
OR2X2 OR2X2_1177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4977_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5192_));
OR2X2 OR2X2_1178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5194_));
OR2X2 OR2X2_1179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4986_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5195_));
OR2X2 OR2X2_118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2568_), .B(AES_CORE_DATAPATH__abc_16009_new_n2569_), .Y(\iv_out[8] ));
OR2X2 OR2X2_1180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5197_));
OR2X2 OR2X2_1181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4995_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5198_));
OR2X2 OR2X2_1182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5200_));
OR2X2 OR2X2_1183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5004_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5201_));
OR2X2 OR2X2_1184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5203_));
OR2X2 OR2X2_1185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5013_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5204_));
OR2X2 OR2X2_1186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5206_));
OR2X2 OR2X2_1187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5022_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5207_));
OR2X2 OR2X2_1188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5209_));
OR2X2 OR2X2_1189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5031_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5210_));
OR2X2 OR2X2_119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2573_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2574_));
OR2X2 OR2X2_1190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5212_));
OR2X2 OR2X2_1191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5040_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5213_));
OR2X2 OR2X2_1192 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5215_));
OR2X2 OR2X2_1193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5049_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5216_));
OR2X2 OR2X2_1194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5218_));
OR2X2 OR2X2_1195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5058_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5219_));
OR2X2 OR2X2_1196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5221_));
OR2X2 OR2X2_1197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5067_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5222_));
OR2X2 OR2X2_1198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5224_));
OR2X2 OR2X2_1199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5076_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5225_));
OR2X2 OR2X2_12 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n131_), .B(AES_CORE_CONTROL_UNIT_state_15_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n132_));
OR2X2 OR2X2_120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2574_), .B(AES_CORE_DATAPATH__abc_16009_new_n2572_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2575_));
OR2X2 OR2X2_1200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5227_));
OR2X2 OR2X2_1201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5085_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5228_));
OR2X2 OR2X2_1202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5230_));
OR2X2 OR2X2_1203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5094_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5231_));
OR2X2 OR2X2_1204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5233_));
OR2X2 OR2X2_1205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5103_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5234_));
OR2X2 OR2X2_1206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5236_));
OR2X2 OR2X2_1207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5112_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5237_));
OR2X2 OR2X2_1208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5239_));
OR2X2 OR2X2_1209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5121_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5240_));
OR2X2 OR2X2_121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2576_));
OR2X2 OR2X2_1210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5242_));
OR2X2 OR2X2_1211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5130_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5243_));
OR2X2 OR2X2_1212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5245_));
OR2X2 OR2X2_1213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5139_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5246_));
OR2X2 OR2X2_1214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5147_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5248_));
OR2X2 OR2X2_1215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5249_));
OR2X2 OR2X2_1216 ( .A(\key_en[2] ), .B(AES_CORE_DATAPATH_key_host_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5252_));
OR2X2 OR2X2_1217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5253_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n5254_));
OR2X2 OR2X2_1218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5256_), .B(AES_CORE_DATAPATH__abc_16009_new_n5251_), .Y(AES_CORE_DATAPATH__0key_host_2__31_0__0_));
OR2X2 OR2X2_1219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5258_));
OR2X2 OR2X2_122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2578_), .B(AES_CORE_DATAPATH__abc_16009_new_n2579_), .Y(\iv_out[9] ));
OR2X2 OR2X2_1220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5259_), .B(AES_CORE_DATAPATH__abc_16009_new_n5260_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5261_));
OR2X2 OR2X2_1221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5261_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5262_));
OR2X2 OR2X2_1222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5264_));
OR2X2 OR2X2_1223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5265_), .B(AES_CORE_DATAPATH__abc_16009_new_n5266_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5267_));
OR2X2 OR2X2_1224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5267_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5268_));
OR2X2 OR2X2_1225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5270_));
OR2X2 OR2X2_1226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5271_), .B(AES_CORE_DATAPATH__abc_16009_new_n5272_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5273_));
OR2X2 OR2X2_1227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5273_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5274_));
OR2X2 OR2X2_1228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5276_));
OR2X2 OR2X2_1229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5277_), .B(AES_CORE_DATAPATH__abc_16009_new_n5278_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5279_));
OR2X2 OR2X2_123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2583_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2584_));
OR2X2 OR2X2_1230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5279_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5280_));
OR2X2 OR2X2_1231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5282_));
OR2X2 OR2X2_1232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5283_), .B(AES_CORE_DATAPATH__abc_16009_new_n5284_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5285_));
OR2X2 OR2X2_1233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5285_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5286_));
OR2X2 OR2X2_1234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5288_));
OR2X2 OR2X2_1235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5289_), .B(AES_CORE_DATAPATH__abc_16009_new_n5290_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5291_));
OR2X2 OR2X2_1236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5291_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5292_));
OR2X2 OR2X2_1237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5294_));
OR2X2 OR2X2_1238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5295_), .B(AES_CORE_DATAPATH__abc_16009_new_n5296_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5297_));
OR2X2 OR2X2_1239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5297_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5298_));
OR2X2 OR2X2_124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2584_), .B(AES_CORE_DATAPATH__abc_16009_new_n2582_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2585_));
OR2X2 OR2X2_1240 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5300_));
OR2X2 OR2X2_1241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5301_), .B(AES_CORE_DATAPATH__abc_16009_new_n5302_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5303_));
OR2X2 OR2X2_1242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5303_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5304_));
OR2X2 OR2X2_1243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5306_));
OR2X2 OR2X2_1244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5307_), .B(AES_CORE_DATAPATH__abc_16009_new_n5308_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5309_));
OR2X2 OR2X2_1245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5309_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5310_));
OR2X2 OR2X2_1246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5312_));
OR2X2 OR2X2_1247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5313_), .B(AES_CORE_DATAPATH__abc_16009_new_n5314_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5315_));
OR2X2 OR2X2_1248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5315_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5316_));
OR2X2 OR2X2_1249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5318_));
OR2X2 OR2X2_125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2586_));
OR2X2 OR2X2_1250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5319_), .B(AES_CORE_DATAPATH__abc_16009_new_n5320_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5321_));
OR2X2 OR2X2_1251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5321_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5322_));
OR2X2 OR2X2_1252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5324_));
OR2X2 OR2X2_1253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5325_), .B(AES_CORE_DATAPATH__abc_16009_new_n5326_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5327_));
OR2X2 OR2X2_1254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5327_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5328_));
OR2X2 OR2X2_1255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5330_));
OR2X2 OR2X2_1256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5331_), .B(AES_CORE_DATAPATH__abc_16009_new_n5332_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5333_));
OR2X2 OR2X2_1257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5333_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5334_));
OR2X2 OR2X2_1258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5336_));
OR2X2 OR2X2_1259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5337_), .B(AES_CORE_DATAPATH__abc_16009_new_n5338_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5339_));
OR2X2 OR2X2_126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2588_), .B(AES_CORE_DATAPATH__abc_16009_new_n2589_), .Y(\iv_out[10] ));
OR2X2 OR2X2_1260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5339_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5340_));
OR2X2 OR2X2_1261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5342_));
OR2X2 OR2X2_1262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5343_), .B(AES_CORE_DATAPATH__abc_16009_new_n5344_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5345_));
OR2X2 OR2X2_1263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5345_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5346_));
OR2X2 OR2X2_1264 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5348_));
OR2X2 OR2X2_1265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5349_), .B(AES_CORE_DATAPATH__abc_16009_new_n5350_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5351_));
OR2X2 OR2X2_1266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5351_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5352_));
OR2X2 OR2X2_1267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5354_));
OR2X2 OR2X2_1268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5355_), .B(AES_CORE_DATAPATH__abc_16009_new_n5356_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5357_));
OR2X2 OR2X2_1269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5357_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5358_));
OR2X2 OR2X2_127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2593_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2594_));
OR2X2 OR2X2_1270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5360_));
OR2X2 OR2X2_1271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5361_), .B(AES_CORE_DATAPATH__abc_16009_new_n5362_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5363_));
OR2X2 OR2X2_1272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5363_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5364_));
OR2X2 OR2X2_1273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5366_));
OR2X2 OR2X2_1274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5367_), .B(AES_CORE_DATAPATH__abc_16009_new_n5368_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5369_));
OR2X2 OR2X2_1275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5369_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5370_));
OR2X2 OR2X2_1276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5372_));
OR2X2 OR2X2_1277 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5373_), .B(AES_CORE_DATAPATH__abc_16009_new_n5374_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5375_));
OR2X2 OR2X2_1278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5375_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5376_));
OR2X2 OR2X2_1279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5378_));
OR2X2 OR2X2_128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2594_), .B(AES_CORE_DATAPATH__abc_16009_new_n2592_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2595_));
OR2X2 OR2X2_1280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5379_), .B(AES_CORE_DATAPATH__abc_16009_new_n5380_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5381_));
OR2X2 OR2X2_1281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5381_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5382_));
OR2X2 OR2X2_1282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5384_));
OR2X2 OR2X2_1283 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5385_), .B(AES_CORE_DATAPATH__abc_16009_new_n5386_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5387_));
OR2X2 OR2X2_1284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5387_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5388_));
OR2X2 OR2X2_1285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5390_));
OR2X2 OR2X2_1286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5391_), .B(AES_CORE_DATAPATH__abc_16009_new_n5392_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5393_));
OR2X2 OR2X2_1287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5393_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5394_));
OR2X2 OR2X2_1288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5396_));
OR2X2 OR2X2_1289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5397_), .B(AES_CORE_DATAPATH__abc_16009_new_n5398_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5399_));
OR2X2 OR2X2_129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2596_));
OR2X2 OR2X2_1290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5399_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5400_));
OR2X2 OR2X2_1291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5402_));
OR2X2 OR2X2_1292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5403_), .B(AES_CORE_DATAPATH__abc_16009_new_n5404_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5405_));
OR2X2 OR2X2_1293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5405_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5406_));
OR2X2 OR2X2_1294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5408_));
OR2X2 OR2X2_1295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5409_), .B(AES_CORE_DATAPATH__abc_16009_new_n5410_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5411_));
OR2X2 OR2X2_1296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5411_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5412_));
OR2X2 OR2X2_1297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5414_));
OR2X2 OR2X2_1298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5415_), .B(AES_CORE_DATAPATH__abc_16009_new_n5416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5417_));
OR2X2 OR2X2_1299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5417_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5418_));
OR2X2 OR2X2_13 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n133_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n125_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_6_));
OR2X2 OR2X2_130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2598_), .B(AES_CORE_DATAPATH__abc_16009_new_n2599_), .Y(\iv_out[11] ));
OR2X2 OR2X2_1300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5420_));
OR2X2 OR2X2_1301 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5421_), .B(AES_CORE_DATAPATH__abc_16009_new_n5422_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5423_));
OR2X2 OR2X2_1302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5423_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5424_));
OR2X2 OR2X2_1303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5426_));
OR2X2 OR2X2_1304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5427_), .B(AES_CORE_DATAPATH__abc_16009_new_n5428_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5429_));
OR2X2 OR2X2_1305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5429_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5430_));
OR2X2 OR2X2_1306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5432_));
OR2X2 OR2X2_1307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5433_), .B(AES_CORE_DATAPATH__abc_16009_new_n5434_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5435_));
OR2X2 OR2X2_1308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5435_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5436_));
OR2X2 OR2X2_1309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5438_), .B(AES_CORE_DATAPATH__abc_16009_new_n5439_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5440_));
OR2X2 OR2X2_131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2603_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2604_));
OR2X2 OR2X2_1310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5440_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5441_));
OR2X2 OR2X2_1311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5442_));
OR2X2 OR2X2_1312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5445_), .B(AES_CORE_DATAPATH__abc_16009_new_n5444_), .Y(AES_CORE_DATAPATH__0key_host_1__31_0__0_));
OR2X2 OR2X2_1313 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4582_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5447_));
OR2X2 OR2X2_1314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5448_));
OR2X2 OR2X2_1315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4591_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5450_));
OR2X2 OR2X2_1316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5451_));
OR2X2 OR2X2_1317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4600_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5453_));
OR2X2 OR2X2_1318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5454_));
OR2X2 OR2X2_1319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4609_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5456_));
OR2X2 OR2X2_132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2604_), .B(AES_CORE_DATAPATH__abc_16009_new_n2602_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2605_));
OR2X2 OR2X2_1320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5457_));
OR2X2 OR2X2_1321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4618_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5459_));
OR2X2 OR2X2_1322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5460_));
OR2X2 OR2X2_1323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4627_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5462_));
OR2X2 OR2X2_1324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5463_));
OR2X2 OR2X2_1325 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4636_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5465_));
OR2X2 OR2X2_1326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5466_));
OR2X2 OR2X2_1327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4645_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5468_));
OR2X2 OR2X2_1328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5469_));
OR2X2 OR2X2_1329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4654_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5471_));
OR2X2 OR2X2_133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2606_));
OR2X2 OR2X2_1330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5472_));
OR2X2 OR2X2_1331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4663_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5474_));
OR2X2 OR2X2_1332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5475_));
OR2X2 OR2X2_1333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4672_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5477_));
OR2X2 OR2X2_1334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5478_));
OR2X2 OR2X2_1335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4681_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5480_));
OR2X2 OR2X2_1336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5481_));
OR2X2 OR2X2_1337 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4690_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5483_));
OR2X2 OR2X2_1338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5484_));
OR2X2 OR2X2_1339 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4699_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5486_));
OR2X2 OR2X2_134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2608_), .B(AES_CORE_DATAPATH__abc_16009_new_n2609_), .Y(\iv_out[12] ));
OR2X2 OR2X2_1340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5487_));
OR2X2 OR2X2_1341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4708_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5489_));
OR2X2 OR2X2_1342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5490_));
OR2X2 OR2X2_1343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4717_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5492_));
OR2X2 OR2X2_1344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5493_));
OR2X2 OR2X2_1345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4726_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5495_));
OR2X2 OR2X2_1346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5496_));
OR2X2 OR2X2_1347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4735_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5498_));
OR2X2 OR2X2_1348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5499_));
OR2X2 OR2X2_1349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4744_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5501_));
OR2X2 OR2X2_135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2613_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2614_));
OR2X2 OR2X2_1350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5502_));
OR2X2 OR2X2_1351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4753_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5504_));
OR2X2 OR2X2_1352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5505_));
OR2X2 OR2X2_1353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4762_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5507_));
OR2X2 OR2X2_1354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5508_));
OR2X2 OR2X2_1355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4771_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5510_));
OR2X2 OR2X2_1356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5511_));
OR2X2 OR2X2_1357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4780_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5513_));
OR2X2 OR2X2_1358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5514_));
OR2X2 OR2X2_1359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4789_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5516_));
OR2X2 OR2X2_136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2614_), .B(AES_CORE_DATAPATH__abc_16009_new_n2612_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2615_));
OR2X2 OR2X2_1360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5517_));
OR2X2 OR2X2_1361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4798_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5519_));
OR2X2 OR2X2_1362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5520_));
OR2X2 OR2X2_1363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4807_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5522_));
OR2X2 OR2X2_1364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5523_));
OR2X2 OR2X2_1365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4816_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5525_));
OR2X2 OR2X2_1366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5526_));
OR2X2 OR2X2_1367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4825_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5528_));
OR2X2 OR2X2_1368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5529_));
OR2X2 OR2X2_1369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4834_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5531_));
OR2X2 OR2X2_137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2616_));
OR2X2 OR2X2_1370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5532_));
OR2X2 OR2X2_1371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4843_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5534_));
OR2X2 OR2X2_1372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5535_));
OR2X2 OR2X2_1373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5537_));
OR2X2 OR2X2_1374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4851_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n5538_));
OR2X2 OR2X2_1375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5540_), .B(AES_CORE_DATAPATH__abc_16009_new_n5541_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5542_));
OR2X2 OR2X2_1376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5255_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5546_));
OR2X2 OR2X2_1377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_32_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5547_));
OR2X2 OR2X2_1378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5548_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5549_));
OR2X2 OR2X2_1379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5551_));
OR2X2 OR2X2_138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2618_), .B(AES_CORE_DATAPATH__abc_16009_new_n2619_), .Y(\iv_out[13] ));
OR2X2 OR2X2_1380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5261_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5553_));
OR2X2 OR2X2_1381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_33_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5554_));
OR2X2 OR2X2_1382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5555_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5556_));
OR2X2 OR2X2_1383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5557_));
OR2X2 OR2X2_1384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5267_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5559_));
OR2X2 OR2X2_1385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_34_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5560_));
OR2X2 OR2X2_1386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5561_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5562_));
OR2X2 OR2X2_1387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5563_));
OR2X2 OR2X2_1388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_35_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5565_));
OR2X2 OR2X2_1389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5273_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5566_));
OR2X2 OR2X2_139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2623_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2624_));
OR2X2 OR2X2_1390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5568_));
OR2X2 OR2X2_1391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5569_));
OR2X2 OR2X2_1392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_36_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5571_));
OR2X2 OR2X2_1393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5279_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5572_));
OR2X2 OR2X2_1394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5573_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5574_));
OR2X2 OR2X2_1395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5575_));
OR2X2 OR2X2_1396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5285_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5577_));
OR2X2 OR2X2_1397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_37_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5578_));
OR2X2 OR2X2_1398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5580_), .B(AES_CORE_DATAPATH__abc_16009_new_n5581_), .Y(AES_CORE_DATAPATH__0key_2__31_0__5_));
OR2X2 OR2X2_1399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_38_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5583_));
OR2X2 OR2X2_14 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n135_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n136_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_9_));
OR2X2 OR2X2_140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2624_), .B(AES_CORE_DATAPATH__abc_16009_new_n2622_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2625_));
OR2X2 OR2X2_1400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5291_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5584_));
OR2X2 OR2X2_1401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5585_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5586_));
OR2X2 OR2X2_1402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5587_));
OR2X2 OR2X2_1403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5297_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5589_));
OR2X2 OR2X2_1404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_39_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5590_));
OR2X2 OR2X2_1405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5591_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5592_));
OR2X2 OR2X2_1406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5593_));
OR2X2 OR2X2_1407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5303_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5595_));
OR2X2 OR2X2_1408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_40_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5596_));
OR2X2 OR2X2_1409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5597_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5598_));
OR2X2 OR2X2_141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2626_));
OR2X2 OR2X2_1410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5599_));
OR2X2 OR2X2_1411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5309_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5601_));
OR2X2 OR2X2_1412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_41_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5602_));
OR2X2 OR2X2_1413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5604_), .B(AES_CORE_DATAPATH__abc_16009_new_n5605_), .Y(AES_CORE_DATAPATH__0key_2__31_0__9_));
OR2X2 OR2X2_1414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5315_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5607_));
OR2X2 OR2X2_1415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_42_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5608_));
OR2X2 OR2X2_1416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5610_), .B(AES_CORE_DATAPATH__abc_16009_new_n5611_), .Y(AES_CORE_DATAPATH__0key_2__31_0__10_));
OR2X2 OR2X2_1417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5321_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5613_));
OR2X2 OR2X2_1418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_43_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5614_));
OR2X2 OR2X2_1419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5616_), .B(AES_CORE_DATAPATH__abc_16009_new_n5617_), .Y(AES_CORE_DATAPATH__0key_2__31_0__11_));
OR2X2 OR2X2_142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2628_), .B(AES_CORE_DATAPATH__abc_16009_new_n2629_), .Y(\iv_out[14] ));
OR2X2 OR2X2_1420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_44_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5619_));
OR2X2 OR2X2_1421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5327_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5620_));
OR2X2 OR2X2_1422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5621_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5622_));
OR2X2 OR2X2_1423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5623_));
OR2X2 OR2X2_1424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_45_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5625_));
OR2X2 OR2X2_1425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5333_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5626_));
OR2X2 OR2X2_1426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5627_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5628_));
OR2X2 OR2X2_1427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5629_));
OR2X2 OR2X2_1428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5339_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5631_));
OR2X2 OR2X2_1429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_46_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5632_));
OR2X2 OR2X2_143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2633_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2634_));
OR2X2 OR2X2_1430 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5634_), .B(AES_CORE_DATAPATH__abc_16009_new_n5635_), .Y(AES_CORE_DATAPATH__0key_2__31_0__14_));
OR2X2 OR2X2_1431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5345_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5637_));
OR2X2 OR2X2_1432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_47_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5638_));
OR2X2 OR2X2_1433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5640_), .B(AES_CORE_DATAPATH__abc_16009_new_n5641_), .Y(AES_CORE_DATAPATH__0key_2__31_0__15_));
OR2X2 OR2X2_1434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_48_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5643_));
OR2X2 OR2X2_1435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5351_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5644_));
OR2X2 OR2X2_1436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5645_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5646_));
OR2X2 OR2X2_1437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5647_));
OR2X2 OR2X2_1438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5357_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5649_));
OR2X2 OR2X2_1439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_49_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5650_));
OR2X2 OR2X2_144 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2634_), .B(AES_CORE_DATAPATH__abc_16009_new_n2632_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2635_));
OR2X2 OR2X2_1440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5652_), .B(AES_CORE_DATAPATH__abc_16009_new_n5653_), .Y(AES_CORE_DATAPATH__0key_2__31_0__17_));
OR2X2 OR2X2_1441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5363_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5655_));
OR2X2 OR2X2_1442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_50_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5656_));
OR2X2 OR2X2_1443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5658_), .B(AES_CORE_DATAPATH__abc_16009_new_n5659_), .Y(AES_CORE_DATAPATH__0key_2__31_0__18_));
OR2X2 OR2X2_1444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_51_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5661_));
OR2X2 OR2X2_1445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5369_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5662_));
OR2X2 OR2X2_1446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5663_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5664_));
OR2X2 OR2X2_1447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5665_));
OR2X2 OR2X2_1448 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5375_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5667_));
OR2X2 OR2X2_1449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_52_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5668_));
OR2X2 OR2X2_145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2636_));
OR2X2 OR2X2_1450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5670_), .B(AES_CORE_DATAPATH__abc_16009_new_n5671_), .Y(AES_CORE_DATAPATH__0key_2__31_0__20_));
OR2X2 OR2X2_1451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5381_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5673_));
OR2X2 OR2X2_1452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_53_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5674_));
OR2X2 OR2X2_1453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5675_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5676_));
OR2X2 OR2X2_1454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5677_));
OR2X2 OR2X2_1455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5387_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5679_));
OR2X2 OR2X2_1456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_54_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5680_));
OR2X2 OR2X2_1457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5681_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5682_));
OR2X2 OR2X2_1458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5683_));
OR2X2 OR2X2_1459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5393_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5685_));
OR2X2 OR2X2_146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2638_), .B(AES_CORE_DATAPATH__abc_16009_new_n2639_), .Y(\iv_out[15] ));
OR2X2 OR2X2_1460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_55_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5686_));
OR2X2 OR2X2_1461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5687_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5688_));
OR2X2 OR2X2_1462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5689_));
OR2X2 OR2X2_1463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5399_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5691_));
OR2X2 OR2X2_1464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_56_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5692_));
OR2X2 OR2X2_1465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5693_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5694_));
OR2X2 OR2X2_1466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5695_));
OR2X2 OR2X2_1467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5405_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5697_));
OR2X2 OR2X2_1468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_57_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5698_));
OR2X2 OR2X2_1469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5700_), .B(AES_CORE_DATAPATH__abc_16009_new_n5701_), .Y(AES_CORE_DATAPATH__0key_2__31_0__25_));
OR2X2 OR2X2_147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2643_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2644_));
OR2X2 OR2X2_1470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5411_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5703_));
OR2X2 OR2X2_1471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_58_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5704_));
OR2X2 OR2X2_1472 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5706_), .B(AES_CORE_DATAPATH__abc_16009_new_n5707_), .Y(AES_CORE_DATAPATH__0key_2__31_0__26_));
OR2X2 OR2X2_1473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5709_));
OR2X2 OR2X2_1474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_59_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5710_));
OR2X2 OR2X2_1475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5711_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5712_));
OR2X2 OR2X2_1476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5713_));
OR2X2 OR2X2_1477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_60_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5715_));
OR2X2 OR2X2_1478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5423_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5716_));
OR2X2 OR2X2_1479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5717_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5718_));
OR2X2 OR2X2_148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2644_), .B(AES_CORE_DATAPATH__abc_16009_new_n2642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2645_));
OR2X2 OR2X2_1480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5719_));
OR2X2 OR2X2_1481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5429_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5721_));
OR2X2 OR2X2_1482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_61_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5722_));
OR2X2 OR2X2_1483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5723_), .B(AES_CORE_DATAPATH__abc_16009_new_n5545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5724_));
OR2X2 OR2X2_1484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5550_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5725_));
OR2X2 OR2X2_1485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5435_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5727_));
OR2X2 OR2X2_1486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_62_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5728_));
OR2X2 OR2X2_1487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5730_), .B(AES_CORE_DATAPATH__abc_16009_new_n5731_), .Y(AES_CORE_DATAPATH__0key_2__31_0__30_));
OR2X2 OR2X2_1488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n5440_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5733_));
OR2X2 OR2X2_1489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_63_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5734_));
OR2X2 OR2X2_149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2646_));
OR2X2 OR2X2_1490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5736_), .B(AES_CORE_DATAPATH__abc_16009_new_n5737_), .Y(AES_CORE_DATAPATH__0key_2__31_0__31_));
OR2X2 OR2X2_1491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5741_), .B(AES_CORE_DATAPATH__abc_16009_new_n5742_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5743_));
OR2X2 OR2X2_1492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5745_), .B(AES_CORE_DATAPATH__abc_16009_new_n5746_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5747_));
OR2X2 OR2X2_1493 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5750_), .B(AES_CORE_DATAPATH__abc_16009_new_n5751_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5752_));
OR2X2 OR2X2_1494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5760_), .B(AES_CORE_DATAPATH__abc_16009_new_n5761_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5762_));
OR2X2 OR2X2_1495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5767_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5768_));
OR2X2 OR2X2_1496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5768_), .B(AES_CORE_DATAPATH__abc_16009_new_n5766_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5769_));
OR2X2 OR2X2_1497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5770_));
OR2X2 OR2X2_1498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5772_), .B(AES_CORE_DATAPATH__abc_16009_new_n5773_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5774_));
OR2X2 OR2X2_1499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5776_), .B(AES_CORE_DATAPATH__abc_16009_new_n5775_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5777_));
OR2X2 OR2X2_15 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT_state_4_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n138_));
OR2X2 OR2X2_150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2648_), .B(AES_CORE_DATAPATH__abc_16009_new_n2649_), .Y(\iv_out[16] ));
OR2X2 OR2X2_1500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5762_), .B(AES_CORE_DATAPATH__abc_16009_new_n5777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5778_));
OR2X2 OR2X2_1501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5781_), .B(AES_CORE_DATAPATH__abc_16009_new_n5782_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5783_));
OR2X2 OR2X2_1502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5783_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5784_));
OR2X2 OR2X2_1503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5786_), .B(AES_CORE_DATAPATH__abc_16009_new_n5787_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5788_));
OR2X2 OR2X2_1504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5789_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5790_));
OR2X2 OR2X2_1505 ( .A(\iv_out[0] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n5791_));
OR2X2 OR2X2_1506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5789_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5797_));
OR2X2 OR2X2_1507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5799_));
OR2X2 OR2X2_1508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5801_), .B(AES_CORE_DATAPATH__abc_16009_new_n5803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5804_));
OR2X2 OR2X2_1509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5804_), .B(AES_CORE_DATAPATH__abc_16009_new_n5795_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5805_));
OR2X2 OR2X2_151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2653_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2654_));
OR2X2 OR2X2_1510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5806_), .B(AES_CORE_DATAPATH__abc_16009_new_n5755_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5807_));
OR2X2 OR2X2_1511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5807_), .B(AES_CORE_DATAPATH__abc_16009_new_n5753_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5808_));
OR2X2 OR2X2_1512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5809_), .B(AES_CORE_DATAPATH__abc_16009_new_n5740_), .Y(AES_CORE_DATAPATH__0col_0__31_0__0_));
OR2X2 OR2X2_1513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5812_), .B(AES_CORE_DATAPATH__abc_16009_new_n5813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5814_));
OR2X2 OR2X2_1514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5818_), .B(AES_CORE_DATAPATH__abc_16009_new_n5819_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5820_));
OR2X2 OR2X2_1515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5822_));
OR2X2 OR2X2_1516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5821_), .B(AES_CORE_DATAPATH__abc_16009_new_n5823_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5824_));
OR2X2 OR2X2_1517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5827_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5828_));
OR2X2 OR2X2_1518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5828_), .B(AES_CORE_DATAPATH__abc_16009_new_n5826_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5829_));
OR2X2 OR2X2_1519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5830_));
OR2X2 OR2X2_152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2654_), .B(AES_CORE_DATAPATH__abc_16009_new_n2652_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2655_));
OR2X2 OR2X2_1520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5832_), .B(AES_CORE_DATAPATH__abc_16009_new_n5833_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5834_));
OR2X2 OR2X2_1521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5834_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5835_));
OR2X2 OR2X2_1522 ( .A(\iv_out[1] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5836_));
OR2X2 OR2X2_1523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5824_), .B(AES_CORE_DATAPATH__abc_16009_new_n5838_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5839_));
OR2X2 OR2X2_1524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3496_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5840_));
OR2X2 OR2X2_1525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5841_), .B(AES_CORE_DATAPATH__abc_16009_new_n5837_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5842_));
OR2X2 OR2X2_1526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5843_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5844_));
OR2X2 OR2X2_1527 ( .A(\iv_out[1] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n5845_));
OR2X2 OR2X2_1528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5843_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5848_));
OR2X2 OR2X2_1529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5849_));
OR2X2 OR2X2_153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2656_));
OR2X2 OR2X2_1530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5851_), .B(AES_CORE_DATAPATH__abc_16009_new_n5852_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5853_));
OR2X2 OR2X2_1531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5853_), .B(AES_CORE_DATAPATH__abc_16009_new_n5847_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5854_));
OR2X2 OR2X2_1532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5855_), .B(AES_CORE_DATAPATH__abc_16009_new_n5856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5857_));
OR2X2 OR2X2_1533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5857_), .B(AES_CORE_DATAPATH__abc_16009_new_n5815_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5858_));
OR2X2 OR2X2_1534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5859_), .B(AES_CORE_DATAPATH__abc_16009_new_n5811_), .Y(AES_CORE_DATAPATH__0col_0__31_0__1_));
OR2X2 OR2X2_1535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5862_), .B(AES_CORE_DATAPATH__abc_16009_new_n5863_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5864_));
OR2X2 OR2X2_1536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5866_), .B(AES_CORE_DATAPATH__abc_16009_new_n5867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5868_));
OR2X2 OR2X2_1537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5871_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5872_));
OR2X2 OR2X2_1538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5872_), .B(AES_CORE_DATAPATH__abc_16009_new_n5870_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5873_));
OR2X2 OR2X2_1539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5874_));
OR2X2 OR2X2_154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2658_), .B(AES_CORE_DATAPATH__abc_16009_new_n2659_), .Y(\iv_out[17] ));
OR2X2 OR2X2_1540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5876_), .B(AES_CORE_DATAPATH__abc_16009_new_n5877_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5878_));
OR2X2 OR2X2_1541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5878_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5879_));
OR2X2 OR2X2_1542 ( .A(\iv_out[2] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5880_));
OR2X2 OR2X2_1543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5868_), .B(AES_CORE_DATAPATH__abc_16009_new_n5881_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5882_));
OR2X2 OR2X2_1544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5885_), .B(AES_CORE_DATAPATH__abc_16009_new_n5886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5887_));
OR2X2 OR2X2_1545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5887_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5888_));
OR2X2 OR2X2_1546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5890_), .B(AES_CORE_DATAPATH__abc_16009_new_n5891_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5892_));
OR2X2 OR2X2_1547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5893_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5894_));
OR2X2 OR2X2_1548 ( .A(\iv_out[2] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n5895_));
OR2X2 OR2X2_1549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5893_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5898_));
OR2X2 OR2X2_155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2663_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2664_));
OR2X2 OR2X2_1550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5899_));
OR2X2 OR2X2_1551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5901_), .B(AES_CORE_DATAPATH__abc_16009_new_n5902_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5903_));
OR2X2 OR2X2_1552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5903_), .B(AES_CORE_DATAPATH__abc_16009_new_n5897_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5904_));
OR2X2 OR2X2_1553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5905_), .B(AES_CORE_DATAPATH__abc_16009_new_n5906_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5907_));
OR2X2 OR2X2_1554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5907_), .B(AES_CORE_DATAPATH__abc_16009_new_n5865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5908_));
OR2X2 OR2X2_1555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5909_), .B(AES_CORE_DATAPATH__abc_16009_new_n5861_), .Y(AES_CORE_DATAPATH__0col_0__31_0__2_));
OR2X2 OR2X2_1556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5912_), .B(AES_CORE_DATAPATH__abc_16009_new_n5913_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5914_));
OR2X2 OR2X2_1557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5918_), .B(AES_CORE_DATAPATH__abc_16009_new_n5919_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5920_));
OR2X2 OR2X2_1558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5922_));
OR2X2 OR2X2_1559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5921_), .B(AES_CORE_DATAPATH__abc_16009_new_n5923_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5924_));
OR2X2 OR2X2_156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2664_), .B(AES_CORE_DATAPATH__abc_16009_new_n2662_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2665_));
OR2X2 OR2X2_1560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5927_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5928_));
OR2X2 OR2X2_1561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5928_), .B(AES_CORE_DATAPATH__abc_16009_new_n5926_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5929_));
OR2X2 OR2X2_1562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5930_));
OR2X2 OR2X2_1563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5932_), .B(AES_CORE_DATAPATH__abc_16009_new_n5933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5934_));
OR2X2 OR2X2_1564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5934_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5935_));
OR2X2 OR2X2_1565 ( .A(\iv_out[3] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5936_));
OR2X2 OR2X2_1566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5924_), .B(AES_CORE_DATAPATH__abc_16009_new_n5938_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5939_));
OR2X2 OR2X2_1567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3560_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5940_));
OR2X2 OR2X2_1568 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5941_), .B(AES_CORE_DATAPATH__abc_16009_new_n5937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5942_));
OR2X2 OR2X2_1569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5943_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5944_));
OR2X2 OR2X2_157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2666_));
OR2X2 OR2X2_1570 ( .A(\iv_out[3] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n5945_));
OR2X2 OR2X2_1571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5943_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5948_));
OR2X2 OR2X2_1572 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5949_));
OR2X2 OR2X2_1573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5951_), .B(AES_CORE_DATAPATH__abc_16009_new_n5952_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5953_));
OR2X2 OR2X2_1574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5953_), .B(AES_CORE_DATAPATH__abc_16009_new_n5947_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5954_));
OR2X2 OR2X2_1575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5955_), .B(AES_CORE_DATAPATH__abc_16009_new_n5956_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5957_));
OR2X2 OR2X2_1576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5957_), .B(AES_CORE_DATAPATH__abc_16009_new_n5915_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5958_));
OR2X2 OR2X2_1577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5959_), .B(AES_CORE_DATAPATH__abc_16009_new_n5911_), .Y(AES_CORE_DATAPATH__0col_0__31_0__3_));
OR2X2 OR2X2_1578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5962_), .B(AES_CORE_DATAPATH__abc_16009_new_n5963_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5964_));
OR2X2 OR2X2_1579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5966_), .B(AES_CORE_DATAPATH__abc_16009_new_n5967_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5968_));
OR2X2 OR2X2_158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2668_), .B(AES_CORE_DATAPATH__abc_16009_new_n2669_), .Y(\iv_out[18] ));
OR2X2 OR2X2_1580 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5971_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5972_));
OR2X2 OR2X2_1581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5972_), .B(AES_CORE_DATAPATH__abc_16009_new_n5970_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5973_));
OR2X2 OR2X2_1582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5974_));
OR2X2 OR2X2_1583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5976_), .B(AES_CORE_DATAPATH__abc_16009_new_n5977_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5978_));
OR2X2 OR2X2_1584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5978_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5979_));
OR2X2 OR2X2_1585 ( .A(\iv_out[4] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5980_));
OR2X2 OR2X2_1586 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5968_), .B(AES_CORE_DATAPATH__abc_16009_new_n5981_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5982_));
OR2X2 OR2X2_1587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5985_), .B(AES_CORE_DATAPATH__abc_16009_new_n5986_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5987_));
OR2X2 OR2X2_1588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5987_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5988_));
OR2X2 OR2X2_1589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5990_), .B(AES_CORE_DATAPATH__abc_16009_new_n5991_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5992_));
OR2X2 OR2X2_159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2673_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2674_));
OR2X2 OR2X2_1590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5993_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5994_));
OR2X2 OR2X2_1591 ( .A(\iv_out[4] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n5995_));
OR2X2 OR2X2_1592 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5993_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5998_));
OR2X2 OR2X2_1593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n5999_));
OR2X2 OR2X2_1594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6001_), .B(AES_CORE_DATAPATH__abc_16009_new_n6002_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6003_));
OR2X2 OR2X2_1595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6003_), .B(AES_CORE_DATAPATH__abc_16009_new_n5997_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6004_));
OR2X2 OR2X2_1596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6005_), .B(AES_CORE_DATAPATH__abc_16009_new_n6006_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6007_));
OR2X2 OR2X2_1597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6007_), .B(AES_CORE_DATAPATH__abc_16009_new_n5965_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6008_));
OR2X2 OR2X2_1598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6009_), .B(AES_CORE_DATAPATH__abc_16009_new_n5961_), .Y(AES_CORE_DATAPATH__0col_0__31_0__4_));
OR2X2 OR2X2_1599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6012_), .B(AES_CORE_DATAPATH__abc_16009_new_n6013_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6014_));
OR2X2 OR2X2_16 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n138_), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n139_));
OR2X2 OR2X2_160 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2674_), .B(AES_CORE_DATAPATH__abc_16009_new_n2672_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2675_));
OR2X2 OR2X2_1600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6016_), .B(AES_CORE_DATAPATH__abc_16009_new_n6017_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6018_));
OR2X2 OR2X2_1601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6021_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6022_));
OR2X2 OR2X2_1602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6022_), .B(AES_CORE_DATAPATH__abc_16009_new_n6020_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6023_));
OR2X2 OR2X2_1603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6024_));
OR2X2 OR2X2_1604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6026_), .B(AES_CORE_DATAPATH__abc_16009_new_n6027_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6028_));
OR2X2 OR2X2_1605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6028_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6029_));
OR2X2 OR2X2_1606 ( .A(\iv_out[5] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6030_));
OR2X2 OR2X2_1607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6018_), .B(AES_CORE_DATAPATH__abc_16009_new_n6031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6032_));
OR2X2 OR2X2_1608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6035_), .B(AES_CORE_DATAPATH__abc_16009_new_n6036_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6037_));
OR2X2 OR2X2_1609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6037_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6038_));
OR2X2 OR2X2_161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2676_));
OR2X2 OR2X2_1610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6040_), .B(AES_CORE_DATAPATH__abc_16009_new_n6041_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6042_));
OR2X2 OR2X2_1611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6043_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6044_));
OR2X2 OR2X2_1612 ( .A(\iv_out[5] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6045_));
OR2X2 OR2X2_1613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6043_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6048_));
OR2X2 OR2X2_1614 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6049_));
OR2X2 OR2X2_1615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6051_), .B(AES_CORE_DATAPATH__abc_16009_new_n6052_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6053_));
OR2X2 OR2X2_1616 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6053_), .B(AES_CORE_DATAPATH__abc_16009_new_n6047_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6054_));
OR2X2 OR2X2_1617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6055_), .B(AES_CORE_DATAPATH__abc_16009_new_n6056_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6057_));
OR2X2 OR2X2_1618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6057_), .B(AES_CORE_DATAPATH__abc_16009_new_n6015_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6058_));
OR2X2 OR2X2_1619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6059_), .B(AES_CORE_DATAPATH__abc_16009_new_n6011_), .Y(AES_CORE_DATAPATH__0col_0__31_0__5_));
OR2X2 OR2X2_162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2678_), .B(AES_CORE_DATAPATH__abc_16009_new_n2679_), .Y(\iv_out[19] ));
OR2X2 OR2X2_1620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6062_), .B(AES_CORE_DATAPATH__abc_16009_new_n6063_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6064_));
OR2X2 OR2X2_1621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6066_), .B(AES_CORE_DATAPATH__abc_16009_new_n6067_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6068_));
OR2X2 OR2X2_1622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6071_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6072_));
OR2X2 OR2X2_1623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6072_), .B(AES_CORE_DATAPATH__abc_16009_new_n6070_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6073_));
OR2X2 OR2X2_1624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6074_));
OR2X2 OR2X2_1625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6076_), .B(AES_CORE_DATAPATH__abc_16009_new_n6077_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6078_));
OR2X2 OR2X2_1626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6078_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6079_));
OR2X2 OR2X2_1627 ( .A(\iv_out[6] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6080_));
OR2X2 OR2X2_1628 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6068_), .B(AES_CORE_DATAPATH__abc_16009_new_n6081_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6082_));
OR2X2 OR2X2_1629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6085_), .B(AES_CORE_DATAPATH__abc_16009_new_n6086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6087_));
OR2X2 OR2X2_163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2683_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2684_));
OR2X2 OR2X2_1630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6087_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6088_));
OR2X2 OR2X2_1631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6090_), .B(AES_CORE_DATAPATH__abc_16009_new_n6091_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6092_));
OR2X2 OR2X2_1632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6093_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6094_));
OR2X2 OR2X2_1633 ( .A(\iv_out[6] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6095_));
OR2X2 OR2X2_1634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6093_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6098_));
OR2X2 OR2X2_1635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6099_));
OR2X2 OR2X2_1636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6101_), .B(AES_CORE_DATAPATH__abc_16009_new_n6102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6103_));
OR2X2 OR2X2_1637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6103_), .B(AES_CORE_DATAPATH__abc_16009_new_n6097_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6104_));
OR2X2 OR2X2_1638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6105_), .B(AES_CORE_DATAPATH__abc_16009_new_n6106_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6107_));
OR2X2 OR2X2_1639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6107_), .B(AES_CORE_DATAPATH__abc_16009_new_n6065_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6108_));
OR2X2 OR2X2_164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2684_), .B(AES_CORE_DATAPATH__abc_16009_new_n2682_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2685_));
OR2X2 OR2X2_1640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6109_), .B(AES_CORE_DATAPATH__abc_16009_new_n6061_), .Y(AES_CORE_DATAPATH__0col_0__31_0__6_));
OR2X2 OR2X2_1641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6112_), .B(AES_CORE_DATAPATH__abc_16009_new_n6113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6114_));
OR2X2 OR2X2_1642 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6118_), .B(AES_CORE_DATAPATH__abc_16009_new_n6119_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6120_));
OR2X2 OR2X2_1643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6122_));
OR2X2 OR2X2_1644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6121_), .B(AES_CORE_DATAPATH__abc_16009_new_n6123_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6124_));
OR2X2 OR2X2_1645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6127_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6128_));
OR2X2 OR2X2_1646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6128_), .B(AES_CORE_DATAPATH__abc_16009_new_n6126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6129_));
OR2X2 OR2X2_1647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6130_));
OR2X2 OR2X2_1648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6132_), .B(AES_CORE_DATAPATH__abc_16009_new_n6133_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6134_));
OR2X2 OR2X2_1649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6134_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6135_));
OR2X2 OR2X2_165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2686_));
OR2X2 OR2X2_1650 ( .A(\iv_out[7] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6136_));
OR2X2 OR2X2_1651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6124_), .B(AES_CORE_DATAPATH__abc_16009_new_n6138_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6139_));
OR2X2 OR2X2_1652 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3688_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6140_));
OR2X2 OR2X2_1653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6141_), .B(AES_CORE_DATAPATH__abc_16009_new_n6137_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6142_));
OR2X2 OR2X2_1654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6143_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6144_));
OR2X2 OR2X2_1655 ( .A(\iv_out[7] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6145_));
OR2X2 OR2X2_1656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6143_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6148_));
OR2X2 OR2X2_1657 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6149_));
OR2X2 OR2X2_1658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6151_), .B(AES_CORE_DATAPATH__abc_16009_new_n6152_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6153_));
OR2X2 OR2X2_1659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6153_), .B(AES_CORE_DATAPATH__abc_16009_new_n6147_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6154_));
OR2X2 OR2X2_166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2688_), .B(AES_CORE_DATAPATH__abc_16009_new_n2689_), .Y(\iv_out[20] ));
OR2X2 OR2X2_1660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6155_), .B(AES_CORE_DATAPATH__abc_16009_new_n6156_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6157_));
OR2X2 OR2X2_1661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6157_), .B(AES_CORE_DATAPATH__abc_16009_new_n6115_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6158_));
OR2X2 OR2X2_1662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6159_), .B(AES_CORE_DATAPATH__abc_16009_new_n6111_), .Y(AES_CORE_DATAPATH__0col_0__31_0__7_));
OR2X2 OR2X2_1663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6162_), .B(AES_CORE_DATAPATH__abc_16009_new_n6163_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6164_));
OR2X2 OR2X2_1664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6166_), .B(AES_CORE_DATAPATH__abc_16009_new_n6167_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6168_));
OR2X2 OR2X2_1665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6171_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6172_));
OR2X2 OR2X2_1666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6172_), .B(AES_CORE_DATAPATH__abc_16009_new_n6170_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6173_));
OR2X2 OR2X2_1667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6174_));
OR2X2 OR2X2_1668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6176_), .B(AES_CORE_DATAPATH__abc_16009_new_n6177_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6178_));
OR2X2 OR2X2_1669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6178_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6179_));
OR2X2 OR2X2_167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2693_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2694_));
OR2X2 OR2X2_1670 ( .A(\iv_out[8] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6180_));
OR2X2 OR2X2_1671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6168_), .B(AES_CORE_DATAPATH__abc_16009_new_n6181_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6182_));
OR2X2 OR2X2_1672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6185_), .B(AES_CORE_DATAPATH__abc_16009_new_n6186_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6187_));
OR2X2 OR2X2_1673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6187_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6188_));
OR2X2 OR2X2_1674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6190_), .B(AES_CORE_DATAPATH__abc_16009_new_n6191_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6192_));
OR2X2 OR2X2_1675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6193_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6194_));
OR2X2 OR2X2_1676 ( .A(\iv_out[8] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6195_));
OR2X2 OR2X2_1677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6193_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6198_));
OR2X2 OR2X2_1678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6199_));
OR2X2 OR2X2_1679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6201_), .B(AES_CORE_DATAPATH__abc_16009_new_n6202_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6203_));
OR2X2 OR2X2_168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2694_), .B(AES_CORE_DATAPATH__abc_16009_new_n2692_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2695_));
OR2X2 OR2X2_1680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6203_), .B(AES_CORE_DATAPATH__abc_16009_new_n6197_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6204_));
OR2X2 OR2X2_1681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6205_), .B(AES_CORE_DATAPATH__abc_16009_new_n6206_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6207_));
OR2X2 OR2X2_1682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6207_), .B(AES_CORE_DATAPATH__abc_16009_new_n6165_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6208_));
OR2X2 OR2X2_1683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6209_), .B(AES_CORE_DATAPATH__abc_16009_new_n6161_), .Y(AES_CORE_DATAPATH__0col_0__31_0__8_));
OR2X2 OR2X2_1684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6212_), .B(AES_CORE_DATAPATH__abc_16009_new_n6213_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6214_));
OR2X2 OR2X2_1685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6218_), .B(AES_CORE_DATAPATH__abc_16009_new_n6219_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6220_));
OR2X2 OR2X2_1686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6222_));
OR2X2 OR2X2_1687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6221_), .B(AES_CORE_DATAPATH__abc_16009_new_n6223_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6224_));
OR2X2 OR2X2_1688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6227_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6228_));
OR2X2 OR2X2_1689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6228_), .B(AES_CORE_DATAPATH__abc_16009_new_n6226_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6229_));
OR2X2 OR2X2_169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2696_));
OR2X2 OR2X2_1690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6230_));
OR2X2 OR2X2_1691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6232_), .B(AES_CORE_DATAPATH__abc_16009_new_n6233_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6234_));
OR2X2 OR2X2_1692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6234_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6235_));
OR2X2 OR2X2_1693 ( .A(\iv_out[9] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6236_));
OR2X2 OR2X2_1694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6224_), .B(AES_CORE_DATAPATH__abc_16009_new_n6238_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6239_));
OR2X2 OR2X2_1695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3752_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6240_));
OR2X2 OR2X2_1696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6241_), .B(AES_CORE_DATAPATH__abc_16009_new_n6237_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6242_));
OR2X2 OR2X2_1697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6243_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6244_));
OR2X2 OR2X2_1698 ( .A(\iv_out[9] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6245_));
OR2X2 OR2X2_1699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6243_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6248_));
OR2X2 OR2X2_17 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n139_), .B(AES_CORE_CONTROL_UNIT_state_8_), .Y(AES_CORE_CONTROL_UNIT_bypass_rk));
OR2X2 OR2X2_170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2698_), .B(AES_CORE_DATAPATH__abc_16009_new_n2699_), .Y(\iv_out[21] ));
OR2X2 OR2X2_1700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6249_));
OR2X2 OR2X2_1701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6251_), .B(AES_CORE_DATAPATH__abc_16009_new_n6252_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6253_));
OR2X2 OR2X2_1702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6253_), .B(AES_CORE_DATAPATH__abc_16009_new_n6247_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6254_));
OR2X2 OR2X2_1703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6255_), .B(AES_CORE_DATAPATH__abc_16009_new_n6256_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6257_));
OR2X2 OR2X2_1704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6257_), .B(AES_CORE_DATAPATH__abc_16009_new_n6215_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6258_));
OR2X2 OR2X2_1705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6259_), .B(AES_CORE_DATAPATH__abc_16009_new_n6211_), .Y(AES_CORE_DATAPATH__0col_0__31_0__9_));
OR2X2 OR2X2_1706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6262_), .B(AES_CORE_DATAPATH__abc_16009_new_n6263_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6264_));
OR2X2 OR2X2_1707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6266_), .B(AES_CORE_DATAPATH__abc_16009_new_n6267_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6268_));
OR2X2 OR2X2_1708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6271_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6272_));
OR2X2 OR2X2_1709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6272_), .B(AES_CORE_DATAPATH__abc_16009_new_n6270_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6273_));
OR2X2 OR2X2_171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2703_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2704_));
OR2X2 OR2X2_1710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6274_));
OR2X2 OR2X2_1711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6276_), .B(AES_CORE_DATAPATH__abc_16009_new_n6277_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6278_));
OR2X2 OR2X2_1712 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6278_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6279_));
OR2X2 OR2X2_1713 ( .A(\iv_out[10] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6280_));
OR2X2 OR2X2_1714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6268_), .B(AES_CORE_DATAPATH__abc_16009_new_n6281_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6282_));
OR2X2 OR2X2_1715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6285_), .B(AES_CORE_DATAPATH__abc_16009_new_n6286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6287_));
OR2X2 OR2X2_1716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6287_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6288_));
OR2X2 OR2X2_1717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6290_), .B(AES_CORE_DATAPATH__abc_16009_new_n6291_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6292_));
OR2X2 OR2X2_1718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6293_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6294_));
OR2X2 OR2X2_1719 ( .A(\iv_out[10] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6295_));
OR2X2 OR2X2_172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2704_), .B(AES_CORE_DATAPATH__abc_16009_new_n2702_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2705_));
OR2X2 OR2X2_1720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6293_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6298_));
OR2X2 OR2X2_1721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6299_));
OR2X2 OR2X2_1722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6301_), .B(AES_CORE_DATAPATH__abc_16009_new_n6302_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6303_));
OR2X2 OR2X2_1723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6303_), .B(AES_CORE_DATAPATH__abc_16009_new_n6297_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6304_));
OR2X2 OR2X2_1724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6305_), .B(AES_CORE_DATAPATH__abc_16009_new_n6306_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6307_));
OR2X2 OR2X2_1725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6307_), .B(AES_CORE_DATAPATH__abc_16009_new_n6265_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6308_));
OR2X2 OR2X2_1726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6309_), .B(AES_CORE_DATAPATH__abc_16009_new_n6261_), .Y(AES_CORE_DATAPATH__0col_0__31_0__10_));
OR2X2 OR2X2_1727 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6312_), .B(AES_CORE_DATAPATH__abc_16009_new_n6313_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6314_));
OR2X2 OR2X2_1728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6318_), .B(AES_CORE_DATAPATH__abc_16009_new_n6319_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6320_));
OR2X2 OR2X2_1729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6322_));
OR2X2 OR2X2_173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2706_));
OR2X2 OR2X2_1730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6321_), .B(AES_CORE_DATAPATH__abc_16009_new_n6323_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6324_));
OR2X2 OR2X2_1731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6327_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6328_));
OR2X2 OR2X2_1732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6328_), .B(AES_CORE_DATAPATH__abc_16009_new_n6326_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6329_));
OR2X2 OR2X2_1733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6330_));
OR2X2 OR2X2_1734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6332_), .B(AES_CORE_DATAPATH__abc_16009_new_n6333_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6334_));
OR2X2 OR2X2_1735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6334_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6335_));
OR2X2 OR2X2_1736 ( .A(\iv_out[11] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6336_));
OR2X2 OR2X2_1737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6324_), .B(AES_CORE_DATAPATH__abc_16009_new_n6338_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6339_));
OR2X2 OR2X2_1738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3816_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6340_));
OR2X2 OR2X2_1739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6341_), .B(AES_CORE_DATAPATH__abc_16009_new_n6337_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6342_));
OR2X2 OR2X2_174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2708_), .B(AES_CORE_DATAPATH__abc_16009_new_n2709_), .Y(\iv_out[22] ));
OR2X2 OR2X2_1740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6343_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6344_));
OR2X2 OR2X2_1741 ( .A(\iv_out[11] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6345_));
OR2X2 OR2X2_1742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6343_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6348_));
OR2X2 OR2X2_1743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6349_));
OR2X2 OR2X2_1744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6351_), .B(AES_CORE_DATAPATH__abc_16009_new_n6352_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6353_));
OR2X2 OR2X2_1745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6353_), .B(AES_CORE_DATAPATH__abc_16009_new_n6347_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6354_));
OR2X2 OR2X2_1746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6355_), .B(AES_CORE_DATAPATH__abc_16009_new_n6356_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6357_));
OR2X2 OR2X2_1747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6357_), .B(AES_CORE_DATAPATH__abc_16009_new_n6315_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6358_));
OR2X2 OR2X2_1748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6359_), .B(AES_CORE_DATAPATH__abc_16009_new_n6311_), .Y(AES_CORE_DATAPATH__0col_0__31_0__11_));
OR2X2 OR2X2_1749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6362_), .B(AES_CORE_DATAPATH__abc_16009_new_n6363_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6364_));
OR2X2 OR2X2_175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2713_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2714_));
OR2X2 OR2X2_1750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6366_), .B(AES_CORE_DATAPATH__abc_16009_new_n6367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6368_));
OR2X2 OR2X2_1751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6371_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6372_));
OR2X2 OR2X2_1752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6372_), .B(AES_CORE_DATAPATH__abc_16009_new_n6370_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6373_));
OR2X2 OR2X2_1753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6374_));
OR2X2 OR2X2_1754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6376_), .B(AES_CORE_DATAPATH__abc_16009_new_n6377_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6378_));
OR2X2 OR2X2_1755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6378_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6379_));
OR2X2 OR2X2_1756 ( .A(\iv_out[12] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6380_));
OR2X2 OR2X2_1757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6368_), .B(AES_CORE_DATAPATH__abc_16009_new_n6381_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6382_));
OR2X2 OR2X2_1758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6385_), .B(AES_CORE_DATAPATH__abc_16009_new_n6386_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6387_));
OR2X2 OR2X2_1759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6387_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6388_));
OR2X2 OR2X2_176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2714_), .B(AES_CORE_DATAPATH__abc_16009_new_n2712_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2715_));
OR2X2 OR2X2_1760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6390_), .B(AES_CORE_DATAPATH__abc_16009_new_n6391_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6392_));
OR2X2 OR2X2_1761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6393_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6394_));
OR2X2 OR2X2_1762 ( .A(\iv_out[12] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6395_));
OR2X2 OR2X2_1763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6393_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6398_));
OR2X2 OR2X2_1764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6399_));
OR2X2 OR2X2_1765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6401_), .B(AES_CORE_DATAPATH__abc_16009_new_n6402_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6403_));
OR2X2 OR2X2_1766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6403_), .B(AES_CORE_DATAPATH__abc_16009_new_n6397_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6404_));
OR2X2 OR2X2_1767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6405_), .B(AES_CORE_DATAPATH__abc_16009_new_n6406_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6407_));
OR2X2 OR2X2_1768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6407_), .B(AES_CORE_DATAPATH__abc_16009_new_n6365_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6408_));
OR2X2 OR2X2_1769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6409_), .B(AES_CORE_DATAPATH__abc_16009_new_n6361_), .Y(AES_CORE_DATAPATH__0col_0__31_0__12_));
OR2X2 OR2X2_177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2716_));
OR2X2 OR2X2_1770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6412_), .B(AES_CORE_DATAPATH__abc_16009_new_n6413_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6414_));
OR2X2 OR2X2_1771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6418_), .B(AES_CORE_DATAPATH__abc_16009_new_n6419_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6420_));
OR2X2 OR2X2_1772 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6422_));
OR2X2 OR2X2_1773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6421_), .B(AES_CORE_DATAPATH__abc_16009_new_n6423_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6424_));
OR2X2 OR2X2_1774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6427_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6428_));
OR2X2 OR2X2_1775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6428_), .B(AES_CORE_DATAPATH__abc_16009_new_n6426_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6429_));
OR2X2 OR2X2_1776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6430_));
OR2X2 OR2X2_1777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6432_), .B(AES_CORE_DATAPATH__abc_16009_new_n6433_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6434_));
OR2X2 OR2X2_1778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6434_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6435_));
OR2X2 OR2X2_1779 ( .A(\iv_out[13] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6436_));
OR2X2 OR2X2_178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2718_), .B(AES_CORE_DATAPATH__abc_16009_new_n2719_), .Y(\iv_out[23] ));
OR2X2 OR2X2_1780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6424_), .B(AES_CORE_DATAPATH__abc_16009_new_n6438_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6439_));
OR2X2 OR2X2_1781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3880_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6440_));
OR2X2 OR2X2_1782 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6441_), .B(AES_CORE_DATAPATH__abc_16009_new_n6437_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6442_));
OR2X2 OR2X2_1783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6443_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6444_));
OR2X2 OR2X2_1784 ( .A(\iv_out[13] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6445_));
OR2X2 OR2X2_1785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6443_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6448_));
OR2X2 OR2X2_1786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6449_));
OR2X2 OR2X2_1787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6451_), .B(AES_CORE_DATAPATH__abc_16009_new_n6452_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6453_));
OR2X2 OR2X2_1788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6453_), .B(AES_CORE_DATAPATH__abc_16009_new_n6447_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6454_));
OR2X2 OR2X2_1789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6455_), .B(AES_CORE_DATAPATH__abc_16009_new_n6456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6457_));
OR2X2 OR2X2_179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2723_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2724_));
OR2X2 OR2X2_1790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6457_), .B(AES_CORE_DATAPATH__abc_16009_new_n6415_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6458_));
OR2X2 OR2X2_1791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6459_), .B(AES_CORE_DATAPATH__abc_16009_new_n6411_), .Y(AES_CORE_DATAPATH__0col_0__31_0__13_));
OR2X2 OR2X2_1792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6462_), .B(AES_CORE_DATAPATH__abc_16009_new_n6463_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6464_));
OR2X2 OR2X2_1793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6466_), .B(AES_CORE_DATAPATH__abc_16009_new_n6467_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6468_));
OR2X2 OR2X2_1794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6471_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6472_));
OR2X2 OR2X2_1795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6472_), .B(AES_CORE_DATAPATH__abc_16009_new_n6470_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6473_));
OR2X2 OR2X2_1796 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6474_));
OR2X2 OR2X2_1797 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6476_), .B(AES_CORE_DATAPATH__abc_16009_new_n6477_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6478_));
OR2X2 OR2X2_1798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6478_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6479_));
OR2X2 OR2X2_1799 ( .A(\iv_out[14] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6480_));
OR2X2 OR2X2_18 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n144_));
OR2X2 OR2X2_180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2724_), .B(AES_CORE_DATAPATH__abc_16009_new_n2722_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2725_));
OR2X2 OR2X2_1800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6468_), .B(AES_CORE_DATAPATH__abc_16009_new_n6481_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6482_));
OR2X2 OR2X2_1801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6485_), .B(AES_CORE_DATAPATH__abc_16009_new_n6486_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6487_));
OR2X2 OR2X2_1802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6487_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6488_));
OR2X2 OR2X2_1803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6490_), .B(AES_CORE_DATAPATH__abc_16009_new_n6491_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6492_));
OR2X2 OR2X2_1804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6493_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6494_));
OR2X2 OR2X2_1805 ( .A(\iv_out[14] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6495_));
OR2X2 OR2X2_1806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6493_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6498_));
OR2X2 OR2X2_1807 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6499_));
OR2X2 OR2X2_1808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6501_), .B(AES_CORE_DATAPATH__abc_16009_new_n6502_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6503_));
OR2X2 OR2X2_1809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6503_), .B(AES_CORE_DATAPATH__abc_16009_new_n6497_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6504_));
OR2X2 OR2X2_181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2726_));
OR2X2 OR2X2_1810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6505_), .B(AES_CORE_DATAPATH__abc_16009_new_n6506_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6507_));
OR2X2 OR2X2_1811 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6507_), .B(AES_CORE_DATAPATH__abc_16009_new_n6465_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6508_));
OR2X2 OR2X2_1812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6509_), .B(AES_CORE_DATAPATH__abc_16009_new_n6461_), .Y(AES_CORE_DATAPATH__0col_0__31_0__14_));
OR2X2 OR2X2_1813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6512_), .B(AES_CORE_DATAPATH__abc_16009_new_n6513_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6514_));
OR2X2 OR2X2_1814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6518_), .B(AES_CORE_DATAPATH__abc_16009_new_n6519_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6520_));
OR2X2 OR2X2_1815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6522_));
OR2X2 OR2X2_1816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6521_), .B(AES_CORE_DATAPATH__abc_16009_new_n6523_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6524_));
OR2X2 OR2X2_1817 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6527_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6528_));
OR2X2 OR2X2_1818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6528_), .B(AES_CORE_DATAPATH__abc_16009_new_n6526_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6529_));
OR2X2 OR2X2_1819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6530_));
OR2X2 OR2X2_182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2728_), .B(AES_CORE_DATAPATH__abc_16009_new_n2729_), .Y(\iv_out[24] ));
OR2X2 OR2X2_1820 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6532_), .B(AES_CORE_DATAPATH__abc_16009_new_n6533_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6534_));
OR2X2 OR2X2_1821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6534_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6535_));
OR2X2 OR2X2_1822 ( .A(\iv_out[15] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6536_));
OR2X2 OR2X2_1823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6524_), .B(AES_CORE_DATAPATH__abc_16009_new_n6538_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6539_));
OR2X2 OR2X2_1824 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3944_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6540_));
OR2X2 OR2X2_1825 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6541_), .B(AES_CORE_DATAPATH__abc_16009_new_n6537_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6542_));
OR2X2 OR2X2_1826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6543_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6544_));
OR2X2 OR2X2_1827 ( .A(\iv_out[15] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6545_));
OR2X2 OR2X2_1828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6543_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6548_));
OR2X2 OR2X2_1829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6549_));
OR2X2 OR2X2_183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2733_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2734_));
OR2X2 OR2X2_1830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6551_), .B(AES_CORE_DATAPATH__abc_16009_new_n6552_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6553_));
OR2X2 OR2X2_1831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6553_), .B(AES_CORE_DATAPATH__abc_16009_new_n6547_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6554_));
OR2X2 OR2X2_1832 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6555_), .B(AES_CORE_DATAPATH__abc_16009_new_n6556_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6557_));
OR2X2 OR2X2_1833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6557_), .B(AES_CORE_DATAPATH__abc_16009_new_n6515_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6558_));
OR2X2 OR2X2_1834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6559_), .B(AES_CORE_DATAPATH__abc_16009_new_n6511_), .Y(AES_CORE_DATAPATH__0col_0__31_0__15_));
OR2X2 OR2X2_1835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6562_), .B(AES_CORE_DATAPATH__abc_16009_new_n6563_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6564_));
OR2X2 OR2X2_1836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6566_), .B(AES_CORE_DATAPATH__abc_16009_new_n6567_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6568_));
OR2X2 OR2X2_1837 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6571_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6572_));
OR2X2 OR2X2_1838 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6572_), .B(AES_CORE_DATAPATH__abc_16009_new_n6570_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6573_));
OR2X2 OR2X2_1839 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6574_));
OR2X2 OR2X2_184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2734_), .B(AES_CORE_DATAPATH__abc_16009_new_n2732_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2735_));
OR2X2 OR2X2_1840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6576_), .B(AES_CORE_DATAPATH__abc_16009_new_n6577_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6578_));
OR2X2 OR2X2_1841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6578_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6579_));
OR2X2 OR2X2_1842 ( .A(\iv_out[16] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6580_));
OR2X2 OR2X2_1843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6568_), .B(AES_CORE_DATAPATH__abc_16009_new_n6581_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6582_));
OR2X2 OR2X2_1844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6585_), .B(AES_CORE_DATAPATH__abc_16009_new_n6586_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6587_));
OR2X2 OR2X2_1845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6587_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6588_));
OR2X2 OR2X2_1846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6590_), .B(AES_CORE_DATAPATH__abc_16009_new_n6591_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6592_));
OR2X2 OR2X2_1847 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6593_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6594_));
OR2X2 OR2X2_1848 ( .A(\iv_out[16] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6595_));
OR2X2 OR2X2_1849 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6593_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6598_));
OR2X2 OR2X2_185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2736_));
OR2X2 OR2X2_1850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6599_));
OR2X2 OR2X2_1851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6601_), .B(AES_CORE_DATAPATH__abc_16009_new_n6602_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6603_));
OR2X2 OR2X2_1852 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6603_), .B(AES_CORE_DATAPATH__abc_16009_new_n6597_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6604_));
OR2X2 OR2X2_1853 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6605_), .B(AES_CORE_DATAPATH__abc_16009_new_n6606_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6607_));
OR2X2 OR2X2_1854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6607_), .B(AES_CORE_DATAPATH__abc_16009_new_n6565_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6608_));
OR2X2 OR2X2_1855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6609_), .B(AES_CORE_DATAPATH__abc_16009_new_n6561_), .Y(AES_CORE_DATAPATH__0col_0__31_0__16_));
OR2X2 OR2X2_1856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6612_), .B(AES_CORE_DATAPATH__abc_16009_new_n6613_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6614_));
OR2X2 OR2X2_1857 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6618_), .B(AES_CORE_DATAPATH__abc_16009_new_n6619_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6620_));
OR2X2 OR2X2_1858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6622_));
OR2X2 OR2X2_1859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6621_), .B(AES_CORE_DATAPATH__abc_16009_new_n6623_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6624_));
OR2X2 OR2X2_186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2738_), .B(AES_CORE_DATAPATH__abc_16009_new_n2739_), .Y(\iv_out[25] ));
OR2X2 OR2X2_1860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6627_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6628_));
OR2X2 OR2X2_1861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6628_), .B(AES_CORE_DATAPATH__abc_16009_new_n6626_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6629_));
OR2X2 OR2X2_1862 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6630_));
OR2X2 OR2X2_1863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6632_), .B(AES_CORE_DATAPATH__abc_16009_new_n6633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6634_));
OR2X2 OR2X2_1864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6634_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6635_));
OR2X2 OR2X2_1865 ( .A(\iv_out[17] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6636_));
OR2X2 OR2X2_1866 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6624_), .B(AES_CORE_DATAPATH__abc_16009_new_n6638_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6639_));
OR2X2 OR2X2_1867 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4008_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6640_));
OR2X2 OR2X2_1868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6641_), .B(AES_CORE_DATAPATH__abc_16009_new_n6637_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6642_));
OR2X2 OR2X2_1869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6643_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6644_));
OR2X2 OR2X2_187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2743_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2744_));
OR2X2 OR2X2_1870 ( .A(\iv_out[17] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6645_));
OR2X2 OR2X2_1871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6643_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6648_));
OR2X2 OR2X2_1872 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6649_));
OR2X2 OR2X2_1873 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6651_), .B(AES_CORE_DATAPATH__abc_16009_new_n6652_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6653_));
OR2X2 OR2X2_1874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6653_), .B(AES_CORE_DATAPATH__abc_16009_new_n6647_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6654_));
OR2X2 OR2X2_1875 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6655_), .B(AES_CORE_DATAPATH__abc_16009_new_n6656_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6657_));
OR2X2 OR2X2_1876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6657_), .B(AES_CORE_DATAPATH__abc_16009_new_n6615_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6658_));
OR2X2 OR2X2_1877 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6659_), .B(AES_CORE_DATAPATH__abc_16009_new_n6611_), .Y(AES_CORE_DATAPATH__0col_0__31_0__17_));
OR2X2 OR2X2_1878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6662_), .B(AES_CORE_DATAPATH__abc_16009_new_n6663_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6664_));
OR2X2 OR2X2_1879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6668_), .B(AES_CORE_DATAPATH__abc_16009_new_n6669_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6670_));
OR2X2 OR2X2_188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2744_), .B(AES_CORE_DATAPATH__abc_16009_new_n2742_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2745_));
OR2X2 OR2X2_1880 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6672_));
OR2X2 OR2X2_1881 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6671_), .B(AES_CORE_DATAPATH__abc_16009_new_n6673_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6674_));
OR2X2 OR2X2_1882 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6677_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6678_));
OR2X2 OR2X2_1883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6678_), .B(AES_CORE_DATAPATH__abc_16009_new_n6676_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6679_));
OR2X2 OR2X2_1884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6680_));
OR2X2 OR2X2_1885 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6682_), .B(AES_CORE_DATAPATH__abc_16009_new_n6683_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6684_));
OR2X2 OR2X2_1886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6684_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6685_));
OR2X2 OR2X2_1887 ( .A(\iv_out[18] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6686_));
OR2X2 OR2X2_1888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6674_), .B(AES_CORE_DATAPATH__abc_16009_new_n6688_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6689_));
OR2X2 OR2X2_1889 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4040_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6690_));
OR2X2 OR2X2_189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2746_));
OR2X2 OR2X2_1890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6691_), .B(AES_CORE_DATAPATH__abc_16009_new_n6687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6692_));
OR2X2 OR2X2_1891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6693_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6694_));
OR2X2 OR2X2_1892 ( .A(\iv_out[18] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6695_));
OR2X2 OR2X2_1893 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6693_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6698_));
OR2X2 OR2X2_1894 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6699_));
OR2X2 OR2X2_1895 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6701_), .B(AES_CORE_DATAPATH__abc_16009_new_n6702_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6703_));
OR2X2 OR2X2_1896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6703_), .B(AES_CORE_DATAPATH__abc_16009_new_n6697_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6704_));
OR2X2 OR2X2_1897 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6705_), .B(AES_CORE_DATAPATH__abc_16009_new_n6706_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6707_));
OR2X2 OR2X2_1898 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6707_), .B(AES_CORE_DATAPATH__abc_16009_new_n6665_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6708_));
OR2X2 OR2X2_1899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6709_), .B(AES_CORE_DATAPATH__abc_16009_new_n6661_), .Y(AES_CORE_DATAPATH__0col_0__31_0__18_));
OR2X2 OR2X2_19 ( .A(AES_CORE_CONTROL_UNIT_state_8_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_));
OR2X2 OR2X2_190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2748_), .B(AES_CORE_DATAPATH__abc_16009_new_n2749_), .Y(\iv_out[26] ));
OR2X2 OR2X2_1900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6712_), .B(AES_CORE_DATAPATH__abc_16009_new_n6713_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6714_));
OR2X2 OR2X2_1901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6718_), .B(AES_CORE_DATAPATH__abc_16009_new_n6719_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6720_));
OR2X2 OR2X2_1902 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6722_));
OR2X2 OR2X2_1903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6721_), .B(AES_CORE_DATAPATH__abc_16009_new_n6723_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6724_));
OR2X2 OR2X2_1904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6727_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6728_));
OR2X2 OR2X2_1905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6728_), .B(AES_CORE_DATAPATH__abc_16009_new_n6726_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6729_));
OR2X2 OR2X2_1906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6730_));
OR2X2 OR2X2_1907 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6732_), .B(AES_CORE_DATAPATH__abc_16009_new_n6733_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6734_));
OR2X2 OR2X2_1908 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6734_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6735_));
OR2X2 OR2X2_1909 ( .A(\iv_out[19] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6736_));
OR2X2 OR2X2_191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2753_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2754_));
OR2X2 OR2X2_1910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6724_), .B(AES_CORE_DATAPATH__abc_16009_new_n6738_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6739_));
OR2X2 OR2X2_1911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4072_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6740_));
OR2X2 OR2X2_1912 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6741_), .B(AES_CORE_DATAPATH__abc_16009_new_n6737_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6742_));
OR2X2 OR2X2_1913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6743_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6744_));
OR2X2 OR2X2_1914 ( .A(\iv_out[19] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6745_));
OR2X2 OR2X2_1915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6743_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6748_));
OR2X2 OR2X2_1916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6749_));
OR2X2 OR2X2_1917 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6751_), .B(AES_CORE_DATAPATH__abc_16009_new_n6752_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6753_));
OR2X2 OR2X2_1918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6753_), .B(AES_CORE_DATAPATH__abc_16009_new_n6747_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6754_));
OR2X2 OR2X2_1919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6755_), .B(AES_CORE_DATAPATH__abc_16009_new_n6756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6757_));
OR2X2 OR2X2_192 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2754_), .B(AES_CORE_DATAPATH__abc_16009_new_n2752_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2755_));
OR2X2 OR2X2_1920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6757_), .B(AES_CORE_DATAPATH__abc_16009_new_n6715_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6758_));
OR2X2 OR2X2_1921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6759_), .B(AES_CORE_DATAPATH__abc_16009_new_n6711_), .Y(AES_CORE_DATAPATH__0col_0__31_0__19_));
OR2X2 OR2X2_1922 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6762_), .B(AES_CORE_DATAPATH__abc_16009_new_n6763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6764_));
OR2X2 OR2X2_1923 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6766_), .B(AES_CORE_DATAPATH__abc_16009_new_n6767_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6768_));
OR2X2 OR2X2_1924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6771_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6772_));
OR2X2 OR2X2_1925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6772_), .B(AES_CORE_DATAPATH__abc_16009_new_n6770_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6773_));
OR2X2 OR2X2_1926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6774_));
OR2X2 OR2X2_1927 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6776_), .B(AES_CORE_DATAPATH__abc_16009_new_n6777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6778_));
OR2X2 OR2X2_1928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6778_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6779_));
OR2X2 OR2X2_1929 ( .A(\iv_out[20] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6780_));
OR2X2 OR2X2_193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2756_));
OR2X2 OR2X2_1930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6768_), .B(AES_CORE_DATAPATH__abc_16009_new_n6781_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6782_));
OR2X2 OR2X2_1931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6785_), .B(AES_CORE_DATAPATH__abc_16009_new_n6786_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6787_));
OR2X2 OR2X2_1932 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6787_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6788_));
OR2X2 OR2X2_1933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6790_), .B(AES_CORE_DATAPATH__abc_16009_new_n6791_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6792_));
OR2X2 OR2X2_1934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6793_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6794_));
OR2X2 OR2X2_1935 ( .A(\iv_out[20] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6795_));
OR2X2 OR2X2_1936 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6793_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6798_));
OR2X2 OR2X2_1937 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6799_));
OR2X2 OR2X2_1938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6801_), .B(AES_CORE_DATAPATH__abc_16009_new_n6802_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6803_));
OR2X2 OR2X2_1939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6803_), .B(AES_CORE_DATAPATH__abc_16009_new_n6797_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6804_));
OR2X2 OR2X2_194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2758_), .B(AES_CORE_DATAPATH__abc_16009_new_n2759_), .Y(\iv_out[27] ));
OR2X2 OR2X2_1940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6805_), .B(AES_CORE_DATAPATH__abc_16009_new_n6806_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6807_));
OR2X2 OR2X2_1941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6807_), .B(AES_CORE_DATAPATH__abc_16009_new_n6765_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6808_));
OR2X2 OR2X2_1942 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6809_), .B(AES_CORE_DATAPATH__abc_16009_new_n6761_), .Y(AES_CORE_DATAPATH__0col_0__31_0__20_));
OR2X2 OR2X2_1943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6812_), .B(AES_CORE_DATAPATH__abc_16009_new_n6813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6814_));
OR2X2 OR2X2_1944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6818_), .B(AES_CORE_DATAPATH__abc_16009_new_n6819_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6820_));
OR2X2 OR2X2_1945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6822_));
OR2X2 OR2X2_1946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6821_), .B(AES_CORE_DATAPATH__abc_16009_new_n6823_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6824_));
OR2X2 OR2X2_1947 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6827_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6828_));
OR2X2 OR2X2_1948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6828_), .B(AES_CORE_DATAPATH__abc_16009_new_n6826_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6829_));
OR2X2 OR2X2_1949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6830_));
OR2X2 OR2X2_195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2763_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2764_));
OR2X2 OR2X2_1950 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6832_), .B(AES_CORE_DATAPATH__abc_16009_new_n6833_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6834_));
OR2X2 OR2X2_1951 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6834_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6835_));
OR2X2 OR2X2_1952 ( .A(\iv_out[21] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6836_));
OR2X2 OR2X2_1953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6824_), .B(AES_CORE_DATAPATH__abc_16009_new_n6838_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6839_));
OR2X2 OR2X2_1954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4136_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6840_));
OR2X2 OR2X2_1955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6841_), .B(AES_CORE_DATAPATH__abc_16009_new_n6837_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6842_));
OR2X2 OR2X2_1956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6843_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6844_));
OR2X2 OR2X2_1957 ( .A(\iv_out[21] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6845_));
OR2X2 OR2X2_1958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6843_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6848_));
OR2X2 OR2X2_1959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6849_));
OR2X2 OR2X2_196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2764_), .B(AES_CORE_DATAPATH__abc_16009_new_n2762_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2765_));
OR2X2 OR2X2_1960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6851_), .B(AES_CORE_DATAPATH__abc_16009_new_n6852_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6853_));
OR2X2 OR2X2_1961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6853_), .B(AES_CORE_DATAPATH__abc_16009_new_n6847_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6854_));
OR2X2 OR2X2_1962 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6855_), .B(AES_CORE_DATAPATH__abc_16009_new_n6856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6857_));
OR2X2 OR2X2_1963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6857_), .B(AES_CORE_DATAPATH__abc_16009_new_n6815_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6858_));
OR2X2 OR2X2_1964 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6859_), .B(AES_CORE_DATAPATH__abc_16009_new_n6811_), .Y(AES_CORE_DATAPATH__0col_0__31_0__21_));
OR2X2 OR2X2_1965 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6862_), .B(AES_CORE_DATAPATH__abc_16009_new_n6863_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6864_));
OR2X2 OR2X2_1966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6866_), .B(AES_CORE_DATAPATH__abc_16009_new_n6867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6868_));
OR2X2 OR2X2_1967 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6871_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6872_));
OR2X2 OR2X2_1968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6872_), .B(AES_CORE_DATAPATH__abc_16009_new_n6870_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6873_));
OR2X2 OR2X2_1969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6874_));
OR2X2 OR2X2_197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2766_));
OR2X2 OR2X2_1970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6876_), .B(AES_CORE_DATAPATH__abc_16009_new_n6877_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6878_));
OR2X2 OR2X2_1971 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6878_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6879_));
OR2X2 OR2X2_1972 ( .A(\iv_out[22] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6880_));
OR2X2 OR2X2_1973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6868_), .B(AES_CORE_DATAPATH__abc_16009_new_n6881_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6882_));
OR2X2 OR2X2_1974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6885_), .B(AES_CORE_DATAPATH__abc_16009_new_n6886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6887_));
OR2X2 OR2X2_1975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6887_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6888_));
OR2X2 OR2X2_1976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6890_), .B(AES_CORE_DATAPATH__abc_16009_new_n6891_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6892_));
OR2X2 OR2X2_1977 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6893_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6894_));
OR2X2 OR2X2_1978 ( .A(\iv_out[22] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6895_));
OR2X2 OR2X2_1979 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6893_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6898_));
OR2X2 OR2X2_198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2768_), .B(AES_CORE_DATAPATH__abc_16009_new_n2769_), .Y(\iv_out[28] ));
OR2X2 OR2X2_1980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6899_));
OR2X2 OR2X2_1981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6901_), .B(AES_CORE_DATAPATH__abc_16009_new_n6902_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6903_));
OR2X2 OR2X2_1982 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6903_), .B(AES_CORE_DATAPATH__abc_16009_new_n6897_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6904_));
OR2X2 OR2X2_1983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6905_), .B(AES_CORE_DATAPATH__abc_16009_new_n6906_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6907_));
OR2X2 OR2X2_1984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6907_), .B(AES_CORE_DATAPATH__abc_16009_new_n6865_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6908_));
OR2X2 OR2X2_1985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6909_), .B(AES_CORE_DATAPATH__abc_16009_new_n6861_), .Y(AES_CORE_DATAPATH__0col_0__31_0__22_));
OR2X2 OR2X2_1986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6912_), .B(AES_CORE_DATAPATH__abc_16009_new_n6913_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6914_));
OR2X2 OR2X2_1987 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6918_), .B(AES_CORE_DATAPATH__abc_16009_new_n6919_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6920_));
OR2X2 OR2X2_1988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6922_));
OR2X2 OR2X2_1989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6921_), .B(AES_CORE_DATAPATH__abc_16009_new_n6923_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6924_));
OR2X2 OR2X2_199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2773_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2774_));
OR2X2 OR2X2_1990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6927_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6928_));
OR2X2 OR2X2_1991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6928_), .B(AES_CORE_DATAPATH__abc_16009_new_n6926_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6929_));
OR2X2 OR2X2_1992 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6930_));
OR2X2 OR2X2_1993 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6932_), .B(AES_CORE_DATAPATH__abc_16009_new_n6933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6934_));
OR2X2 OR2X2_1994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6934_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6935_));
OR2X2 OR2X2_1995 ( .A(\iv_out[23] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6936_));
OR2X2 OR2X2_1996 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6924_), .B(AES_CORE_DATAPATH__abc_16009_new_n6938_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6939_));
OR2X2 OR2X2_1997 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4200_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6940_));
OR2X2 OR2X2_1998 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6941_), .B(AES_CORE_DATAPATH__abc_16009_new_n6937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6942_));
OR2X2 OR2X2_1999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6943_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6944_));
OR2X2 OR2X2_2 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n95_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n96_));
OR2X2 OR2X2_20 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n144_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n146_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n147_));
OR2X2 OR2X2_200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2774_), .B(AES_CORE_DATAPATH__abc_16009_new_n2772_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2775_));
OR2X2 OR2X2_2000 ( .A(\iv_out[23] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6945_));
OR2X2 OR2X2_2001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6943_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6948_));
OR2X2 OR2X2_2002 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6949_));
OR2X2 OR2X2_2003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6951_), .B(AES_CORE_DATAPATH__abc_16009_new_n6952_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6953_));
OR2X2 OR2X2_2004 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6953_), .B(AES_CORE_DATAPATH__abc_16009_new_n6947_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6954_));
OR2X2 OR2X2_2005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6955_), .B(AES_CORE_DATAPATH__abc_16009_new_n6956_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6957_));
OR2X2 OR2X2_2006 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6957_), .B(AES_CORE_DATAPATH__abc_16009_new_n6915_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6958_));
OR2X2 OR2X2_2007 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6959_), .B(AES_CORE_DATAPATH__abc_16009_new_n6911_), .Y(AES_CORE_DATAPATH__0col_0__31_0__23_));
OR2X2 OR2X2_2008 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6962_), .B(AES_CORE_DATAPATH__abc_16009_new_n6963_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6964_));
OR2X2 OR2X2_2009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6966_), .B(AES_CORE_DATAPATH__abc_16009_new_n6967_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6968_));
OR2X2 OR2X2_201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2776_));
OR2X2 OR2X2_2010 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6971_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6972_));
OR2X2 OR2X2_2011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6972_), .B(AES_CORE_DATAPATH__abc_16009_new_n6970_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6973_));
OR2X2 OR2X2_2012 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6974_));
OR2X2 OR2X2_2013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6976_), .B(AES_CORE_DATAPATH__abc_16009_new_n6977_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6978_));
OR2X2 OR2X2_2014 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6978_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6979_));
OR2X2 OR2X2_2015 ( .A(\iv_out[24] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6980_));
OR2X2 OR2X2_2016 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6968_), .B(AES_CORE_DATAPATH__abc_16009_new_n6981_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6982_));
OR2X2 OR2X2_2017 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6985_), .B(AES_CORE_DATAPATH__abc_16009_new_n6986_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6987_));
OR2X2 OR2X2_2018 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6987_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6988_));
OR2X2 OR2X2_2019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6990_), .B(AES_CORE_DATAPATH__abc_16009_new_n6991_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6992_));
OR2X2 OR2X2_202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2778_), .B(AES_CORE_DATAPATH__abc_16009_new_n2779_), .Y(\iv_out[29] ));
OR2X2 OR2X2_2020 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6993_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6994_));
OR2X2 OR2X2_2021 ( .A(\iv_out[24] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n6995_));
OR2X2 OR2X2_2022 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6993_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6998_));
OR2X2 OR2X2_2023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n6999_));
OR2X2 OR2X2_2024 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7001_), .B(AES_CORE_DATAPATH__abc_16009_new_n7002_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7003_));
OR2X2 OR2X2_2025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7003_), .B(AES_CORE_DATAPATH__abc_16009_new_n6997_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7004_));
OR2X2 OR2X2_2026 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7005_), .B(AES_CORE_DATAPATH__abc_16009_new_n7006_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7007_));
OR2X2 OR2X2_2027 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7007_), .B(AES_CORE_DATAPATH__abc_16009_new_n6965_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7008_));
OR2X2 OR2X2_2028 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7009_), .B(AES_CORE_DATAPATH__abc_16009_new_n6961_), .Y(AES_CORE_DATAPATH__0col_0__31_0__24_));
OR2X2 OR2X2_2029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7012_), .B(AES_CORE_DATAPATH__abc_16009_new_n7013_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7014_));
OR2X2 OR2X2_203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2783_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2784_));
OR2X2 OR2X2_2030 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7018_), .B(AES_CORE_DATAPATH__abc_16009_new_n7019_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7020_));
OR2X2 OR2X2_2031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7022_));
OR2X2 OR2X2_2032 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7021_), .B(AES_CORE_DATAPATH__abc_16009_new_n7023_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7024_));
OR2X2 OR2X2_2033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7027_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7028_));
OR2X2 OR2X2_2034 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7028_), .B(AES_CORE_DATAPATH__abc_16009_new_n7026_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7029_));
OR2X2 OR2X2_2035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7030_));
OR2X2 OR2X2_2036 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7032_), .B(AES_CORE_DATAPATH__abc_16009_new_n7033_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7034_));
OR2X2 OR2X2_2037 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7034_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7035_));
OR2X2 OR2X2_2038 ( .A(\iv_out[25] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7036_));
OR2X2 OR2X2_2039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7024_), .B(AES_CORE_DATAPATH__abc_16009_new_n7038_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7039_));
OR2X2 OR2X2_204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2784_), .B(AES_CORE_DATAPATH__abc_16009_new_n2782_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2785_));
OR2X2 OR2X2_2040 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4264_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7040_));
OR2X2 OR2X2_2041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7041_), .B(AES_CORE_DATAPATH__abc_16009_new_n7037_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7042_));
OR2X2 OR2X2_2042 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7043_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7044_));
OR2X2 OR2X2_2043 ( .A(\iv_out[25] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7045_));
OR2X2 OR2X2_2044 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7043_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7048_));
OR2X2 OR2X2_2045 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7049_));
OR2X2 OR2X2_2046 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7051_), .B(AES_CORE_DATAPATH__abc_16009_new_n7052_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7053_));
OR2X2 OR2X2_2047 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7053_), .B(AES_CORE_DATAPATH__abc_16009_new_n7047_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7054_));
OR2X2 OR2X2_2048 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7055_), .B(AES_CORE_DATAPATH__abc_16009_new_n7056_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7057_));
OR2X2 OR2X2_2049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7057_), .B(AES_CORE_DATAPATH__abc_16009_new_n7015_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7058_));
OR2X2 OR2X2_205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2786_));
OR2X2 OR2X2_2050 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7059_), .B(AES_CORE_DATAPATH__abc_16009_new_n7011_), .Y(AES_CORE_DATAPATH__0col_0__31_0__25_));
OR2X2 OR2X2_2051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7062_), .B(AES_CORE_DATAPATH__abc_16009_new_n7063_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7064_));
OR2X2 OR2X2_2052 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7068_), .B(AES_CORE_DATAPATH__abc_16009_new_n7069_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7070_));
OR2X2 OR2X2_2053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7072_));
OR2X2 OR2X2_2054 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7071_), .B(AES_CORE_DATAPATH__abc_16009_new_n7073_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7074_));
OR2X2 OR2X2_2055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7077_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7078_));
OR2X2 OR2X2_2056 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7078_), .B(AES_CORE_DATAPATH__abc_16009_new_n7076_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7079_));
OR2X2 OR2X2_2057 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7080_));
OR2X2 OR2X2_2058 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7082_), .B(AES_CORE_DATAPATH__abc_16009_new_n7083_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7084_));
OR2X2 OR2X2_2059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7084_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7085_));
OR2X2 OR2X2_206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2788_), .B(AES_CORE_DATAPATH__abc_16009_new_n2789_), .Y(\iv_out[30] ));
OR2X2 OR2X2_2060 ( .A(\iv_out[26] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7086_));
OR2X2 OR2X2_2061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7074_), .B(AES_CORE_DATAPATH__abc_16009_new_n7088_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7089_));
OR2X2 OR2X2_2062 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4296_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7090_));
OR2X2 OR2X2_2063 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7091_), .B(AES_CORE_DATAPATH__abc_16009_new_n7087_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7092_));
OR2X2 OR2X2_2064 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7093_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7094_));
OR2X2 OR2X2_2065 ( .A(\iv_out[26] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7095_));
OR2X2 OR2X2_2066 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7093_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7098_));
OR2X2 OR2X2_2067 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7099_));
OR2X2 OR2X2_2068 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7101_), .B(AES_CORE_DATAPATH__abc_16009_new_n7102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7103_));
OR2X2 OR2X2_2069 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7103_), .B(AES_CORE_DATAPATH__abc_16009_new_n7097_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7104_));
OR2X2 OR2X2_207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2793_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2794_));
OR2X2 OR2X2_2070 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7105_), .B(AES_CORE_DATAPATH__abc_16009_new_n7106_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7107_));
OR2X2 OR2X2_2071 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7107_), .B(AES_CORE_DATAPATH__abc_16009_new_n7065_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7108_));
OR2X2 OR2X2_2072 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7109_), .B(AES_CORE_DATAPATH__abc_16009_new_n7061_), .Y(AES_CORE_DATAPATH__0col_0__31_0__26_));
OR2X2 OR2X2_2073 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7112_), .B(AES_CORE_DATAPATH__abc_16009_new_n7113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7114_));
OR2X2 OR2X2_2074 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7116_), .B(AES_CORE_DATAPATH__abc_16009_new_n7117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7118_));
OR2X2 OR2X2_2075 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7121_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7122_));
OR2X2 OR2X2_2076 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7122_), .B(AES_CORE_DATAPATH__abc_16009_new_n7120_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7123_));
OR2X2 OR2X2_2077 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7124_));
OR2X2 OR2X2_2078 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7126_), .B(AES_CORE_DATAPATH__abc_16009_new_n7127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7128_));
OR2X2 OR2X2_2079 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7128_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7129_));
OR2X2 OR2X2_208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2794_), .B(AES_CORE_DATAPATH__abc_16009_new_n2792_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2795_));
OR2X2 OR2X2_2080 ( .A(\iv_out[27] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7130_));
OR2X2 OR2X2_2081 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7118_), .B(AES_CORE_DATAPATH__abc_16009_new_n7131_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7132_));
OR2X2 OR2X2_2082 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7135_), .B(AES_CORE_DATAPATH__abc_16009_new_n7136_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7137_));
OR2X2 OR2X2_2083 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7137_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7138_));
OR2X2 OR2X2_2084 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7140_), .B(AES_CORE_DATAPATH__abc_16009_new_n7141_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7142_));
OR2X2 OR2X2_2085 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7143_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7144_));
OR2X2 OR2X2_2086 ( .A(\iv_out[27] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7145_));
OR2X2 OR2X2_2087 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7143_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7148_));
OR2X2 OR2X2_2088 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7149_));
OR2X2 OR2X2_2089 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7151_), .B(AES_CORE_DATAPATH__abc_16009_new_n7152_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7153_));
OR2X2 OR2X2_209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2796_));
OR2X2 OR2X2_2090 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7153_), .B(AES_CORE_DATAPATH__abc_16009_new_n7147_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7154_));
OR2X2 OR2X2_2091 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7155_), .B(AES_CORE_DATAPATH__abc_16009_new_n7156_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7157_));
OR2X2 OR2X2_2092 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7157_), .B(AES_CORE_DATAPATH__abc_16009_new_n7115_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7158_));
OR2X2 OR2X2_2093 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7159_), .B(AES_CORE_DATAPATH__abc_16009_new_n7111_), .Y(AES_CORE_DATAPATH__0col_0__31_0__27_));
OR2X2 OR2X2_2094 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7162_), .B(AES_CORE_DATAPATH__abc_16009_new_n7163_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7164_));
OR2X2 OR2X2_2095 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7168_), .B(AES_CORE_DATAPATH__abc_16009_new_n7169_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7170_));
OR2X2 OR2X2_2096 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7172_));
OR2X2 OR2X2_2097 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7171_), .B(AES_CORE_DATAPATH__abc_16009_new_n7173_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7174_));
OR2X2 OR2X2_2098 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7177_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7178_));
OR2X2 OR2X2_2099 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7178_), .B(AES_CORE_DATAPATH__abc_16009_new_n7176_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7179_));
OR2X2 OR2X2_21 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n149_), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_));
OR2X2 OR2X2_210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2798_), .B(AES_CORE_DATAPATH__abc_16009_new_n2799_), .Y(\iv_out[31] ));
OR2X2 OR2X2_2100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7180_));
OR2X2 OR2X2_2101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7182_), .B(AES_CORE_DATAPATH__abc_16009_new_n7183_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7184_));
OR2X2 OR2X2_2102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7184_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7185_));
OR2X2 OR2X2_2103 ( .A(\iv_out[28] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7186_));
OR2X2 OR2X2_2104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7174_), .B(AES_CORE_DATAPATH__abc_16009_new_n7188_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7189_));
OR2X2 OR2X2_2105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4360_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7190_));
OR2X2 OR2X2_2106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7191_), .B(AES_CORE_DATAPATH__abc_16009_new_n7187_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7192_));
OR2X2 OR2X2_2107 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7193_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7194_));
OR2X2 OR2X2_2108 ( .A(\iv_out[28] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7195_));
OR2X2 OR2X2_2109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7193_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7198_));
OR2X2 OR2X2_211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2804_));
OR2X2 OR2X2_2110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7199_));
OR2X2 OR2X2_2111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7201_), .B(AES_CORE_DATAPATH__abc_16009_new_n7202_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7203_));
OR2X2 OR2X2_2112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7203_), .B(AES_CORE_DATAPATH__abc_16009_new_n7197_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7204_));
OR2X2 OR2X2_2113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7205_), .B(AES_CORE_DATAPATH__abc_16009_new_n7206_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7207_));
OR2X2 OR2X2_2114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7207_), .B(AES_CORE_DATAPATH__abc_16009_new_n7165_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7208_));
OR2X2 OR2X2_2115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7209_), .B(AES_CORE_DATAPATH__abc_16009_new_n7161_), .Y(AES_CORE_DATAPATH__0col_0__31_0__28_));
OR2X2 OR2X2_2116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7212_), .B(AES_CORE_DATAPATH__abc_16009_new_n7213_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7214_));
OR2X2 OR2X2_2117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7216_), .B(AES_CORE_DATAPATH__abc_16009_new_n7217_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7218_));
OR2X2 OR2X2_2118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7221_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7222_));
OR2X2 OR2X2_2119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7222_), .B(AES_CORE_DATAPATH__abc_16009_new_n7220_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7223_));
OR2X2 OR2X2_212 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_mode_ctr), .Y(AES_CORE_DATAPATH__abc_16009_new_n2805_));
OR2X2 OR2X2_2120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7224_));
OR2X2 OR2X2_2121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7226_), .B(AES_CORE_DATAPATH__abc_16009_new_n7227_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7228_));
OR2X2 OR2X2_2122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7228_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7229_));
OR2X2 OR2X2_2123 ( .A(\iv_out[29] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7230_));
OR2X2 OR2X2_2124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7218_), .B(AES_CORE_DATAPATH__abc_16009_new_n7231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7232_));
OR2X2 OR2X2_2125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7235_), .B(AES_CORE_DATAPATH__abc_16009_new_n7236_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7237_));
OR2X2 OR2X2_2126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7237_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7238_));
OR2X2 OR2X2_2127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7240_), .B(AES_CORE_DATAPATH__abc_16009_new_n7241_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7242_));
OR2X2 OR2X2_2128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7243_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7244_));
OR2X2 OR2X2_2129 ( .A(\iv_out[29] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7245_));
OR2X2 OR2X2_213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2808_), .B(AES_CORE_DATAPATH__abc_16009_new_n2809_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2810_));
OR2X2 OR2X2_2130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7243_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7248_));
OR2X2 OR2X2_2131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7249_));
OR2X2 OR2X2_2132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7251_), .B(AES_CORE_DATAPATH__abc_16009_new_n7252_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7253_));
OR2X2 OR2X2_2133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7253_), .B(AES_CORE_DATAPATH__abc_16009_new_n7247_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7254_));
OR2X2 OR2X2_2134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7255_), .B(AES_CORE_DATAPATH__abc_16009_new_n7256_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7257_));
OR2X2 OR2X2_2135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7257_), .B(AES_CORE_DATAPATH__abc_16009_new_n7215_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7258_));
OR2X2 OR2X2_2136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7259_), .B(AES_CORE_DATAPATH__abc_16009_new_n7211_), .Y(AES_CORE_DATAPATH__0col_0__31_0__29_));
OR2X2 OR2X2_2137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7262_), .B(AES_CORE_DATAPATH__abc_16009_new_n7263_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7264_));
OR2X2 OR2X2_2138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7266_), .B(AES_CORE_DATAPATH__abc_16009_new_n7267_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7268_));
OR2X2 OR2X2_2139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7271_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7272_));
OR2X2 OR2X2_214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2812_), .B(\key_sel_rd[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2813_));
OR2X2 OR2X2_2140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7272_), .B(AES_CORE_DATAPATH__abc_16009_new_n7270_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7273_));
OR2X2 OR2X2_2141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7274_));
OR2X2 OR2X2_2142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7276_), .B(AES_CORE_DATAPATH__abc_16009_new_n7277_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7278_));
OR2X2 OR2X2_2143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7278_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7279_));
OR2X2 OR2X2_2144 ( .A(\iv_out[30] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7280_));
OR2X2 OR2X2_2145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7268_), .B(AES_CORE_DATAPATH__abc_16009_new_n7281_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7282_));
OR2X2 OR2X2_2146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7285_), .B(AES_CORE_DATAPATH__abc_16009_new_n7286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7287_));
OR2X2 OR2X2_2147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7287_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7288_));
OR2X2 OR2X2_2148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7290_), .B(AES_CORE_DATAPATH__abc_16009_new_n7291_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7292_));
OR2X2 OR2X2_2149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7293_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7294_));
OR2X2 OR2X2_215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2811_), .B(AES_CORE_DATAPATH__abc_16009_new_n2813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2814_));
OR2X2 OR2X2_2150 ( .A(\iv_out[30] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7295_));
OR2X2 OR2X2_2151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7293_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7298_));
OR2X2 OR2X2_2152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7299_));
OR2X2 OR2X2_2153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7301_), .B(AES_CORE_DATAPATH__abc_16009_new_n7302_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7303_));
OR2X2 OR2X2_2154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7303_), .B(AES_CORE_DATAPATH__abc_16009_new_n7297_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7304_));
OR2X2 OR2X2_2155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7305_), .B(AES_CORE_DATAPATH__abc_16009_new_n7306_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7307_));
OR2X2 OR2X2_2156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7307_), .B(AES_CORE_DATAPATH__abc_16009_new_n7265_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7308_));
OR2X2 OR2X2_2157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7309_), .B(AES_CORE_DATAPATH__abc_16009_new_n7261_), .Y(AES_CORE_DATAPATH__0col_0__31_0__30_));
OR2X2 OR2X2_2158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7312_), .B(AES_CORE_DATAPATH__abc_16009_new_n7313_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7314_));
OR2X2 OR2X2_2159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7318_), .B(AES_CORE_DATAPATH__abc_16009_new_n7319_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7320_));
OR2X2 OR2X2_216 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2815_), .B(AES_CORE_DATAPATH__abc_16009_new_n2816_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2817_));
OR2X2 OR2X2_2160 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5759_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7322_));
OR2X2 OR2X2_2161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7321_), .B(AES_CORE_DATAPATH__abc_16009_new_n7323_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7324_));
OR2X2 OR2X2_2162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7327_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7328_));
OR2X2 OR2X2_2163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7328_), .B(AES_CORE_DATAPATH__abc_16009_new_n7326_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7329_));
OR2X2 OR2X2_2164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_bkp_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7330_));
OR2X2 OR2X2_2165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7332_), .B(AES_CORE_DATAPATH__abc_16009_new_n7333_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7334_));
OR2X2 OR2X2_2166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7334_), .B(AES_CORE_DATAPATH__abc_16009_new_n5763_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7335_));
OR2X2 OR2X2_2167 ( .A(\iv_out[31] ), .B(AES_CORE_DATAPATH__abc_16009_new_n5764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7336_));
OR2X2 OR2X2_2168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7324_), .B(AES_CORE_DATAPATH__abc_16009_new_n7338_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7339_));
OR2X2 OR2X2_2169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4456_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7340_));
OR2X2 OR2X2_217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2819_), .B(\key_sel_rd[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2820_));
OR2X2 OR2X2_2170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7341_), .B(AES_CORE_DATAPATH__abc_16009_new_n7337_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7342_));
OR2X2 OR2X2_2171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7343_), .B(AES_CORE_DATAPATH__abc_16009_new_n5757_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7344_));
OR2X2 OR2X2_2172 ( .A(\iv_out[31] ), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_DATAPATH__abc_16009_new_n7345_));
OR2X2 OR2X2_2173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7343_), .B(AES_CORE_DATAPATH__abc_16009_new_n5796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7348_));
OR2X2 OR2X2_2174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5798_), .B(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7349_));
OR2X2 OR2X2_2175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7351_), .B(AES_CORE_DATAPATH__abc_16009_new_n7352_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7353_));
OR2X2 OR2X2_2176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7353_), .B(AES_CORE_DATAPATH__abc_16009_new_n7347_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7354_));
OR2X2 OR2X2_2177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7355_), .B(AES_CORE_DATAPATH__abc_16009_new_n7356_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7357_));
OR2X2 OR2X2_2178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7357_), .B(AES_CORE_DATAPATH__abc_16009_new_n7315_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7358_));
OR2X2 OR2X2_2179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7359_), .B(AES_CORE_DATAPATH__abc_16009_new_n7311_), .Y(AES_CORE_DATAPATH__0col_0__31_0__31_));
OR2X2 OR2X2_218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2818_), .B(AES_CORE_DATAPATH__abc_16009_new_n2820_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2821_));
OR2X2 OR2X2_2180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7361_), .B(AES_CORE_DATAPATH__abc_16009_new_n7362_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7363_));
OR2X2 OR2X2_2181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7369_), .B(AES_CORE_DATAPATH__abc_16009_new_n7368_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7370_));
OR2X2 OR2X2_2182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7370_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7371_));
OR2X2 OR2X2_2183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7372_));
OR2X2 OR2X2_2184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7373_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7374_));
OR2X2 OR2X2_2185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7376_));
OR2X2 OR2X2_2186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7378_));
OR2X2 OR2X2_2187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7379_), .B(AES_CORE_DATAPATH__abc_16009_new_n7380_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7381_));
OR2X2 OR2X2_2188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7381_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7382_));
OR2X2 OR2X2_2189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7383_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7384_));
OR2X2 OR2X2_219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2814_), .B(AES_CORE_DATAPATH__abc_16009_new_n2821_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2822_));
OR2X2 OR2X2_2190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7385_));
OR2X2 OR2X2_2191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7387_));
OR2X2 OR2X2_2192 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7388_), .B(AES_CORE_DATAPATH__abc_16009_new_n7389_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7390_));
OR2X2 OR2X2_2193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7390_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7391_));
OR2X2 OR2X2_2194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7392_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7393_));
OR2X2 OR2X2_2195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7394_));
OR2X2 OR2X2_2196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7396_));
OR2X2 OR2X2_2197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7397_), .B(AES_CORE_DATAPATH__abc_16009_new_n7398_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7399_));
OR2X2 OR2X2_2198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7399_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7400_));
OR2X2 OR2X2_2199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7401_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7402_));
OR2X2 OR2X2_22 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_), .Y(AES_CORE_CONTROL_UNIT_bypass_key_en));
OR2X2 OR2X2_220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2823_));
OR2X2 OR2X2_2200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7403_));
OR2X2 OR2X2_2201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7405_));
OR2X2 OR2X2_2202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7406_), .B(AES_CORE_DATAPATH__abc_16009_new_n7407_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7408_));
OR2X2 OR2X2_2203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7408_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7409_));
OR2X2 OR2X2_2204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7411_), .B(AES_CORE_DATAPATH__abc_16009_new_n7412_), .Y(AES_CORE_DATAPATH__0key_3__31_0__4_));
OR2X2 OR2X2_2205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7414_));
OR2X2 OR2X2_2206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7415_), .B(AES_CORE_DATAPATH__abc_16009_new_n7416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7417_));
OR2X2 OR2X2_2207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7418_));
OR2X2 OR2X2_2208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7420_), .B(AES_CORE_DATAPATH__abc_16009_new_n7421_), .Y(AES_CORE_DATAPATH__0key_3__31_0__5_));
OR2X2 OR2X2_2209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7423_));
OR2X2 OR2X2_221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2824_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2825_));
OR2X2 OR2X2_2210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7424_), .B(AES_CORE_DATAPATH__abc_16009_new_n7425_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7426_));
OR2X2 OR2X2_2211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7426_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7427_));
OR2X2 OR2X2_2212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7428_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7429_));
OR2X2 OR2X2_2213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7430_));
OR2X2 OR2X2_2214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7432_));
OR2X2 OR2X2_2215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7433_), .B(AES_CORE_DATAPATH__abc_16009_new_n7434_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7435_));
OR2X2 OR2X2_2216 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7435_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7436_));
OR2X2 OR2X2_2217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7437_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7438_));
OR2X2 OR2X2_2218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7439_));
OR2X2 OR2X2_2219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7441_));
OR2X2 OR2X2_222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_DATAPATH__abc_16009_new_n2830_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2831_));
OR2X2 OR2X2_2220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7442_), .B(AES_CORE_DATAPATH__abc_16009_new_n7443_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7444_));
OR2X2 OR2X2_2221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7444_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7445_));
OR2X2 OR2X2_2222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7447_), .B(AES_CORE_DATAPATH__abc_16009_new_n7448_), .Y(AES_CORE_DATAPATH__0key_3__31_0__8_));
OR2X2 OR2X2_2223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7450_));
OR2X2 OR2X2_2224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7451_), .B(AES_CORE_DATAPATH__abc_16009_new_n7452_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7453_));
OR2X2 OR2X2_2225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7453_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7454_));
OR2X2 OR2X2_2226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7456_), .B(AES_CORE_DATAPATH__abc_16009_new_n7457_), .Y(AES_CORE_DATAPATH__0key_3__31_0__9_));
OR2X2 OR2X2_2227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7459_));
OR2X2 OR2X2_2228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7460_), .B(AES_CORE_DATAPATH__abc_16009_new_n7461_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7462_));
OR2X2 OR2X2_2229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7463_));
OR2X2 OR2X2_223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH__abc_16009_new_n2832_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2833_));
OR2X2 OR2X2_2230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7465_), .B(AES_CORE_DATAPATH__abc_16009_new_n7466_), .Y(AES_CORE_DATAPATH__0key_3__31_0__10_));
OR2X2 OR2X2_2231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7468_));
OR2X2 OR2X2_2232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7469_), .B(AES_CORE_DATAPATH__abc_16009_new_n7470_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7471_));
OR2X2 OR2X2_2233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7471_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7472_));
OR2X2 OR2X2_2234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7474_), .B(AES_CORE_DATAPATH__abc_16009_new_n7475_), .Y(AES_CORE_DATAPATH__0key_3__31_0__11_));
OR2X2 OR2X2_2235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7477_));
OR2X2 OR2X2_2236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7478_), .B(AES_CORE_DATAPATH__abc_16009_new_n7479_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7480_));
OR2X2 OR2X2_2237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7480_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7481_));
OR2X2 OR2X2_2238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7483_), .B(AES_CORE_DATAPATH__abc_16009_new_n7484_), .Y(AES_CORE_DATAPATH__0key_3__31_0__12_));
OR2X2 OR2X2_2239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7486_));
OR2X2 OR2X2_224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2834_), .B(AES_CORE_CONTROL_UNIT_bypass_key_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n2835_));
OR2X2 OR2X2_2240 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7487_), .B(AES_CORE_DATAPATH__abc_16009_new_n7488_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7489_));
OR2X2 OR2X2_2241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7489_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7490_));
OR2X2 OR2X2_2242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7492_), .B(AES_CORE_DATAPATH__abc_16009_new_n7493_), .Y(AES_CORE_DATAPATH__0key_3__31_0__13_));
OR2X2 OR2X2_2243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7495_));
OR2X2 OR2X2_2244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7496_), .B(AES_CORE_DATAPATH__abc_16009_new_n7497_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7498_));
OR2X2 OR2X2_2245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7498_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7499_));
OR2X2 OR2X2_2246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7501_), .B(AES_CORE_DATAPATH__abc_16009_new_n7502_), .Y(AES_CORE_DATAPATH__0key_3__31_0__14_));
OR2X2 OR2X2_2247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7504_));
OR2X2 OR2X2_2248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7505_), .B(AES_CORE_DATAPATH__abc_16009_new_n7506_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7507_));
OR2X2 OR2X2_2249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7507_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7508_));
OR2X2 OR2X2_225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2829_), .B(AES_CORE_DATAPATH__abc_16009_new_n2839_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2840_));
OR2X2 OR2X2_2250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7510_), .B(AES_CORE_DATAPATH__abc_16009_new_n7511_), .Y(AES_CORE_DATAPATH__0key_3__31_0__15_));
OR2X2 OR2X2_2251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7513_));
OR2X2 OR2X2_2252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7514_), .B(AES_CORE_DATAPATH__abc_16009_new_n7515_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7516_));
OR2X2 OR2X2_2253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7516_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7517_));
OR2X2 OR2X2_2254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7519_), .B(AES_CORE_DATAPATH__abc_16009_new_n7520_), .Y(AES_CORE_DATAPATH__0key_3__31_0__16_));
OR2X2 OR2X2_2255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7522_));
OR2X2 OR2X2_2256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7523_), .B(AES_CORE_DATAPATH__abc_16009_new_n7524_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7525_));
OR2X2 OR2X2_2257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7525_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7526_));
OR2X2 OR2X2_2258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7527_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7528_));
OR2X2 OR2X2_2259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7529_));
OR2X2 OR2X2_226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2840_), .B(AES_CORE_DATAPATH__abc_16009_new_n2827_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2841_));
OR2X2 OR2X2_2260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7531_));
OR2X2 OR2X2_2261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7532_), .B(AES_CORE_DATAPATH__abc_16009_new_n7533_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7534_));
OR2X2 OR2X2_2262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7534_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7535_));
OR2X2 OR2X2_2263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7536_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7537_));
OR2X2 OR2X2_2264 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7538_));
OR2X2 OR2X2_2265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7540_));
OR2X2 OR2X2_2266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7541_), .B(AES_CORE_DATAPATH__abc_16009_new_n7542_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7543_));
OR2X2 OR2X2_2267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7543_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7544_));
OR2X2 OR2X2_2268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7545_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7546_));
OR2X2 OR2X2_2269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7547_));
OR2X2 OR2X2_227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2845_), .B(AES_CORE_DATAPATH__abc_16009_new_n2843_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2846_));
OR2X2 OR2X2_2270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7549_));
OR2X2 OR2X2_2271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7550_), .B(AES_CORE_DATAPATH__abc_16009_new_n7551_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7552_));
OR2X2 OR2X2_2272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7552_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7553_));
OR2X2 OR2X2_2273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7555_), .B(AES_CORE_DATAPATH__abc_16009_new_n7556_), .Y(AES_CORE_DATAPATH__0key_3__31_0__20_));
OR2X2 OR2X2_2274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7558_));
OR2X2 OR2X2_2275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7559_), .B(AES_CORE_DATAPATH__abc_16009_new_n7560_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7561_));
OR2X2 OR2X2_2276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7561_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7562_));
OR2X2 OR2X2_2277 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7564_), .B(AES_CORE_DATAPATH__abc_16009_new_n7565_), .Y(AES_CORE_DATAPATH__0key_3__31_0__21_));
OR2X2 OR2X2_2278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7567_));
OR2X2 OR2X2_2279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7568_), .B(AES_CORE_DATAPATH__abc_16009_new_n7569_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7570_));
OR2X2 OR2X2_228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2846_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2847_));
OR2X2 OR2X2_2280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7570_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7571_));
OR2X2 OR2X2_2281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7572_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7573_));
OR2X2 OR2X2_2282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7574_));
OR2X2 OR2X2_2283 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7576_));
OR2X2 OR2X2_2284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7577_), .B(AES_CORE_DATAPATH__abc_16009_new_n7578_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7579_));
OR2X2 OR2X2_2285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7579_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7580_));
OR2X2 OR2X2_2286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7581_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7582_));
OR2X2 OR2X2_2287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7583_));
OR2X2 OR2X2_2288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7585_));
OR2X2 OR2X2_2289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7586_), .B(AES_CORE_DATAPATH__abc_16009_new_n7587_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7588_));
OR2X2 OR2X2_229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2849_));
OR2X2 OR2X2_2290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7588_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7589_));
OR2X2 OR2X2_2291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7590_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7591_));
OR2X2 OR2X2_2292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7592_));
OR2X2 OR2X2_2293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7594_));
OR2X2 OR2X2_2294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7595_), .B(AES_CORE_DATAPATH__abc_16009_new_n7596_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7597_));
OR2X2 OR2X2_2295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7597_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7598_));
OR2X2 OR2X2_2296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7599_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7600_));
OR2X2 OR2X2_2297 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7601_));
OR2X2 OR2X2_2298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7603_));
OR2X2 OR2X2_2299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7604_), .B(AES_CORE_DATAPATH__abc_16009_new_n7605_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7606_));
OR2X2 OR2X2_23 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n152_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n153_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n154_));
OR2X2 OR2X2_230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2851_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2852_));
OR2X2 OR2X2_2300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7606_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7607_));
OR2X2 OR2X2_2301 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7608_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7609_));
OR2X2 OR2X2_2302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7610_));
OR2X2 OR2X2_2303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7612_));
OR2X2 OR2X2_2304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7613_), .B(AES_CORE_DATAPATH__abc_16009_new_n7614_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7615_));
OR2X2 OR2X2_2305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7615_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7616_));
OR2X2 OR2X2_2306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7618_), .B(AES_CORE_DATAPATH__abc_16009_new_n7619_), .Y(AES_CORE_DATAPATH__0key_3__31_0__27_));
OR2X2 OR2X2_2307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7621_));
OR2X2 OR2X2_2308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7622_), .B(AES_CORE_DATAPATH__abc_16009_new_n7623_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7624_));
OR2X2 OR2X2_2309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7624_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7625_));
OR2X2 OR2X2_231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2855_), .B(AES_CORE_DATAPATH__abc_16009_new_n2856_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2857_));
OR2X2 OR2X2_2310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7627_), .B(AES_CORE_DATAPATH__abc_16009_new_n7628_), .Y(AES_CORE_DATAPATH__0key_3__31_0__28_));
OR2X2 OR2X2_2311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7630_));
OR2X2 OR2X2_2312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7631_), .B(AES_CORE_DATAPATH__abc_16009_new_n7632_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7633_));
OR2X2 OR2X2_2313 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7634_));
OR2X2 OR2X2_2314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7635_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7636_));
OR2X2 OR2X2_2315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7637_));
OR2X2 OR2X2_2316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7639_));
OR2X2 OR2X2_2317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7640_), .B(AES_CORE_DATAPATH__abc_16009_new_n7641_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7642_));
OR2X2 OR2X2_2318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7643_));
OR2X2 OR2X2_2319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7645_), .B(AES_CORE_DATAPATH__abc_16009_new_n7646_), .Y(AES_CORE_DATAPATH__0key_3__31_0__30_));
OR2X2 OR2X2_232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2857_), .B(AES_CORE_DATAPATH__abc_16009_new_n2854_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2858_));
OR2X2 OR2X2_2320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7648_));
OR2X2 OR2X2_2321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7649_), .B(AES_CORE_DATAPATH__abc_16009_new_n7650_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7651_));
OR2X2 OR2X2_2322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n7651_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7652_));
OR2X2 OR2X2_2323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7653_), .B(AES_CORE_DATAPATH__abc_16009_new_n7367_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7654_));
OR2X2 OR2X2_2324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7655_));
OR2X2 OR2X2_2325 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7658_), .B(AES_CORE_DATAPATH__abc_16009_new_n7657_), .Y(AES_CORE_DATAPATH__0key_host_3__31_0__0_));
OR2X2 OR2X2_2326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7381_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7660_));
OR2X2 OR2X2_2327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7661_));
OR2X2 OR2X2_2328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7390_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7663_));
OR2X2 OR2X2_2329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7664_));
OR2X2 OR2X2_233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2859_));
OR2X2 OR2X2_2330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7399_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7666_));
OR2X2 OR2X2_2331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7667_));
OR2X2 OR2X2_2332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7408_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7669_));
OR2X2 OR2X2_2333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7670_));
OR2X2 OR2X2_2334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7417_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7672_));
OR2X2 OR2X2_2335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7673_));
OR2X2 OR2X2_2336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7426_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7675_));
OR2X2 OR2X2_2337 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7676_));
OR2X2 OR2X2_2338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7435_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7678_));
OR2X2 OR2X2_2339 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7679_));
OR2X2 OR2X2_234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2863_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2864_));
OR2X2 OR2X2_2340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7444_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7681_));
OR2X2 OR2X2_2341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7682_));
OR2X2 OR2X2_2342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7453_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7684_));
OR2X2 OR2X2_2343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7685_));
OR2X2 OR2X2_2344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7462_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7687_));
OR2X2 OR2X2_2345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7688_));
OR2X2 OR2X2_2346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7471_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7690_));
OR2X2 OR2X2_2347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7691_));
OR2X2 OR2X2_2348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7480_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7693_));
OR2X2 OR2X2_2349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7694_));
OR2X2 OR2X2_235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2864_), .B(AES_CORE_DATAPATH__abc_16009_new_n2861_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2865_));
OR2X2 OR2X2_2350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7489_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7696_));
OR2X2 OR2X2_2351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7697_));
OR2X2 OR2X2_2352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7498_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7699_));
OR2X2 OR2X2_2353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7700_));
OR2X2 OR2X2_2354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7507_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7702_));
OR2X2 OR2X2_2355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7703_));
OR2X2 OR2X2_2356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7516_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7705_));
OR2X2 OR2X2_2357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7706_));
OR2X2 OR2X2_2358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7525_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7708_));
OR2X2 OR2X2_2359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7709_));
OR2X2 OR2X2_236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2867_));
OR2X2 OR2X2_2360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7534_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7711_));
OR2X2 OR2X2_2361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7712_));
OR2X2 OR2X2_2362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7543_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7714_));
OR2X2 OR2X2_2363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7715_));
OR2X2 OR2X2_2364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7552_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7717_));
OR2X2 OR2X2_2365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7718_));
OR2X2 OR2X2_2366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7561_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7720_));
OR2X2 OR2X2_2367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7721_));
OR2X2 OR2X2_2368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7570_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7723_));
OR2X2 OR2X2_2369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7724_));
OR2X2 OR2X2_237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2869_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2870_));
OR2X2 OR2X2_2370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7579_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7726_));
OR2X2 OR2X2_2371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7727_));
OR2X2 OR2X2_2372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7588_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7729_));
OR2X2 OR2X2_2373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7730_));
OR2X2 OR2X2_2374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7597_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7732_));
OR2X2 OR2X2_2375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7733_));
OR2X2 OR2X2_2376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7606_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7735_));
OR2X2 OR2X2_2377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7736_));
OR2X2 OR2X2_2378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7615_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7738_));
OR2X2 OR2X2_2379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7739_));
OR2X2 OR2X2_238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2873_), .B(AES_CORE_DATAPATH__abc_16009_new_n2874_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2875_));
OR2X2 OR2X2_2380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7624_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7741_));
OR2X2 OR2X2_2381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7742_));
OR2X2 OR2X2_2382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7633_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7744_));
OR2X2 OR2X2_2383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7745_));
OR2X2 OR2X2_2384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7642_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7747_));
OR2X2 OR2X2_2385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7748_));
OR2X2 OR2X2_2386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5155_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7750_));
OR2X2 OR2X2_2387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7651_), .B(AES_CORE_CONTROL_UNIT_key_derivation_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n7751_));
OR2X2 OR2X2_2388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7755_), .B(AES_CORE_DATAPATH__abc_16009_new_n7756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7757_));
OR2X2 OR2X2_2389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5807_), .B(AES_CORE_DATAPATH__abc_16009_new_n7758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7759_));
OR2X2 OR2X2_239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2875_), .B(AES_CORE_DATAPATH__abc_16009_new_n2872_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2876_));
OR2X2 OR2X2_2390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7760_), .B(AES_CORE_DATAPATH__abc_16009_new_n7754_), .Y(AES_CORE_DATAPATH__0col_3__31_0__0_));
OR2X2 OR2X2_2391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7763_), .B(AES_CORE_DATAPATH__abc_16009_new_n7764_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7765_));
OR2X2 OR2X2_2392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5857_), .B(AES_CORE_DATAPATH__abc_16009_new_n7766_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7767_));
OR2X2 OR2X2_2393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7768_), .B(AES_CORE_DATAPATH__abc_16009_new_n7762_), .Y(AES_CORE_DATAPATH__0col_3__31_0__1_));
OR2X2 OR2X2_2394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7771_), .B(AES_CORE_DATAPATH__abc_16009_new_n7772_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7773_));
OR2X2 OR2X2_2395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5907_), .B(AES_CORE_DATAPATH__abc_16009_new_n7774_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7775_));
OR2X2 OR2X2_2396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7776_), .B(AES_CORE_DATAPATH__abc_16009_new_n7770_), .Y(AES_CORE_DATAPATH__0col_3__31_0__2_));
OR2X2 OR2X2_2397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7779_), .B(AES_CORE_DATAPATH__abc_16009_new_n7780_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7781_));
OR2X2 OR2X2_2398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5957_), .B(AES_CORE_DATAPATH__abc_16009_new_n7782_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7783_));
OR2X2 OR2X2_2399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7784_), .B(AES_CORE_DATAPATH__abc_16009_new_n7778_), .Y(AES_CORE_DATAPATH__0col_3__31_0__3_));
OR2X2 OR2X2_24 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n157_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n156_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_12_));
OR2X2 OR2X2_240 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2877_));
OR2X2 OR2X2_2400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7787_), .B(AES_CORE_DATAPATH__abc_16009_new_n7788_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7789_));
OR2X2 OR2X2_2401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6007_), .B(AES_CORE_DATAPATH__abc_16009_new_n7790_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7791_));
OR2X2 OR2X2_2402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7792_), .B(AES_CORE_DATAPATH__abc_16009_new_n7786_), .Y(AES_CORE_DATAPATH__0col_3__31_0__4_));
OR2X2 OR2X2_2403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7795_), .B(AES_CORE_DATAPATH__abc_16009_new_n7796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7797_));
OR2X2 OR2X2_2404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6057_), .B(AES_CORE_DATAPATH__abc_16009_new_n7798_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7799_));
OR2X2 OR2X2_2405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7800_), .B(AES_CORE_DATAPATH__abc_16009_new_n7794_), .Y(AES_CORE_DATAPATH__0col_3__31_0__5_));
OR2X2 OR2X2_2406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7803_), .B(AES_CORE_DATAPATH__abc_16009_new_n7804_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7805_));
OR2X2 OR2X2_2407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6107_), .B(AES_CORE_DATAPATH__abc_16009_new_n7806_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7807_));
OR2X2 OR2X2_2408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7808_), .B(AES_CORE_DATAPATH__abc_16009_new_n7802_), .Y(AES_CORE_DATAPATH__0col_3__31_0__6_));
OR2X2 OR2X2_2409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7811_), .B(AES_CORE_DATAPATH__abc_16009_new_n7812_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7813_));
OR2X2 OR2X2_241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2881_), .B(AES_CORE_DATAPATH__abc_16009_new_n2879_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2882_));
OR2X2 OR2X2_2410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6157_), .B(AES_CORE_DATAPATH__abc_16009_new_n7814_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7815_));
OR2X2 OR2X2_2411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7816_), .B(AES_CORE_DATAPATH__abc_16009_new_n7810_), .Y(AES_CORE_DATAPATH__0col_3__31_0__7_));
OR2X2 OR2X2_2412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7819_), .B(AES_CORE_DATAPATH__abc_16009_new_n7820_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7821_));
OR2X2 OR2X2_2413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6207_), .B(AES_CORE_DATAPATH__abc_16009_new_n7822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7823_));
OR2X2 OR2X2_2414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7824_), .B(AES_CORE_DATAPATH__abc_16009_new_n7818_), .Y(AES_CORE_DATAPATH__0col_3__31_0__8_));
OR2X2 OR2X2_2415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7827_), .B(AES_CORE_DATAPATH__abc_16009_new_n7828_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7829_));
OR2X2 OR2X2_2416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6257_), .B(AES_CORE_DATAPATH__abc_16009_new_n7830_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7831_));
OR2X2 OR2X2_2417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7832_), .B(AES_CORE_DATAPATH__abc_16009_new_n7826_), .Y(AES_CORE_DATAPATH__0col_3__31_0__9_));
OR2X2 OR2X2_2418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7835_), .B(AES_CORE_DATAPATH__abc_16009_new_n7836_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7837_));
OR2X2 OR2X2_2419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6307_), .B(AES_CORE_DATAPATH__abc_16009_new_n7838_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7839_));
OR2X2 OR2X2_242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2882_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2883_));
OR2X2 OR2X2_2420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7840_), .B(AES_CORE_DATAPATH__abc_16009_new_n7834_), .Y(AES_CORE_DATAPATH__0col_3__31_0__10_));
OR2X2 OR2X2_2421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7843_), .B(AES_CORE_DATAPATH__abc_16009_new_n7844_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7845_));
OR2X2 OR2X2_2422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6357_), .B(AES_CORE_DATAPATH__abc_16009_new_n7846_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7847_));
OR2X2 OR2X2_2423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7848_), .B(AES_CORE_DATAPATH__abc_16009_new_n7842_), .Y(AES_CORE_DATAPATH__0col_3__31_0__11_));
OR2X2 OR2X2_2424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7851_), .B(AES_CORE_DATAPATH__abc_16009_new_n7852_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7853_));
OR2X2 OR2X2_2425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6407_), .B(AES_CORE_DATAPATH__abc_16009_new_n7854_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7855_));
OR2X2 OR2X2_2426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7856_), .B(AES_CORE_DATAPATH__abc_16009_new_n7850_), .Y(AES_CORE_DATAPATH__0col_3__31_0__12_));
OR2X2 OR2X2_2427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7859_), .B(AES_CORE_DATAPATH__abc_16009_new_n7860_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7861_));
OR2X2 OR2X2_2428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6457_), .B(AES_CORE_DATAPATH__abc_16009_new_n7862_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7863_));
OR2X2 OR2X2_2429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7864_), .B(AES_CORE_DATAPATH__abc_16009_new_n7858_), .Y(AES_CORE_DATAPATH__0col_3__31_0__13_));
OR2X2 OR2X2_243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2885_));
OR2X2 OR2X2_2430 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7867_), .B(AES_CORE_DATAPATH__abc_16009_new_n7868_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7869_));
OR2X2 OR2X2_2431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6507_), .B(AES_CORE_DATAPATH__abc_16009_new_n7870_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7871_));
OR2X2 OR2X2_2432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7872_), .B(AES_CORE_DATAPATH__abc_16009_new_n7866_), .Y(AES_CORE_DATAPATH__0col_3__31_0__14_));
OR2X2 OR2X2_2433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7875_), .B(AES_CORE_DATAPATH__abc_16009_new_n7876_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7877_));
OR2X2 OR2X2_2434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6557_), .B(AES_CORE_DATAPATH__abc_16009_new_n7878_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7879_));
OR2X2 OR2X2_2435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7880_), .B(AES_CORE_DATAPATH__abc_16009_new_n7874_), .Y(AES_CORE_DATAPATH__0col_3__31_0__15_));
OR2X2 OR2X2_2436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7883_), .B(AES_CORE_DATAPATH__abc_16009_new_n7884_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7885_));
OR2X2 OR2X2_2437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6607_), .B(AES_CORE_DATAPATH__abc_16009_new_n7886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7887_));
OR2X2 OR2X2_2438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7888_), .B(AES_CORE_DATAPATH__abc_16009_new_n7882_), .Y(AES_CORE_DATAPATH__0col_3__31_0__16_));
OR2X2 OR2X2_2439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7891_), .B(AES_CORE_DATAPATH__abc_16009_new_n7892_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7893_));
OR2X2 OR2X2_244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2887_));
OR2X2 OR2X2_2440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6657_), .B(AES_CORE_DATAPATH__abc_16009_new_n7894_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7895_));
OR2X2 OR2X2_2441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7896_), .B(AES_CORE_DATAPATH__abc_16009_new_n7890_), .Y(AES_CORE_DATAPATH__0col_3__31_0__17_));
OR2X2 OR2X2_2442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7899_), .B(AES_CORE_DATAPATH__abc_16009_new_n7900_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7901_));
OR2X2 OR2X2_2443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6707_), .B(AES_CORE_DATAPATH__abc_16009_new_n7902_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7903_));
OR2X2 OR2X2_2444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7904_), .B(AES_CORE_DATAPATH__abc_16009_new_n7898_), .Y(AES_CORE_DATAPATH__0col_3__31_0__18_));
OR2X2 OR2X2_2445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7907_), .B(AES_CORE_DATAPATH__abc_16009_new_n7908_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7909_));
OR2X2 OR2X2_2446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6757_), .B(AES_CORE_DATAPATH__abc_16009_new_n7910_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7911_));
OR2X2 OR2X2_2447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7912_), .B(AES_CORE_DATAPATH__abc_16009_new_n7906_), .Y(AES_CORE_DATAPATH__0col_3__31_0__19_));
OR2X2 OR2X2_2448 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7915_), .B(AES_CORE_DATAPATH__abc_16009_new_n7916_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7917_));
OR2X2 OR2X2_2449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6807_), .B(AES_CORE_DATAPATH__abc_16009_new_n7918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7919_));
OR2X2 OR2X2_245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2888_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2889_));
OR2X2 OR2X2_2450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7920_), .B(AES_CORE_DATAPATH__abc_16009_new_n7914_), .Y(AES_CORE_DATAPATH__0col_3__31_0__20_));
OR2X2 OR2X2_2451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7923_), .B(AES_CORE_DATAPATH__abc_16009_new_n7924_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7925_));
OR2X2 OR2X2_2452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6857_), .B(AES_CORE_DATAPATH__abc_16009_new_n7926_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7927_));
OR2X2 OR2X2_2453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7928_), .B(AES_CORE_DATAPATH__abc_16009_new_n7922_), .Y(AES_CORE_DATAPATH__0col_3__31_0__21_));
OR2X2 OR2X2_2454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7931_), .B(AES_CORE_DATAPATH__abc_16009_new_n7932_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7933_));
OR2X2 OR2X2_2455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6907_), .B(AES_CORE_DATAPATH__abc_16009_new_n7934_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7935_));
OR2X2 OR2X2_2456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7936_), .B(AES_CORE_DATAPATH__abc_16009_new_n7930_), .Y(AES_CORE_DATAPATH__0col_3__31_0__22_));
OR2X2 OR2X2_2457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7939_), .B(AES_CORE_DATAPATH__abc_16009_new_n7940_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7941_));
OR2X2 OR2X2_2458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6957_), .B(AES_CORE_DATAPATH__abc_16009_new_n7942_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7943_));
OR2X2 OR2X2_2459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7944_), .B(AES_CORE_DATAPATH__abc_16009_new_n7938_), .Y(AES_CORE_DATAPATH__0col_3__31_0__23_));
OR2X2 OR2X2_246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2892_), .B(AES_CORE_DATAPATH__abc_16009_new_n2893_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2894_));
OR2X2 OR2X2_2460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7947_), .B(AES_CORE_DATAPATH__abc_16009_new_n7948_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7949_));
OR2X2 OR2X2_2461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7007_), .B(AES_CORE_DATAPATH__abc_16009_new_n7950_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7951_));
OR2X2 OR2X2_2462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7952_), .B(AES_CORE_DATAPATH__abc_16009_new_n7946_), .Y(AES_CORE_DATAPATH__0col_3__31_0__24_));
OR2X2 OR2X2_2463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7955_), .B(AES_CORE_DATAPATH__abc_16009_new_n7956_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7957_));
OR2X2 OR2X2_2464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7057_), .B(AES_CORE_DATAPATH__abc_16009_new_n7958_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7959_));
OR2X2 OR2X2_2465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7960_), .B(AES_CORE_DATAPATH__abc_16009_new_n7954_), .Y(AES_CORE_DATAPATH__0col_3__31_0__25_));
OR2X2 OR2X2_2466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7963_), .B(AES_CORE_DATAPATH__abc_16009_new_n7964_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7965_));
OR2X2 OR2X2_2467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7107_), .B(AES_CORE_DATAPATH__abc_16009_new_n7966_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7967_));
OR2X2 OR2X2_2468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7968_), .B(AES_CORE_DATAPATH__abc_16009_new_n7962_), .Y(AES_CORE_DATAPATH__0col_3__31_0__26_));
OR2X2 OR2X2_2469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7971_), .B(AES_CORE_DATAPATH__abc_16009_new_n7972_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7973_));
OR2X2 OR2X2_247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2894_), .B(AES_CORE_DATAPATH__abc_16009_new_n2891_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2895_));
OR2X2 OR2X2_2470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7157_), .B(AES_CORE_DATAPATH__abc_16009_new_n7974_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7975_));
OR2X2 OR2X2_2471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7976_), .B(AES_CORE_DATAPATH__abc_16009_new_n7970_), .Y(AES_CORE_DATAPATH__0col_3__31_0__27_));
OR2X2 OR2X2_2472 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7979_), .B(AES_CORE_DATAPATH__abc_16009_new_n7980_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7981_));
OR2X2 OR2X2_2473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7207_), .B(AES_CORE_DATAPATH__abc_16009_new_n7982_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7983_));
OR2X2 OR2X2_2474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7984_), .B(AES_CORE_DATAPATH__abc_16009_new_n7978_), .Y(AES_CORE_DATAPATH__0col_3__31_0__28_));
OR2X2 OR2X2_2475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7987_), .B(AES_CORE_DATAPATH__abc_16009_new_n7988_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7989_));
OR2X2 OR2X2_2476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7257_), .B(AES_CORE_DATAPATH__abc_16009_new_n7990_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7991_));
OR2X2 OR2X2_2477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7992_), .B(AES_CORE_DATAPATH__abc_16009_new_n7986_), .Y(AES_CORE_DATAPATH__0col_3__31_0__29_));
OR2X2 OR2X2_2478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7995_), .B(AES_CORE_DATAPATH__abc_16009_new_n7996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7997_));
OR2X2 OR2X2_2479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7307_), .B(AES_CORE_DATAPATH__abc_16009_new_n7998_), .Y(AES_CORE_DATAPATH__abc_16009_new_n7999_));
OR2X2 OR2X2_248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2899_), .B(AES_CORE_DATAPATH__abc_16009_new_n2897_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2900_));
OR2X2 OR2X2_2480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8000_), .B(AES_CORE_DATAPATH__abc_16009_new_n7994_), .Y(AES_CORE_DATAPATH__0col_3__31_0__30_));
OR2X2 OR2X2_2481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8003_), .B(AES_CORE_DATAPATH__abc_16009_new_n8004_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8005_));
OR2X2 OR2X2_2482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7357_), .B(AES_CORE_DATAPATH__abc_16009_new_n8006_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8007_));
OR2X2 OR2X2_2483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8008_), .B(AES_CORE_DATAPATH__abc_16009_new_n8002_), .Y(AES_CORE_DATAPATH__0col_3__31_0__31_));
OR2X2 OR2X2_2484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8012_), .B(AES_CORE_DATAPATH__abc_16009_new_n8013_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8014_));
OR2X2 OR2X2_2485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5807_), .B(AES_CORE_DATAPATH__abc_16009_new_n8015_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8016_));
OR2X2 OR2X2_2486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8017_), .B(AES_CORE_DATAPATH__abc_16009_new_n8011_), .Y(AES_CORE_DATAPATH__0col_1__31_0__0_));
OR2X2 OR2X2_2487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8020_), .B(AES_CORE_DATAPATH__abc_16009_new_n8021_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8022_));
OR2X2 OR2X2_2488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8023_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8024_));
OR2X2 OR2X2_2489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8025_), .B(AES_CORE_DATAPATH__abc_16009_new_n8019_), .Y(AES_CORE_DATAPATH__0col_1__31_0__1_));
OR2X2 OR2X2_249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2900_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2901_));
OR2X2 OR2X2_2490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8028_), .B(AES_CORE_DATAPATH__abc_16009_new_n8029_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8030_));
OR2X2 OR2X2_2491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5907_), .B(AES_CORE_DATAPATH__abc_16009_new_n8031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8032_));
OR2X2 OR2X2_2492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8033_), .B(AES_CORE_DATAPATH__abc_16009_new_n8027_), .Y(AES_CORE_DATAPATH__0col_1__31_0__2_));
OR2X2 OR2X2_2493 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8036_), .B(AES_CORE_DATAPATH__abc_16009_new_n8037_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8038_));
OR2X2 OR2X2_2494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5957_), .B(AES_CORE_DATAPATH__abc_16009_new_n8039_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8040_));
OR2X2 OR2X2_2495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8041_), .B(AES_CORE_DATAPATH__abc_16009_new_n8035_), .Y(AES_CORE_DATAPATH__0col_1__31_0__3_));
OR2X2 OR2X2_2496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8044_), .B(AES_CORE_DATAPATH__abc_16009_new_n8045_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8046_));
OR2X2 OR2X2_2497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6007_), .B(AES_CORE_DATAPATH__abc_16009_new_n8047_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8048_));
OR2X2 OR2X2_2498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8049_), .B(AES_CORE_DATAPATH__abc_16009_new_n8043_), .Y(AES_CORE_DATAPATH__0col_1__31_0__4_));
OR2X2 OR2X2_2499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8052_), .B(AES_CORE_DATAPATH__abc_16009_new_n8053_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8054_));
OR2X2 OR2X2_25 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n161_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n159_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_13_));
OR2X2 OR2X2_250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2903_));
OR2X2 OR2X2_2500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6057_), .B(AES_CORE_DATAPATH__abc_16009_new_n8055_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8056_));
OR2X2 OR2X2_2501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8057_), .B(AES_CORE_DATAPATH__abc_16009_new_n8051_), .Y(AES_CORE_DATAPATH__0col_1__31_0__5_));
OR2X2 OR2X2_2502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8060_), .B(AES_CORE_DATAPATH__abc_16009_new_n8061_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8062_));
OR2X2 OR2X2_2503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6107_), .B(AES_CORE_DATAPATH__abc_16009_new_n8063_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8064_));
OR2X2 OR2X2_2504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8065_), .B(AES_CORE_DATAPATH__abc_16009_new_n8059_), .Y(AES_CORE_DATAPATH__0col_1__31_0__6_));
OR2X2 OR2X2_2505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8068_), .B(AES_CORE_DATAPATH__abc_16009_new_n8069_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8070_));
OR2X2 OR2X2_2506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6157_), .B(AES_CORE_DATAPATH__abc_16009_new_n8071_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8072_));
OR2X2 OR2X2_2507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8073_), .B(AES_CORE_DATAPATH__abc_16009_new_n8067_), .Y(AES_CORE_DATAPATH__0col_1__31_0__7_));
OR2X2 OR2X2_2508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8076_), .B(AES_CORE_DATAPATH__abc_16009_new_n8077_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8078_));
OR2X2 OR2X2_2509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6207_), .B(AES_CORE_DATAPATH__abc_16009_new_n8079_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8080_));
OR2X2 OR2X2_251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2905_));
OR2X2 OR2X2_2510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8081_), .B(AES_CORE_DATAPATH__abc_16009_new_n8075_), .Y(AES_CORE_DATAPATH__0col_1__31_0__8_));
OR2X2 OR2X2_2511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8084_), .B(AES_CORE_DATAPATH__abc_16009_new_n8085_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8086_));
OR2X2 OR2X2_2512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6257_), .B(AES_CORE_DATAPATH__abc_16009_new_n8087_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8088_));
OR2X2 OR2X2_2513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8089_), .B(AES_CORE_DATAPATH__abc_16009_new_n8083_), .Y(AES_CORE_DATAPATH__0col_1__31_0__9_));
OR2X2 OR2X2_2514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8092_), .B(AES_CORE_DATAPATH__abc_16009_new_n8093_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8094_));
OR2X2 OR2X2_2515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6307_), .B(AES_CORE_DATAPATH__abc_16009_new_n8095_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8096_));
OR2X2 OR2X2_2516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8097_), .B(AES_CORE_DATAPATH__abc_16009_new_n8091_), .Y(AES_CORE_DATAPATH__0col_1__31_0__10_));
OR2X2 OR2X2_2517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8100_), .B(AES_CORE_DATAPATH__abc_16009_new_n8101_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8102_));
OR2X2 OR2X2_2518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6357_), .B(AES_CORE_DATAPATH__abc_16009_new_n8103_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8104_));
OR2X2 OR2X2_2519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8105_), .B(AES_CORE_DATAPATH__abc_16009_new_n8099_), .Y(AES_CORE_DATAPATH__0col_1__31_0__11_));
OR2X2 OR2X2_252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2906_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2907_));
OR2X2 OR2X2_2520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8108_), .B(AES_CORE_DATAPATH__abc_16009_new_n8109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8110_));
OR2X2 OR2X2_2521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6407_), .B(AES_CORE_DATAPATH__abc_16009_new_n8111_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8112_));
OR2X2 OR2X2_2522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8113_), .B(AES_CORE_DATAPATH__abc_16009_new_n8107_), .Y(AES_CORE_DATAPATH__0col_1__31_0__12_));
OR2X2 OR2X2_2523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8116_), .B(AES_CORE_DATAPATH__abc_16009_new_n8117_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8118_));
OR2X2 OR2X2_2524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6457_), .B(AES_CORE_DATAPATH__abc_16009_new_n8119_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8120_));
OR2X2 OR2X2_2525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8121_), .B(AES_CORE_DATAPATH__abc_16009_new_n8115_), .Y(AES_CORE_DATAPATH__0col_1__31_0__13_));
OR2X2 OR2X2_2526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8124_), .B(AES_CORE_DATAPATH__abc_16009_new_n8125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8126_));
OR2X2 OR2X2_2527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6507_), .B(AES_CORE_DATAPATH__abc_16009_new_n8127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8128_));
OR2X2 OR2X2_2528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8129_), .B(AES_CORE_DATAPATH__abc_16009_new_n8123_), .Y(AES_CORE_DATAPATH__0col_1__31_0__14_));
OR2X2 OR2X2_2529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8132_), .B(AES_CORE_DATAPATH__abc_16009_new_n8133_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8134_));
OR2X2 OR2X2_253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2910_), .B(AES_CORE_DATAPATH__abc_16009_new_n2911_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2912_));
OR2X2 OR2X2_2530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6557_), .B(AES_CORE_DATAPATH__abc_16009_new_n8135_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8136_));
OR2X2 OR2X2_2531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8137_), .B(AES_CORE_DATAPATH__abc_16009_new_n8131_), .Y(AES_CORE_DATAPATH__0col_1__31_0__15_));
OR2X2 OR2X2_2532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8140_), .B(AES_CORE_DATAPATH__abc_16009_new_n8141_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8142_));
OR2X2 OR2X2_2533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6607_), .B(AES_CORE_DATAPATH__abc_16009_new_n8143_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8144_));
OR2X2 OR2X2_2534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8145_), .B(AES_CORE_DATAPATH__abc_16009_new_n8139_), .Y(AES_CORE_DATAPATH__0col_1__31_0__16_));
OR2X2 OR2X2_2535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8148_), .B(AES_CORE_DATAPATH__abc_16009_new_n8149_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8150_));
OR2X2 OR2X2_2536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6657_), .B(AES_CORE_DATAPATH__abc_16009_new_n8151_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8152_));
OR2X2 OR2X2_2537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8153_), .B(AES_CORE_DATAPATH__abc_16009_new_n8147_), .Y(AES_CORE_DATAPATH__0col_1__31_0__17_));
OR2X2 OR2X2_2538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8156_), .B(AES_CORE_DATAPATH__abc_16009_new_n8157_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8158_));
OR2X2 OR2X2_2539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6707_), .B(AES_CORE_DATAPATH__abc_16009_new_n8159_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8160_));
OR2X2 OR2X2_254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2912_), .B(AES_CORE_DATAPATH__abc_16009_new_n2909_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2913_));
OR2X2 OR2X2_2540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8161_), .B(AES_CORE_DATAPATH__abc_16009_new_n8155_), .Y(AES_CORE_DATAPATH__0col_1__31_0__18_));
OR2X2 OR2X2_2541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8164_), .B(AES_CORE_DATAPATH__abc_16009_new_n8165_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8166_));
OR2X2 OR2X2_2542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6757_), .B(AES_CORE_DATAPATH__abc_16009_new_n8167_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8168_));
OR2X2 OR2X2_2543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8169_), .B(AES_CORE_DATAPATH__abc_16009_new_n8163_), .Y(AES_CORE_DATAPATH__0col_1__31_0__19_));
OR2X2 OR2X2_2544 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8172_), .B(AES_CORE_DATAPATH__abc_16009_new_n8173_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8174_));
OR2X2 OR2X2_2545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6807_), .B(AES_CORE_DATAPATH__abc_16009_new_n8175_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8176_));
OR2X2 OR2X2_2546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8177_), .B(AES_CORE_DATAPATH__abc_16009_new_n8171_), .Y(AES_CORE_DATAPATH__0col_1__31_0__20_));
OR2X2 OR2X2_2547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8180_), .B(AES_CORE_DATAPATH__abc_16009_new_n8181_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8182_));
OR2X2 OR2X2_2548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8183_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8184_));
OR2X2 OR2X2_2549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8185_), .B(AES_CORE_DATAPATH__abc_16009_new_n8179_), .Y(AES_CORE_DATAPATH__0col_1__31_0__21_));
OR2X2 OR2X2_255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2917_), .B(AES_CORE_DATAPATH__abc_16009_new_n2915_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2918_));
OR2X2 OR2X2_2550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8188_), .B(AES_CORE_DATAPATH__abc_16009_new_n8189_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8190_));
OR2X2 OR2X2_2551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6907_), .B(AES_CORE_DATAPATH__abc_16009_new_n8191_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8192_));
OR2X2 OR2X2_2552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8193_), .B(AES_CORE_DATAPATH__abc_16009_new_n8187_), .Y(AES_CORE_DATAPATH__0col_1__31_0__22_));
OR2X2 OR2X2_2553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8196_), .B(AES_CORE_DATAPATH__abc_16009_new_n8197_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8198_));
OR2X2 OR2X2_2554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6957_), .B(AES_CORE_DATAPATH__abc_16009_new_n8199_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8200_));
OR2X2 OR2X2_2555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8201_), .B(AES_CORE_DATAPATH__abc_16009_new_n8195_), .Y(AES_CORE_DATAPATH__0col_1__31_0__23_));
OR2X2 OR2X2_2556 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8204_), .B(AES_CORE_DATAPATH__abc_16009_new_n8205_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8206_));
OR2X2 OR2X2_2557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7007_), .B(AES_CORE_DATAPATH__abc_16009_new_n8207_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8208_));
OR2X2 OR2X2_2558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8209_), .B(AES_CORE_DATAPATH__abc_16009_new_n8203_), .Y(AES_CORE_DATAPATH__0col_1__31_0__24_));
OR2X2 OR2X2_2559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8212_), .B(AES_CORE_DATAPATH__abc_16009_new_n8213_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8214_));
OR2X2 OR2X2_256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2918_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2919_));
OR2X2 OR2X2_2560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7057_), .B(AES_CORE_DATAPATH__abc_16009_new_n8215_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8216_));
OR2X2 OR2X2_2561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8217_), .B(AES_CORE_DATAPATH__abc_16009_new_n8211_), .Y(AES_CORE_DATAPATH__0col_1__31_0__25_));
OR2X2 OR2X2_2562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8220_), .B(AES_CORE_DATAPATH__abc_16009_new_n8221_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8222_));
OR2X2 OR2X2_2563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7107_), .B(AES_CORE_DATAPATH__abc_16009_new_n8223_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8224_));
OR2X2 OR2X2_2564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8225_), .B(AES_CORE_DATAPATH__abc_16009_new_n8219_), .Y(AES_CORE_DATAPATH__0col_1__31_0__26_));
OR2X2 OR2X2_2565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8228_), .B(AES_CORE_DATAPATH__abc_16009_new_n8229_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8230_));
OR2X2 OR2X2_2566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7157_), .B(AES_CORE_DATAPATH__abc_16009_new_n8231_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8232_));
OR2X2 OR2X2_2567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8233_), .B(AES_CORE_DATAPATH__abc_16009_new_n8227_), .Y(AES_CORE_DATAPATH__0col_1__31_0__27_));
OR2X2 OR2X2_2568 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8236_), .B(AES_CORE_DATAPATH__abc_16009_new_n8237_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8238_));
OR2X2 OR2X2_2569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7207_), .B(AES_CORE_DATAPATH__abc_16009_new_n8239_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8240_));
OR2X2 OR2X2_257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2921_));
OR2X2 OR2X2_2570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8241_), .B(AES_CORE_DATAPATH__abc_16009_new_n8235_), .Y(AES_CORE_DATAPATH__0col_1__31_0__28_));
OR2X2 OR2X2_2571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8244_), .B(AES_CORE_DATAPATH__abc_16009_new_n8245_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8246_));
OR2X2 OR2X2_2572 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7257_), .B(AES_CORE_DATAPATH__abc_16009_new_n8247_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8248_));
OR2X2 OR2X2_2573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8249_), .B(AES_CORE_DATAPATH__abc_16009_new_n8243_), .Y(AES_CORE_DATAPATH__0col_1__31_0__29_));
OR2X2 OR2X2_2574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8252_), .B(AES_CORE_DATAPATH__abc_16009_new_n8253_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8254_));
OR2X2 OR2X2_2575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7307_), .B(AES_CORE_DATAPATH__abc_16009_new_n8255_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8256_));
OR2X2 OR2X2_2576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8257_), .B(AES_CORE_DATAPATH__abc_16009_new_n8251_), .Y(AES_CORE_DATAPATH__0col_1__31_0__30_));
OR2X2 OR2X2_2577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8260_), .B(AES_CORE_DATAPATH__abc_16009_new_n8261_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8262_));
OR2X2 OR2X2_2578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7357_), .B(AES_CORE_DATAPATH__abc_16009_new_n8263_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8264_));
OR2X2 OR2X2_2579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8265_), .B(AES_CORE_DATAPATH__abc_16009_new_n8259_), .Y(AES_CORE_DATAPATH__0col_1__31_0__31_));
OR2X2 OR2X2_258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2923_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2924_));
OR2X2 OR2X2_2580 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8269_), .B(AES_CORE_DATAPATH__abc_16009_new_n8270_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8271_));
OR2X2 OR2X2_2581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5807_), .B(AES_CORE_DATAPATH__abc_16009_new_n8272_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8273_));
OR2X2 OR2X2_2582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8274_), .B(AES_CORE_DATAPATH__abc_16009_new_n8268_), .Y(AES_CORE_DATAPATH__0col_2__31_0__0_));
OR2X2 OR2X2_2583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8277_), .B(AES_CORE_DATAPATH__abc_16009_new_n8278_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8279_));
OR2X2 OR2X2_2584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8280_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8281_));
OR2X2 OR2X2_2585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8282_), .B(AES_CORE_DATAPATH__abc_16009_new_n8276_), .Y(AES_CORE_DATAPATH__0col_2__31_0__1_));
OR2X2 OR2X2_2586 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8285_), .B(AES_CORE_DATAPATH__abc_16009_new_n8286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8287_));
OR2X2 OR2X2_2587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5907_), .B(AES_CORE_DATAPATH__abc_16009_new_n8288_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8289_));
OR2X2 OR2X2_2588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8290_), .B(AES_CORE_DATAPATH__abc_16009_new_n8284_), .Y(AES_CORE_DATAPATH__0col_2__31_0__2_));
OR2X2 OR2X2_2589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8293_), .B(AES_CORE_DATAPATH__abc_16009_new_n8294_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8295_));
OR2X2 OR2X2_259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2927_), .B(AES_CORE_DATAPATH__abc_16009_new_n2928_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2929_));
OR2X2 OR2X2_2590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5957_), .B(AES_CORE_DATAPATH__abc_16009_new_n8296_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8297_));
OR2X2 OR2X2_2591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8298_), .B(AES_CORE_DATAPATH__abc_16009_new_n8292_), .Y(AES_CORE_DATAPATH__0col_2__31_0__3_));
OR2X2 OR2X2_2592 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8301_), .B(AES_CORE_DATAPATH__abc_16009_new_n8302_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8303_));
OR2X2 OR2X2_2593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6007_), .B(AES_CORE_DATAPATH__abc_16009_new_n8304_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8305_));
OR2X2 OR2X2_2594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8306_), .B(AES_CORE_DATAPATH__abc_16009_new_n8300_), .Y(AES_CORE_DATAPATH__0col_2__31_0__4_));
OR2X2 OR2X2_2595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8309_), .B(AES_CORE_DATAPATH__abc_16009_new_n8310_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8311_));
OR2X2 OR2X2_2596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6057_), .B(AES_CORE_DATAPATH__abc_16009_new_n8312_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8313_));
OR2X2 OR2X2_2597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8314_), .B(AES_CORE_DATAPATH__abc_16009_new_n8308_), .Y(AES_CORE_DATAPATH__0col_2__31_0__5_));
OR2X2 OR2X2_2598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8317_), .B(AES_CORE_DATAPATH__abc_16009_new_n8318_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8319_));
OR2X2 OR2X2_2599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6107_), .B(AES_CORE_DATAPATH__abc_16009_new_n8320_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8321_));
OR2X2 OR2X2_26 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n164_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n163_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_14_));
OR2X2 OR2X2_260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2929_), .B(AES_CORE_DATAPATH__abc_16009_new_n2926_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2930_));
OR2X2 OR2X2_2600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8322_), .B(AES_CORE_DATAPATH__abc_16009_new_n8316_), .Y(AES_CORE_DATAPATH__0col_2__31_0__6_));
OR2X2 OR2X2_2601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8325_), .B(AES_CORE_DATAPATH__abc_16009_new_n8326_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8327_));
OR2X2 OR2X2_2602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6157_), .B(AES_CORE_DATAPATH__abc_16009_new_n8328_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8329_));
OR2X2 OR2X2_2603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8330_), .B(AES_CORE_DATAPATH__abc_16009_new_n8324_), .Y(AES_CORE_DATAPATH__0col_2__31_0__7_));
OR2X2 OR2X2_2604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8333_), .B(AES_CORE_DATAPATH__abc_16009_new_n8334_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8335_));
OR2X2 OR2X2_2605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6207_), .B(AES_CORE_DATAPATH__abc_16009_new_n8336_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8337_));
OR2X2 OR2X2_2606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8338_), .B(AES_CORE_DATAPATH__abc_16009_new_n8332_), .Y(AES_CORE_DATAPATH__0col_2__31_0__8_));
OR2X2 OR2X2_2607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8341_), .B(AES_CORE_DATAPATH__abc_16009_new_n8342_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8343_));
OR2X2 OR2X2_2608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6257_), .B(AES_CORE_DATAPATH__abc_16009_new_n8344_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8345_));
OR2X2 OR2X2_2609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8346_), .B(AES_CORE_DATAPATH__abc_16009_new_n8340_), .Y(AES_CORE_DATAPATH__0col_2__31_0__9_));
OR2X2 OR2X2_261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2931_));
OR2X2 OR2X2_2610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8349_), .B(AES_CORE_DATAPATH__abc_16009_new_n8350_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8351_));
OR2X2 OR2X2_2611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6307_), .B(AES_CORE_DATAPATH__abc_16009_new_n8352_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8353_));
OR2X2 OR2X2_2612 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8354_), .B(AES_CORE_DATAPATH__abc_16009_new_n8348_), .Y(AES_CORE_DATAPATH__0col_2__31_0__10_));
OR2X2 OR2X2_2613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8357_), .B(AES_CORE_DATAPATH__abc_16009_new_n8358_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8359_));
OR2X2 OR2X2_2614 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6357_), .B(AES_CORE_DATAPATH__abc_16009_new_n8360_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8361_));
OR2X2 OR2X2_2615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8362_), .B(AES_CORE_DATAPATH__abc_16009_new_n8356_), .Y(AES_CORE_DATAPATH__0col_2__31_0__11_));
OR2X2 OR2X2_2616 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8365_), .B(AES_CORE_DATAPATH__abc_16009_new_n8366_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8367_));
OR2X2 OR2X2_2617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6407_), .B(AES_CORE_DATAPATH__abc_16009_new_n8368_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8369_));
OR2X2 OR2X2_2618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8370_), .B(AES_CORE_DATAPATH__abc_16009_new_n8364_), .Y(AES_CORE_DATAPATH__0col_2__31_0__12_));
OR2X2 OR2X2_2619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8373_), .B(AES_CORE_DATAPATH__abc_16009_new_n8374_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8375_));
OR2X2 OR2X2_262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2935_), .B(AES_CORE_DATAPATH__abc_16009_new_n2933_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2936_));
OR2X2 OR2X2_2620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6457_), .B(AES_CORE_DATAPATH__abc_16009_new_n8376_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8377_));
OR2X2 OR2X2_2621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8378_), .B(AES_CORE_DATAPATH__abc_16009_new_n8372_), .Y(AES_CORE_DATAPATH__0col_2__31_0__13_));
OR2X2 OR2X2_2622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8381_), .B(AES_CORE_DATAPATH__abc_16009_new_n8382_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8383_));
OR2X2 OR2X2_2623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6507_), .B(AES_CORE_DATAPATH__abc_16009_new_n8384_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8385_));
OR2X2 OR2X2_2624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8386_), .B(AES_CORE_DATAPATH__abc_16009_new_n8380_), .Y(AES_CORE_DATAPATH__0col_2__31_0__14_));
OR2X2 OR2X2_2625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8389_), .B(AES_CORE_DATAPATH__abc_16009_new_n8390_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8391_));
OR2X2 OR2X2_2626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6557_), .B(AES_CORE_DATAPATH__abc_16009_new_n8392_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8393_));
OR2X2 OR2X2_2627 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8394_), .B(AES_CORE_DATAPATH__abc_16009_new_n8388_), .Y(AES_CORE_DATAPATH__0col_2__31_0__15_));
OR2X2 OR2X2_2628 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8397_), .B(AES_CORE_DATAPATH__abc_16009_new_n8398_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8399_));
OR2X2 OR2X2_2629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6607_), .B(AES_CORE_DATAPATH__abc_16009_new_n8400_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8401_));
OR2X2 OR2X2_263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2936_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2937_));
OR2X2 OR2X2_2630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8402_), .B(AES_CORE_DATAPATH__abc_16009_new_n8396_), .Y(AES_CORE_DATAPATH__0col_2__31_0__16_));
OR2X2 OR2X2_2631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8405_), .B(AES_CORE_DATAPATH__abc_16009_new_n8406_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8407_));
OR2X2 OR2X2_2632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6657_), .B(AES_CORE_DATAPATH__abc_16009_new_n8408_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8409_));
OR2X2 OR2X2_2633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8410_), .B(AES_CORE_DATAPATH__abc_16009_new_n8404_), .Y(AES_CORE_DATAPATH__0col_2__31_0__17_));
OR2X2 OR2X2_2634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8413_), .B(AES_CORE_DATAPATH__abc_16009_new_n8414_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8415_));
OR2X2 OR2X2_2635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6707_), .B(AES_CORE_DATAPATH__abc_16009_new_n8416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8417_));
OR2X2 OR2X2_2636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8418_), .B(AES_CORE_DATAPATH__abc_16009_new_n8412_), .Y(AES_CORE_DATAPATH__0col_2__31_0__18_));
OR2X2 OR2X2_2637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8421_), .B(AES_CORE_DATAPATH__abc_16009_new_n8422_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8423_));
OR2X2 OR2X2_2638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6757_), .B(AES_CORE_DATAPATH__abc_16009_new_n8424_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8425_));
OR2X2 OR2X2_2639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8426_), .B(AES_CORE_DATAPATH__abc_16009_new_n8420_), .Y(AES_CORE_DATAPATH__0col_2__31_0__19_));
OR2X2 OR2X2_264 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2939_));
OR2X2 OR2X2_2640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8429_), .B(AES_CORE_DATAPATH__abc_16009_new_n8430_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8431_));
OR2X2 OR2X2_2641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6807_), .B(AES_CORE_DATAPATH__abc_16009_new_n8432_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8433_));
OR2X2 OR2X2_2642 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8434_), .B(AES_CORE_DATAPATH__abc_16009_new_n8428_), .Y(AES_CORE_DATAPATH__0col_2__31_0__20_));
OR2X2 OR2X2_2643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8437_), .B(AES_CORE_DATAPATH__abc_16009_new_n8438_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8439_));
OR2X2 OR2X2_2644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8440_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8441_));
OR2X2 OR2X2_2645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8442_), .B(AES_CORE_DATAPATH__abc_16009_new_n8436_), .Y(AES_CORE_DATAPATH__0col_2__31_0__21_));
OR2X2 OR2X2_2646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8445_), .B(AES_CORE_DATAPATH__abc_16009_new_n8446_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8447_));
OR2X2 OR2X2_2647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6907_), .B(AES_CORE_DATAPATH__abc_16009_new_n8448_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8449_));
OR2X2 OR2X2_2648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8450_), .B(AES_CORE_DATAPATH__abc_16009_new_n8444_), .Y(AES_CORE_DATAPATH__0col_2__31_0__22_));
OR2X2 OR2X2_2649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8453_), .B(AES_CORE_DATAPATH__abc_16009_new_n8454_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8455_));
OR2X2 OR2X2_265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2941_));
OR2X2 OR2X2_2650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6957_), .B(AES_CORE_DATAPATH__abc_16009_new_n8456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8457_));
OR2X2 OR2X2_2651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8458_), .B(AES_CORE_DATAPATH__abc_16009_new_n8452_), .Y(AES_CORE_DATAPATH__0col_2__31_0__23_));
OR2X2 OR2X2_2652 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8461_), .B(AES_CORE_DATAPATH__abc_16009_new_n8462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8463_));
OR2X2 OR2X2_2653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7007_), .B(AES_CORE_DATAPATH__abc_16009_new_n8464_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8465_));
OR2X2 OR2X2_2654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8466_), .B(AES_CORE_DATAPATH__abc_16009_new_n8460_), .Y(AES_CORE_DATAPATH__0col_2__31_0__24_));
OR2X2 OR2X2_2655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8469_), .B(AES_CORE_DATAPATH__abc_16009_new_n8470_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8471_));
OR2X2 OR2X2_2656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7057_), .B(AES_CORE_DATAPATH__abc_16009_new_n8472_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8473_));
OR2X2 OR2X2_2657 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8474_), .B(AES_CORE_DATAPATH__abc_16009_new_n8468_), .Y(AES_CORE_DATAPATH__0col_2__31_0__25_));
OR2X2 OR2X2_2658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8477_), .B(AES_CORE_DATAPATH__abc_16009_new_n8478_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8479_));
OR2X2 OR2X2_2659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7107_), .B(AES_CORE_DATAPATH__abc_16009_new_n8480_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8481_));
OR2X2 OR2X2_266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2942_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2943_));
OR2X2 OR2X2_2660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8482_), .B(AES_CORE_DATAPATH__abc_16009_new_n8476_), .Y(AES_CORE_DATAPATH__0col_2__31_0__26_));
OR2X2 OR2X2_2661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8485_), .B(AES_CORE_DATAPATH__abc_16009_new_n8486_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8487_));
OR2X2 OR2X2_2662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7157_), .B(AES_CORE_DATAPATH__abc_16009_new_n8488_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8489_));
OR2X2 OR2X2_2663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8490_), .B(AES_CORE_DATAPATH__abc_16009_new_n8484_), .Y(AES_CORE_DATAPATH__0col_2__31_0__27_));
OR2X2 OR2X2_2664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8493_), .B(AES_CORE_DATAPATH__abc_16009_new_n8494_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8495_));
OR2X2 OR2X2_2665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7207_), .B(AES_CORE_DATAPATH__abc_16009_new_n8496_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8497_));
OR2X2 OR2X2_2666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8498_), .B(AES_CORE_DATAPATH__abc_16009_new_n8492_), .Y(AES_CORE_DATAPATH__0col_2__31_0__28_));
OR2X2 OR2X2_2667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8501_), .B(AES_CORE_DATAPATH__abc_16009_new_n8502_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8503_));
OR2X2 OR2X2_2668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7257_), .B(AES_CORE_DATAPATH__abc_16009_new_n8504_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8505_));
OR2X2 OR2X2_2669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8506_), .B(AES_CORE_DATAPATH__abc_16009_new_n8500_), .Y(AES_CORE_DATAPATH__0col_2__31_0__29_));
OR2X2 OR2X2_267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2946_), .B(AES_CORE_DATAPATH__abc_16009_new_n2947_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2948_));
OR2X2 OR2X2_2670 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8509_), .B(AES_CORE_DATAPATH__abc_16009_new_n8510_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8511_));
OR2X2 OR2X2_2671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7307_), .B(AES_CORE_DATAPATH__abc_16009_new_n8512_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8513_));
OR2X2 OR2X2_2672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8514_), .B(AES_CORE_DATAPATH__abc_16009_new_n8508_), .Y(AES_CORE_DATAPATH__0col_2__31_0__30_));
OR2X2 OR2X2_2673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8517_), .B(AES_CORE_DATAPATH__abc_16009_new_n8518_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8519_));
OR2X2 OR2X2_2674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7357_), .B(AES_CORE_DATAPATH__abc_16009_new_n8520_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8521_));
OR2X2 OR2X2_2675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8522_), .B(AES_CORE_DATAPATH__abc_16009_new_n8516_), .Y(AES_CORE_DATAPATH__0col_2__31_0__31_));
OR2X2 OR2X2_2676 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5802_), .B(AES_CORE_DATAPATH__abc_16009_new_n5758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8524_));
OR2X2 OR2X2_2677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8526_), .B(AES_CORE_DATAPATH__abc_16009_new_n8529_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8530_));
OR2X2 OR2X2_2678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8533_), .B(AES_CORE_DATAPATH__abc_16009_new_n8532_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__0_));
OR2X2 OR2X2_2679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8536_), .B(AES_CORE_DATAPATH__abc_16009_new_n8535_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__1_));
OR2X2 OR2X2_268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2948_), .B(AES_CORE_DATAPATH__abc_16009_new_n2945_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2949_));
OR2X2 OR2X2_2680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8539_), .B(AES_CORE_DATAPATH__abc_16009_new_n8538_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__2_));
OR2X2 OR2X2_2681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8542_), .B(AES_CORE_DATAPATH__abc_16009_new_n8541_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__3_));
OR2X2 OR2X2_2682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8545_), .B(AES_CORE_DATAPATH__abc_16009_new_n8544_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__4_));
OR2X2 OR2X2_2683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8548_), .B(AES_CORE_DATAPATH__abc_16009_new_n8547_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__5_));
OR2X2 OR2X2_2684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8551_), .B(AES_CORE_DATAPATH__abc_16009_new_n8550_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__6_));
OR2X2 OR2X2_2685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8554_), .B(AES_CORE_DATAPATH__abc_16009_new_n8553_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__7_));
OR2X2 OR2X2_2686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8557_), .B(AES_CORE_DATAPATH__abc_16009_new_n8556_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__8_));
OR2X2 OR2X2_2687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8560_), .B(AES_CORE_DATAPATH__abc_16009_new_n8559_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__9_));
OR2X2 OR2X2_2688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8563_), .B(AES_CORE_DATAPATH__abc_16009_new_n8562_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__10_));
OR2X2 OR2X2_2689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8566_), .B(AES_CORE_DATAPATH__abc_16009_new_n8565_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__11_));
OR2X2 OR2X2_269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2953_), .B(AES_CORE_DATAPATH__abc_16009_new_n2951_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2954_));
OR2X2 OR2X2_2690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8569_), .B(AES_CORE_DATAPATH__abc_16009_new_n8568_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__12_));
OR2X2 OR2X2_2691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8572_), .B(AES_CORE_DATAPATH__abc_16009_new_n8571_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__13_));
OR2X2 OR2X2_2692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8575_), .B(AES_CORE_DATAPATH__abc_16009_new_n8574_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__14_));
OR2X2 OR2X2_2693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8578_), .B(AES_CORE_DATAPATH__abc_16009_new_n8577_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__15_));
OR2X2 OR2X2_2694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8581_), .B(AES_CORE_DATAPATH__abc_16009_new_n8580_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__16_));
OR2X2 OR2X2_2695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8584_), .B(AES_CORE_DATAPATH__abc_16009_new_n8583_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__17_));
OR2X2 OR2X2_2696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8587_), .B(AES_CORE_DATAPATH__abc_16009_new_n8586_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__18_));
OR2X2 OR2X2_2697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8590_), .B(AES_CORE_DATAPATH__abc_16009_new_n8589_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__19_));
OR2X2 OR2X2_2698 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8593_), .B(AES_CORE_DATAPATH__abc_16009_new_n8592_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__20_));
OR2X2 OR2X2_2699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8596_), .B(AES_CORE_DATAPATH__abc_16009_new_n8595_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__21_));
OR2X2 OR2X2_27 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT_state_13_), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_2_));
OR2X2 OR2X2_270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2954_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2955_));
OR2X2 OR2X2_2700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8599_), .B(AES_CORE_DATAPATH__abc_16009_new_n8598_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__22_));
OR2X2 OR2X2_2701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8602_), .B(AES_CORE_DATAPATH__abc_16009_new_n8601_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__23_));
OR2X2 OR2X2_2702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8605_), .B(AES_CORE_DATAPATH__abc_16009_new_n8604_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__24_));
OR2X2 OR2X2_2703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8608_), .B(AES_CORE_DATAPATH__abc_16009_new_n8607_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__25_));
OR2X2 OR2X2_2704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8611_), .B(AES_CORE_DATAPATH__abc_16009_new_n8610_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__26_));
OR2X2 OR2X2_2705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8614_), .B(AES_CORE_DATAPATH__abc_16009_new_n8613_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__27_));
OR2X2 OR2X2_2706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8617_), .B(AES_CORE_DATAPATH__abc_16009_new_n8616_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__28_));
OR2X2 OR2X2_2707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8620_), .B(AES_CORE_DATAPATH__abc_16009_new_n8619_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__29_));
OR2X2 OR2X2_2708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8623_), .B(AES_CORE_DATAPATH__abc_16009_new_n8622_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__30_));
OR2X2 OR2X2_2709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8626_), .B(AES_CORE_DATAPATH__abc_16009_new_n8625_), .Y(AES_CORE_DATAPATH__0bkp_1_3__31_0__31_));
OR2X2 OR2X2_271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2957_));
OR2X2 OR2X2_2710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5808_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8629_));
OR2X2 OR2X2_2711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8630_));
OR2X2 OR2X2_2712 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8634_));
OR2X2 OR2X2_2713 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8632_), .B(AES_CORE_DATAPATH__abc_16009_new_n8634_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8635_));
OR2X2 OR2X2_2714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8636_));
OR2X2 OR2X2_2715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5858_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8638_));
OR2X2 OR2X2_2716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8639_));
OR2X2 OR2X2_2717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8643_));
OR2X2 OR2X2_2718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8641_), .B(AES_CORE_DATAPATH__abc_16009_new_n8643_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8644_));
OR2X2 OR2X2_2719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8645_));
OR2X2 OR2X2_272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2959_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2960_));
OR2X2 OR2X2_2720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5908_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8647_));
OR2X2 OR2X2_2721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8648_));
OR2X2 OR2X2_2722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8651_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8652_));
OR2X2 OR2X2_2723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8650_), .B(AES_CORE_DATAPATH__abc_16009_new_n8652_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8653_));
OR2X2 OR2X2_2724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8654_));
OR2X2 OR2X2_2725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n5958_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8656_));
OR2X2 OR2X2_2726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8657_));
OR2X2 OR2X2_2727 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8660_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8661_));
OR2X2 OR2X2_2728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8659_), .B(AES_CORE_DATAPATH__abc_16009_new_n8661_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8662_));
OR2X2 OR2X2_2729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8663_));
OR2X2 OR2X2_273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2963_), .B(AES_CORE_DATAPATH__abc_16009_new_n2964_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2965_));
OR2X2 OR2X2_2730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6008_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8665_));
OR2X2 OR2X2_2731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8666_));
OR2X2 OR2X2_2732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8669_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8670_));
OR2X2 OR2X2_2733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8668_), .B(AES_CORE_DATAPATH__abc_16009_new_n8670_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8671_));
OR2X2 OR2X2_2734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8672_));
OR2X2 OR2X2_2735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6058_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8674_));
OR2X2 OR2X2_2736 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8675_));
OR2X2 OR2X2_2737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8678_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8679_));
OR2X2 OR2X2_2738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8677_), .B(AES_CORE_DATAPATH__abc_16009_new_n8679_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8680_));
OR2X2 OR2X2_2739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8681_));
OR2X2 OR2X2_274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2965_), .B(AES_CORE_DATAPATH__abc_16009_new_n2962_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2966_));
OR2X2 OR2X2_2740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6108_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8683_));
OR2X2 OR2X2_2741 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8684_));
OR2X2 OR2X2_2742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8688_));
OR2X2 OR2X2_2743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8686_), .B(AES_CORE_DATAPATH__abc_16009_new_n8688_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8689_));
OR2X2 OR2X2_2744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8690_));
OR2X2 OR2X2_2745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6158_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8692_));
OR2X2 OR2X2_2746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8693_));
OR2X2 OR2X2_2747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8696_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8697_));
OR2X2 OR2X2_2748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8695_), .B(AES_CORE_DATAPATH__abc_16009_new_n8697_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8698_));
OR2X2 OR2X2_2749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8699_));
OR2X2 OR2X2_275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2967_));
OR2X2 OR2X2_2750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6208_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8701_));
OR2X2 OR2X2_2751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8702_));
OR2X2 OR2X2_2752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8705_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8706_));
OR2X2 OR2X2_2753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8704_), .B(AES_CORE_DATAPATH__abc_16009_new_n8706_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8707_));
OR2X2 OR2X2_2754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8708_));
OR2X2 OR2X2_2755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6258_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8710_));
OR2X2 OR2X2_2756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8711_));
OR2X2 OR2X2_2757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8714_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8715_));
OR2X2 OR2X2_2758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8713_), .B(AES_CORE_DATAPATH__abc_16009_new_n8715_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8716_));
OR2X2 OR2X2_2759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8717_));
OR2X2 OR2X2_276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2971_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2972_));
OR2X2 OR2X2_2760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6308_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8719_));
OR2X2 OR2X2_2761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8720_));
OR2X2 OR2X2_2762 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8723_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8724_));
OR2X2 OR2X2_2763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8722_), .B(AES_CORE_DATAPATH__abc_16009_new_n8724_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8725_));
OR2X2 OR2X2_2764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8726_));
OR2X2 OR2X2_2765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6358_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8728_));
OR2X2 OR2X2_2766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8729_));
OR2X2 OR2X2_2767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8732_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8733_));
OR2X2 OR2X2_2768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8731_), .B(AES_CORE_DATAPATH__abc_16009_new_n8733_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8734_));
OR2X2 OR2X2_2769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8735_));
OR2X2 OR2X2_277 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2972_), .B(AES_CORE_DATAPATH__abc_16009_new_n2969_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2973_));
OR2X2 OR2X2_2770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6408_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8737_));
OR2X2 OR2X2_2771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8738_));
OR2X2 OR2X2_2772 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8741_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8742_));
OR2X2 OR2X2_2773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8740_), .B(AES_CORE_DATAPATH__abc_16009_new_n8742_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8743_));
OR2X2 OR2X2_2774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8744_));
OR2X2 OR2X2_2775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6458_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8746_));
OR2X2 OR2X2_2776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8747_));
OR2X2 OR2X2_2777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8750_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8751_));
OR2X2 OR2X2_2778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8749_), .B(AES_CORE_DATAPATH__abc_16009_new_n8751_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8752_));
OR2X2 OR2X2_2779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8753_));
OR2X2 OR2X2_278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2977_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2978_));
OR2X2 OR2X2_2780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6508_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8755_));
OR2X2 OR2X2_2781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8756_));
OR2X2 OR2X2_2782 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8760_));
OR2X2 OR2X2_2783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8758_), .B(AES_CORE_DATAPATH__abc_16009_new_n8760_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8761_));
OR2X2 OR2X2_2784 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8762_));
OR2X2 OR2X2_2785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6558_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8764_));
OR2X2 OR2X2_2786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8765_));
OR2X2 OR2X2_2787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8768_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8769_));
OR2X2 OR2X2_2788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8767_), .B(AES_CORE_DATAPATH__abc_16009_new_n8769_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8770_));
OR2X2 OR2X2_2789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8771_));
OR2X2 OR2X2_279 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2981_), .B(AES_CORE_DATAPATH__abc_16009_new_n2982_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2983_));
OR2X2 OR2X2_2790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6608_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8773_));
OR2X2 OR2X2_2791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8774_));
OR2X2 OR2X2_2792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8778_));
OR2X2 OR2X2_2793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8776_), .B(AES_CORE_DATAPATH__abc_16009_new_n8778_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8779_));
OR2X2 OR2X2_2794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8780_));
OR2X2 OR2X2_2795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6658_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8782_));
OR2X2 OR2X2_2796 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8783_));
OR2X2 OR2X2_2797 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8786_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8787_));
OR2X2 OR2X2_2798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8785_), .B(AES_CORE_DATAPATH__abc_16009_new_n8787_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8788_));
OR2X2 OR2X2_2799 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8789_));
OR2X2 OR2X2_28 ( .A(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .B(AES_CORE_CONTROL_UNIT_rd_count_0_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n172_));
OR2X2 OR2X2_280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2983_), .B(AES_CORE_DATAPATH__abc_16009_new_n2980_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2984_));
OR2X2 OR2X2_2800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6708_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8791_));
OR2X2 OR2X2_2801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8792_));
OR2X2 OR2X2_2802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8795_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8796_));
OR2X2 OR2X2_2803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8794_), .B(AES_CORE_DATAPATH__abc_16009_new_n8796_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8797_));
OR2X2 OR2X2_2804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8798_));
OR2X2 OR2X2_2805 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6758_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8800_));
OR2X2 OR2X2_2806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8801_));
OR2X2 OR2X2_2807 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8804_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8805_));
OR2X2 OR2X2_2808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8803_), .B(AES_CORE_DATAPATH__abc_16009_new_n8805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8806_));
OR2X2 OR2X2_2809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8807_));
OR2X2 OR2X2_281 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2985_));
OR2X2 OR2X2_2810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6808_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8809_));
OR2X2 OR2X2_2811 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8810_));
OR2X2 OR2X2_2812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8814_));
OR2X2 OR2X2_2813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8812_), .B(AES_CORE_DATAPATH__abc_16009_new_n8814_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8815_));
OR2X2 OR2X2_2814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8816_));
OR2X2 OR2X2_2815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6858_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8818_));
OR2X2 OR2X2_2816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8819_));
OR2X2 OR2X2_2817 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8823_));
OR2X2 OR2X2_2818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8821_), .B(AES_CORE_DATAPATH__abc_16009_new_n8823_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8824_));
OR2X2 OR2X2_2819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8825_));
OR2X2 OR2X2_282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2987_), .B(AES_CORE_DATAPATH__abc_16009_new_n2976_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2988_));
OR2X2 OR2X2_2820 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6908_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8827_));
OR2X2 OR2X2_2821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8828_));
OR2X2 OR2X2_2822 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8832_));
OR2X2 OR2X2_2823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8830_), .B(AES_CORE_DATAPATH__abc_16009_new_n8832_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8833_));
OR2X2 OR2X2_2824 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8834_));
OR2X2 OR2X2_2825 ( .A(AES_CORE_DATAPATH__abc_16009_new_n6958_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8836_));
OR2X2 OR2X2_2826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8837_));
OR2X2 OR2X2_2827 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8840_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8841_));
OR2X2 OR2X2_2828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8839_), .B(AES_CORE_DATAPATH__abc_16009_new_n8841_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8842_));
OR2X2 OR2X2_2829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8843_));
OR2X2 OR2X2_283 ( .A(\key_out[8] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2989_));
OR2X2 OR2X2_2830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7008_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8845_));
OR2X2 OR2X2_2831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8846_));
OR2X2 OR2X2_2832 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8849_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8850_));
OR2X2 OR2X2_2833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8848_), .B(AES_CORE_DATAPATH__abc_16009_new_n8850_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8851_));
OR2X2 OR2X2_2834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8852_));
OR2X2 OR2X2_2835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7058_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8854_));
OR2X2 OR2X2_2836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8855_));
OR2X2 OR2X2_2837 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8858_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8859_));
OR2X2 OR2X2_2838 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8859_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8860_));
OR2X2 OR2X2_2839 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8861_));
OR2X2 OR2X2_284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2991_), .B(AES_CORE_DATAPATH__abc_16009_new_n2975_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__8_));
OR2X2 OR2X2_2840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7108_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8863_));
OR2X2 OR2X2_2841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8864_));
OR2X2 OR2X2_2842 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8868_));
OR2X2 OR2X2_2843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8866_), .B(AES_CORE_DATAPATH__abc_16009_new_n8868_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8869_));
OR2X2 OR2X2_2844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8870_));
OR2X2 OR2X2_2845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7158_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8872_));
OR2X2 OR2X2_2846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8873_));
OR2X2 OR2X2_2847 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8876_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8877_));
OR2X2 OR2X2_2848 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8875_), .B(AES_CORE_DATAPATH__abc_16009_new_n8877_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8878_));
OR2X2 OR2X2_2849 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8879_));
OR2X2 OR2X2_285 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2993_));
OR2X2 OR2X2_2850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7208_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8881_));
OR2X2 OR2X2_2851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8882_));
OR2X2 OR2X2_2852 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8885_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8886_));
OR2X2 OR2X2_2853 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8884_), .B(AES_CORE_DATAPATH__abc_16009_new_n8886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8887_));
OR2X2 OR2X2_2854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8888_));
OR2X2 OR2X2_2855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7258_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8890_));
OR2X2 OR2X2_2856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8891_));
OR2X2 OR2X2_2857 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8894_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8895_));
OR2X2 OR2X2_2858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8893_), .B(AES_CORE_DATAPATH__abc_16009_new_n8895_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8896_));
OR2X2 OR2X2_2859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8897_));
OR2X2 OR2X2_286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n2995_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2996_));
OR2X2 OR2X2_2860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7308_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8899_));
OR2X2 OR2X2_2861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8900_));
OR2X2 OR2X2_2862 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8903_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8904_));
OR2X2 OR2X2_2863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8902_), .B(AES_CORE_DATAPATH__abc_16009_new_n8904_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8905_));
OR2X2 OR2X2_2864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8906_));
OR2X2 OR2X2_2865 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7358_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8908_));
OR2X2 OR2X2_2866 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8909_));
OR2X2 OR2X2_2867 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8531_), .B(AES_CORE_DATAPATH__abc_16009_new_n8912_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8913_));
OR2X2 OR2X2_2868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8911_), .B(AES_CORE_DATAPATH__abc_16009_new_n8913_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8914_));
OR2X2 OR2X2_2869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8530_), .B(AES_CORE_DATAPATH_bkp_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8915_));
OR2X2 OR2X2_287 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2999_), .B(AES_CORE_DATAPATH__abc_16009_new_n3000_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3001_));
OR2X2 OR2X2_2870 ( .A(AES_CORE_CONTROL_UNIT_iv_cnt_en), .B(\iv_en[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n8917_));
OR2X2 OR2X2_2871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n8919_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8920_));
OR2X2 OR2X2_2872 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8921_), .B(AES_CORE_DATAPATH_iv_3__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8922_));
OR2X2 OR2X2_2873 ( .A(\bus_in[0] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8923_));
OR2X2 OR2X2_2874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8927_), .B(AES_CORE_DATAPATH__abc_16009_new_n8918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8928_));
OR2X2 OR2X2_2875 ( .A(\bus_in[1] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8930_));
OR2X2 OR2X2_2876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8935_), .B(AES_CORE_DATAPATH__abc_16009_new_n8918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8936_));
OR2X2 OR2X2_2877 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8938_), .B(AES_CORE_DATAPATH__abc_16009_new_n8937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8939_));
OR2X2 OR2X2_2878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8940_), .B(AES_CORE_DATAPATH_iv_3__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8941_));
OR2X2 OR2X2_2879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8932_), .B(AES_CORE_DATAPATH__abc_16009_new_n8937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8943_));
OR2X2 OR2X2_288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3001_), .B(AES_CORE_DATAPATH__abc_16009_new_n2998_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3002_));
OR2X2 OR2X2_2880 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8944_), .B(AES_CORE_DATAPATH_iv_3__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8945_));
OR2X2 OR2X2_2881 ( .A(\bus_in[2] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8946_));
OR2X2 OR2X2_2882 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8950_), .B(AES_CORE_DATAPATH__abc_16009_new_n8918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8951_));
OR2X2 OR2X2_2883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8947_), .B(AES_CORE_DATAPATH__abc_16009_new_n8937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8953_));
OR2X2 OR2X2_2884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8954_), .B(AES_CORE_DATAPATH_iv_3__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8955_));
OR2X2 OR2X2_2885 ( .A(\bus_in[3] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8956_));
OR2X2 OR2X2_2886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8962_), .B(AES_CORE_DATAPATH__abc_16009_new_n8918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8963_));
OR2X2 OR2X2_2887 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8959_), .B(AES_CORE_DATAPATH__abc_16009_new_n8937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8965_));
OR2X2 OR2X2_2888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8966_), .B(AES_CORE_DATAPATH_iv_3__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8967_));
OR2X2 OR2X2_2889 ( .A(\bus_in[4] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8968_));
OR2X2 OR2X2_289 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3003_));
OR2X2 OR2X2_2890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8972_), .B(AES_CORE_DATAPATH__abc_16009_new_n8918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8973_));
OR2X2 OR2X2_2891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8969_), .B(AES_CORE_DATAPATH_iv_3__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8976_));
OR2X2 OR2X2_2892 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8980_), .B(AES_CORE_DATAPATH__abc_16009_new_n8937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8981_));
OR2X2 OR2X2_2893 ( .A(\bus_in[5] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8982_));
OR2X2 OR2X2_2894 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8984_), .B(AES_CORE_DATAPATH__abc_16009_new_n8975_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__5_));
OR2X2 OR2X2_2895 ( .A(\bus_in[6] ), .B(AES_CORE_CONTROL_UNIT_iv_cnt_en), .Y(AES_CORE_DATAPATH__abc_16009_new_n8987_));
OR2X2 OR2X2_2896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8989_), .B(AES_CORE_DATAPATH__abc_16009_new_n8991_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8992_));
OR2X2 OR2X2_2897 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8992_), .B(AES_CORE_DATAPATH__abc_16009_new_n8937_), .Y(AES_CORE_DATAPATH__abc_16009_new_n8993_));
OR2X2 OR2X2_2898 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8994_), .B(AES_CORE_DATAPATH__abc_16009_new_n8986_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__6_));
OR2X2 OR2X2_2899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9002_), .B(AES_CORE_DATAPATH__abc_16009_new_n8996_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9003_));
OR2X2 OR2X2_29 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n173_), .B(AES_CORE_CONTROL_UNIT_rd_count_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n177_));
OR2X2 OR2X2_290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3007_), .B(AES_CORE_DATAPATH__abc_16009_new_n3005_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3008_));
OR2X2 OR2X2_2900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9001_), .B(AES_CORE_DATAPATH__abc_16009_new_n8920_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9005_));
OR2X2 OR2X2_2901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9004_), .B(AES_CORE_DATAPATH__abc_16009_new_n9006_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__7_));
OR2X2 OR2X2_2902 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9012_), .B(AES_CORE_DATAPATH__abc_16009_new_n9008_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9013_));
OR2X2 OR2X2_2903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9011_), .B(AES_CORE_DATAPATH__abc_16009_new_n8920_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9015_));
OR2X2 OR2X2_2904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9014_), .B(AES_CORE_DATAPATH__abc_16009_new_n9016_), .Y(AES_CORE_DATAPATH__0iv_3__31_0__8_));
OR2X2 OR2X2_2905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9018_));
OR2X2 OR2X2_2906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9009_), .B(AES_CORE_DATAPATH_iv_3__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9019_));
OR2X2 OR2X2_2907 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9024_), .B(AES_CORE_DATAPATH__abc_16009_new_n9020_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9025_));
OR2X2 OR2X2_2908 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9027_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9028_));
OR2X2 OR2X2_2909 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9026_), .B(AES_CORE_DATAPATH__abc_16009_new_n9028_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9029_));
OR2X2 OR2X2_291 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3008_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3009_));
OR2X2 OR2X2_2910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9031_));
OR2X2 OR2X2_2911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9022_), .B(AES_CORE_DATAPATH_iv_3__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9032_));
OR2X2 OR2X2_2912 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9037_), .B(AES_CORE_DATAPATH__abc_16009_new_n9038_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9039_));
OR2X2 OR2X2_2913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9039_), .B(AES_CORE_DATAPATH__abc_16009_new_n8918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9040_));
OR2X2 OR2X2_2914 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9036_), .B(AES_CORE_DATAPATH__abc_16009_new_n9040_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9041_));
OR2X2 OR2X2_2915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9043_));
OR2X2 OR2X2_2916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9033_), .B(AES_CORE_DATAPATH_iv_3__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9044_));
OR2X2 OR2X2_2917 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9048_), .B(AES_CORE_DATAPATH__abc_16009_new_n9045_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9049_));
OR2X2 OR2X2_2918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9051_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9052_));
OR2X2 OR2X2_2919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9050_), .B(AES_CORE_DATAPATH__abc_16009_new_n9052_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9053_));
OR2X2 OR2X2_292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3013_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3014_));
OR2X2 OR2X2_2920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9055_));
OR2X2 OR2X2_2921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9046_), .B(AES_CORE_DATAPATH_iv_3__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9058_));
OR2X2 OR2X2_2922 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9062_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9063_));
OR2X2 OR2X2_2923 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9063_), .B(AES_CORE_DATAPATH__abc_16009_new_n9061_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9064_));
OR2X2 OR2X2_2924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9060_), .B(AES_CORE_DATAPATH__abc_16009_new_n9064_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9065_));
OR2X2 OR2X2_2925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9067_));
OR2X2 OR2X2_2926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9056_), .B(AES_CORE_DATAPATH_iv_3__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9070_));
OR2X2 OR2X2_2927 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9074_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9075_));
OR2X2 OR2X2_2928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9075_), .B(AES_CORE_DATAPATH__abc_16009_new_n9073_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9076_));
OR2X2 OR2X2_2929 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9072_), .B(AES_CORE_DATAPATH__abc_16009_new_n9076_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9077_));
OR2X2 OR2X2_293 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3017_), .B(AES_CORE_DATAPATH__abc_16009_new_n3018_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3019_));
OR2X2 OR2X2_2930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9079_));
OR2X2 OR2X2_2931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9068_), .B(AES_CORE_DATAPATH_iv_3__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9082_));
OR2X2 OR2X2_2932 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9087_));
OR2X2 OR2X2_2933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9087_), .B(AES_CORE_DATAPATH__abc_16009_new_n9085_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9088_));
OR2X2 OR2X2_2934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9084_), .B(AES_CORE_DATAPATH__abc_16009_new_n9088_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9089_));
OR2X2 OR2X2_2935 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9091_));
OR2X2 OR2X2_2936 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9080_), .B(AES_CORE_DATAPATH_iv_3__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9094_));
OR2X2 OR2X2_2937 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9098_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9099_));
OR2X2 OR2X2_2938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9099_), .B(AES_CORE_DATAPATH__abc_16009_new_n9097_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9100_));
OR2X2 OR2X2_2939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9096_), .B(AES_CORE_DATAPATH__abc_16009_new_n9100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9101_));
OR2X2 OR2X2_294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3019_), .B(AES_CORE_DATAPATH__abc_16009_new_n3016_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3020_));
OR2X2 OR2X2_2940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9103_));
OR2X2 OR2X2_2941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9092_), .B(AES_CORE_DATAPATH_iv_3__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9106_));
OR2X2 OR2X2_2942 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9111_));
OR2X2 OR2X2_2943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9111_), .B(AES_CORE_DATAPATH__abc_16009_new_n9109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9112_));
OR2X2 OR2X2_2944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9108_), .B(AES_CORE_DATAPATH__abc_16009_new_n9112_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9113_));
OR2X2 OR2X2_2945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9115_));
OR2X2 OR2X2_2946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9104_), .B(AES_CORE_DATAPATH_iv_3__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9118_));
OR2X2 OR2X2_2947 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9123_));
OR2X2 OR2X2_2948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9123_), .B(AES_CORE_DATAPATH__abc_16009_new_n9121_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9124_));
OR2X2 OR2X2_2949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9120_), .B(AES_CORE_DATAPATH__abc_16009_new_n9124_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9125_));
OR2X2 OR2X2_295 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3021_));
OR2X2 OR2X2_2950 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9127_));
OR2X2 OR2X2_2951 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9116_), .B(AES_CORE_DATAPATH_iv_3__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9128_));
OR2X2 OR2X2_2952 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9135_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9136_));
OR2X2 OR2X2_2953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9136_), .B(AES_CORE_DATAPATH__abc_16009_new_n9134_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9137_));
OR2X2 OR2X2_2954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9133_), .B(AES_CORE_DATAPATH__abc_16009_new_n9137_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9138_));
OR2X2 OR2X2_2955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9140_));
OR2X2 OR2X2_2956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9130_), .B(AES_CORE_DATAPATH_iv_3__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9143_));
OR2X2 OR2X2_2957 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9147_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9148_));
OR2X2 OR2X2_2958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9148_), .B(AES_CORE_DATAPATH__abc_16009_new_n9146_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9149_));
OR2X2 OR2X2_2959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9145_), .B(AES_CORE_DATAPATH__abc_16009_new_n9149_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9150_));
OR2X2 OR2X2_296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3023_), .B(AES_CORE_DATAPATH__abc_16009_new_n3012_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3024_));
OR2X2 OR2X2_2960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9152_));
OR2X2 OR2X2_2961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9154_), .B(AES_CORE_DATAPATH_iv_3__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9155_));
OR2X2 OR2X2_2962 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9161_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9162_));
OR2X2 OR2X2_2963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9162_), .B(AES_CORE_DATAPATH__abc_16009_new_n9160_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9163_));
OR2X2 OR2X2_2964 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9159_), .B(AES_CORE_DATAPATH__abc_16009_new_n9163_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9164_));
OR2X2 OR2X2_2965 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9166_));
OR2X2 OR2X2_2966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9167_), .B(AES_CORE_DATAPATH__abc_16009_new_n9169_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9170_));
OR2X2 OR2X2_2967 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9173_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9174_));
OR2X2 OR2X2_2968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9174_), .B(AES_CORE_DATAPATH__abc_16009_new_n9172_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9175_));
OR2X2 OR2X2_2969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9171_), .B(AES_CORE_DATAPATH__abc_16009_new_n9175_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9176_));
OR2X2 OR2X2_297 ( .A(\key_out[10] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3025_));
OR2X2 OR2X2_2970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9178_));
OR2X2 OR2X2_2971 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9179_), .B(AES_CORE_DATAPATH_iv_3__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9180_));
OR2X2 OR2X2_2972 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9188_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9189_));
OR2X2 OR2X2_2973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9189_), .B(AES_CORE_DATAPATH__abc_16009_new_n9187_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9190_));
OR2X2 OR2X2_2974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9186_), .B(AES_CORE_DATAPATH__abc_16009_new_n9190_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9191_));
OR2X2 OR2X2_2975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9193_));
OR2X2 OR2X2_2976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9183_), .B(AES_CORE_DATAPATH_iv_3__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9196_));
OR2X2 OR2X2_2977 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9200_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9201_));
OR2X2 OR2X2_2978 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9201_), .B(AES_CORE_DATAPATH__abc_16009_new_n9199_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9202_));
OR2X2 OR2X2_2979 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9198_), .B(AES_CORE_DATAPATH__abc_16009_new_n9202_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9203_));
OR2X2 OR2X2_298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3027_), .B(AES_CORE_DATAPATH__abc_16009_new_n3011_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__10_));
OR2X2 OR2X2_2980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9205_));
OR2X2 OR2X2_2981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9207_), .B(AES_CORE_DATAPATH_iv_3__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9208_));
OR2X2 OR2X2_2982 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9214_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9215_));
OR2X2 OR2X2_2983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9215_), .B(AES_CORE_DATAPATH__abc_16009_new_n9213_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9216_));
OR2X2 OR2X2_2984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9212_), .B(AES_CORE_DATAPATH__abc_16009_new_n9216_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9217_));
OR2X2 OR2X2_2985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9219_));
OR2X2 OR2X2_2986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9220_), .B(AES_CORE_DATAPATH__abc_16009_new_n9222_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9223_));
OR2X2 OR2X2_2987 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9226_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9227_));
OR2X2 OR2X2_2988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9227_), .B(AES_CORE_DATAPATH__abc_16009_new_n9225_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9228_));
OR2X2 OR2X2_2989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9224_), .B(AES_CORE_DATAPATH__abc_16009_new_n9228_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9229_));
OR2X2 OR2X2_299 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3029_));
OR2X2 OR2X2_2990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9231_));
OR2X2 OR2X2_2991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9232_), .B(AES_CORE_DATAPATH_iv_3__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9233_));
OR2X2 OR2X2_2992 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9239_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9240_));
OR2X2 OR2X2_2993 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9240_), .B(AES_CORE_DATAPATH__abc_16009_new_n9238_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9241_));
OR2X2 OR2X2_2994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9237_), .B(AES_CORE_DATAPATH__abc_16009_new_n9241_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9242_));
OR2X2 OR2X2_2995 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9244_));
OR2X2 OR2X2_2996 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9234_), .B(AES_CORE_DATAPATH_iv_3__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9245_));
OR2X2 OR2X2_2997 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9251_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9252_));
OR2X2 OR2X2_2998 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9252_), .B(AES_CORE_DATAPATH__abc_16009_new_n9250_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9253_));
OR2X2 OR2X2_2999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9249_), .B(AES_CORE_DATAPATH__abc_16009_new_n9253_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9254_));
OR2X2 OR2X2_3 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n96_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n91_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n97_));
OR2X2 OR2X2_30 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n178_), .B(AES_CORE_CONTROL_UNIT_rd_count_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n184_));
OR2X2 OR2X2_300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3031_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3032_));
OR2X2 OR2X2_3000 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9256_));
OR2X2 OR2X2_3001 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9246_), .B(AES_CORE_DATAPATH_iv_3__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9257_));
OR2X2 OR2X2_3002 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9263_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9264_));
OR2X2 OR2X2_3003 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9264_), .B(AES_CORE_DATAPATH__abc_16009_new_n9262_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9265_));
OR2X2 OR2X2_3004 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9261_), .B(AES_CORE_DATAPATH__abc_16009_new_n9265_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9266_));
OR2X2 OR2X2_3005 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9268_));
OR2X2 OR2X2_3006 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9258_), .B(AES_CORE_DATAPATH_iv_3__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9269_));
OR2X2 OR2X2_3007 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9275_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9276_));
OR2X2 OR2X2_3008 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9276_), .B(AES_CORE_DATAPATH__abc_16009_new_n9274_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9277_));
OR2X2 OR2X2_3009 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9273_), .B(AES_CORE_DATAPATH__abc_16009_new_n9277_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9278_));
OR2X2 OR2X2_301 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3035_), .B(AES_CORE_DATAPATH__abc_16009_new_n3036_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3037_));
OR2X2 OR2X2_3010 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9280_));
OR2X2 OR2X2_3011 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9270_), .B(AES_CORE_DATAPATH_iv_3__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9283_));
OR2X2 OR2X2_3012 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9287_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9288_));
OR2X2 OR2X2_3013 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9288_), .B(AES_CORE_DATAPATH__abc_16009_new_n9286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9289_));
OR2X2 OR2X2_3014 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9285_), .B(AES_CORE_DATAPATH__abc_16009_new_n9289_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9290_));
OR2X2 OR2X2_3015 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8917_), .B(AES_CORE_DATAPATH_iv_3__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9292_));
OR2X2 OR2X2_3016 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9293_), .B(AES_CORE_DATAPATH__abc_16009_new_n9295_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9296_));
OR2X2 OR2X2_3017 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8918_), .B(AES_CORE_DATAPATH__abc_16009_new_n9299_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9300_));
OR2X2 OR2X2_3018 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9300_), .B(AES_CORE_DATAPATH__abc_16009_new_n9298_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9301_));
OR2X2 OR2X2_3019 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9297_), .B(AES_CORE_DATAPATH__abc_16009_new_n9301_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9302_));
OR2X2 OR2X2_302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3037_), .B(AES_CORE_DATAPATH__abc_16009_new_n3034_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3038_));
OR2X2 OR2X2_3020 ( .A(AES_CORE_DATAPATH_iv_2__0_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9304_));
OR2X2 OR2X2_3021 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9306_));
OR2X2 OR2X2_3022 ( .A(AES_CORE_DATAPATH_iv_2__1_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9308_));
OR2X2 OR2X2_3023 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9309_));
OR2X2 OR2X2_3024 ( .A(AES_CORE_DATAPATH_iv_2__2_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9311_));
OR2X2 OR2X2_3025 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9312_));
OR2X2 OR2X2_3026 ( .A(AES_CORE_DATAPATH_iv_2__3_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9314_));
OR2X2 OR2X2_3027 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9315_));
OR2X2 OR2X2_3028 ( .A(AES_CORE_DATAPATH_iv_2__4_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9317_));
OR2X2 OR2X2_3029 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9318_));
OR2X2 OR2X2_303 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3039_));
OR2X2 OR2X2_3030 ( .A(AES_CORE_DATAPATH_iv_2__5_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9320_));
OR2X2 OR2X2_3031 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9321_));
OR2X2 OR2X2_3032 ( .A(AES_CORE_DATAPATH_iv_2__6_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9323_));
OR2X2 OR2X2_3033 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9324_));
OR2X2 OR2X2_3034 ( .A(AES_CORE_DATAPATH_iv_2__7_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9326_));
OR2X2 OR2X2_3035 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9327_));
OR2X2 OR2X2_3036 ( .A(AES_CORE_DATAPATH_iv_2__8_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9329_));
OR2X2 OR2X2_3037 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9330_));
OR2X2 OR2X2_3038 ( .A(AES_CORE_DATAPATH_iv_2__9_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9332_));
OR2X2 OR2X2_3039 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9333_));
OR2X2 OR2X2_304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3043_), .B(AES_CORE_DATAPATH__abc_16009_new_n3041_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3044_));
OR2X2 OR2X2_3040 ( .A(AES_CORE_DATAPATH_iv_2__10_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9335_));
OR2X2 OR2X2_3041 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9336_));
OR2X2 OR2X2_3042 ( .A(AES_CORE_DATAPATH_iv_2__11_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9338_));
OR2X2 OR2X2_3043 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9339_));
OR2X2 OR2X2_3044 ( .A(AES_CORE_DATAPATH_iv_2__12_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9341_));
OR2X2 OR2X2_3045 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9342_));
OR2X2 OR2X2_3046 ( .A(AES_CORE_DATAPATH_iv_2__13_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9344_));
OR2X2 OR2X2_3047 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9345_));
OR2X2 OR2X2_3048 ( .A(AES_CORE_DATAPATH_iv_2__14_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9347_));
OR2X2 OR2X2_3049 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9348_));
OR2X2 OR2X2_305 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3044_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3045_));
OR2X2 OR2X2_3050 ( .A(AES_CORE_DATAPATH_iv_2__15_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9350_));
OR2X2 OR2X2_3051 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9351_));
OR2X2 OR2X2_3052 ( .A(AES_CORE_DATAPATH_iv_2__16_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9353_));
OR2X2 OR2X2_3053 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9354_));
OR2X2 OR2X2_3054 ( .A(AES_CORE_DATAPATH_iv_2__17_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9356_));
OR2X2 OR2X2_3055 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9357_));
OR2X2 OR2X2_3056 ( .A(AES_CORE_DATAPATH_iv_2__18_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9359_));
OR2X2 OR2X2_3057 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9360_));
OR2X2 OR2X2_3058 ( .A(AES_CORE_DATAPATH_iv_2__19_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9362_));
OR2X2 OR2X2_3059 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9363_));
OR2X2 OR2X2_306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3047_));
OR2X2 OR2X2_3060 ( .A(AES_CORE_DATAPATH_iv_2__20_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9365_));
OR2X2 OR2X2_3061 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9366_));
OR2X2 OR2X2_3062 ( .A(AES_CORE_DATAPATH_iv_2__21_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9368_));
OR2X2 OR2X2_3063 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9369_));
OR2X2 OR2X2_3064 ( .A(AES_CORE_DATAPATH_iv_2__22_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9371_));
OR2X2 OR2X2_3065 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9372_));
OR2X2 OR2X2_3066 ( .A(AES_CORE_DATAPATH_iv_2__23_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9374_));
OR2X2 OR2X2_3067 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9375_));
OR2X2 OR2X2_3068 ( .A(AES_CORE_DATAPATH_iv_2__24_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9377_));
OR2X2 OR2X2_3069 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9378_));
OR2X2 OR2X2_307 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3049_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3050_));
OR2X2 OR2X2_3070 ( .A(AES_CORE_DATAPATH_iv_2__25_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9380_));
OR2X2 OR2X2_3071 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9381_));
OR2X2 OR2X2_3072 ( .A(AES_CORE_DATAPATH_iv_2__26_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9383_));
OR2X2 OR2X2_3073 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9384_));
OR2X2 OR2X2_3074 ( .A(AES_CORE_DATAPATH_iv_2__27_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9386_));
OR2X2 OR2X2_3075 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9387_));
OR2X2 OR2X2_3076 ( .A(AES_CORE_DATAPATH_iv_2__28_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9389_));
OR2X2 OR2X2_3077 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9390_));
OR2X2 OR2X2_3078 ( .A(AES_CORE_DATAPATH_iv_2__29_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9392_));
OR2X2 OR2X2_3079 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9393_));
OR2X2 OR2X2_308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3053_), .B(AES_CORE_DATAPATH__abc_16009_new_n3054_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3055_));
OR2X2 OR2X2_3080 ( .A(AES_CORE_DATAPATH_iv_2__30_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9395_));
OR2X2 OR2X2_3081 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9396_));
OR2X2 OR2X2_3082 ( .A(AES_CORE_DATAPATH_iv_2__31_), .B(\iv_en[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9398_));
OR2X2 OR2X2_3083 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9305_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9399_));
OR2X2 OR2X2_3084 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9401_), .B(AES_CORE_DATAPATH__abc_16009_new_n9402_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9403_));
OR2X2 OR2X2_3085 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9406_), .B(AES_CORE_DATAPATH__abc_16009_new_n9405_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__0_));
OR2X2 OR2X2_3086 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9409_), .B(AES_CORE_DATAPATH__abc_16009_new_n9408_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__1_));
OR2X2 OR2X2_3087 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9412_), .B(AES_CORE_DATAPATH__abc_16009_new_n9411_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__2_));
OR2X2 OR2X2_3088 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9415_), .B(AES_CORE_DATAPATH__abc_16009_new_n9414_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__3_));
OR2X2 OR2X2_3089 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9418_), .B(AES_CORE_DATAPATH__abc_16009_new_n9417_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__4_));
OR2X2 OR2X2_309 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3055_), .B(AES_CORE_DATAPATH__abc_16009_new_n3052_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3056_));
OR2X2 OR2X2_3090 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9421_), .B(AES_CORE_DATAPATH__abc_16009_new_n9420_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__5_));
OR2X2 OR2X2_3091 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9424_), .B(AES_CORE_DATAPATH__abc_16009_new_n9423_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__6_));
OR2X2 OR2X2_3092 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9427_), .B(AES_CORE_DATAPATH__abc_16009_new_n9426_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__7_));
OR2X2 OR2X2_3093 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9430_), .B(AES_CORE_DATAPATH__abc_16009_new_n9429_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__8_));
OR2X2 OR2X2_3094 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9433_), .B(AES_CORE_DATAPATH__abc_16009_new_n9432_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__9_));
OR2X2 OR2X2_3095 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9436_), .B(AES_CORE_DATAPATH__abc_16009_new_n9435_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__10_));
OR2X2 OR2X2_3096 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9439_), .B(AES_CORE_DATAPATH__abc_16009_new_n9438_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__11_));
OR2X2 OR2X2_3097 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9442_), .B(AES_CORE_DATAPATH__abc_16009_new_n9441_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__12_));
OR2X2 OR2X2_3098 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9445_), .B(AES_CORE_DATAPATH__abc_16009_new_n9444_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__13_));
OR2X2 OR2X2_3099 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9448_), .B(AES_CORE_DATAPATH__abc_16009_new_n9447_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__14_));
OR2X2 OR2X2_31 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n187_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n188_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n189_));
OR2X2 OR2X2_310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3057_));
OR2X2 OR2X2_3100 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9451_), .B(AES_CORE_DATAPATH__abc_16009_new_n9450_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__15_));
OR2X2 OR2X2_3101 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9454_), .B(AES_CORE_DATAPATH__abc_16009_new_n9453_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__16_));
OR2X2 OR2X2_3102 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9457_), .B(AES_CORE_DATAPATH__abc_16009_new_n9456_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__17_));
OR2X2 OR2X2_3103 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9460_), .B(AES_CORE_DATAPATH__abc_16009_new_n9459_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__18_));
OR2X2 OR2X2_3104 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9463_), .B(AES_CORE_DATAPATH__abc_16009_new_n9462_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__19_));
OR2X2 OR2X2_3105 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9466_), .B(AES_CORE_DATAPATH__abc_16009_new_n9465_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__20_));
OR2X2 OR2X2_3106 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9469_), .B(AES_CORE_DATAPATH__abc_16009_new_n9468_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__21_));
OR2X2 OR2X2_3107 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9472_), .B(AES_CORE_DATAPATH__abc_16009_new_n9471_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__22_));
OR2X2 OR2X2_3108 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9475_), .B(AES_CORE_DATAPATH__abc_16009_new_n9474_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__23_));
OR2X2 OR2X2_3109 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9478_), .B(AES_CORE_DATAPATH__abc_16009_new_n9477_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__24_));
OR2X2 OR2X2_311 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3061_), .B(AES_CORE_DATAPATH__abc_16009_new_n3059_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3062_));
OR2X2 OR2X2_3110 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9481_), .B(AES_CORE_DATAPATH__abc_16009_new_n9480_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__25_));
OR2X2 OR2X2_3111 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9484_), .B(AES_CORE_DATAPATH__abc_16009_new_n9483_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__26_));
OR2X2 OR2X2_3112 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9487_), .B(AES_CORE_DATAPATH__abc_16009_new_n9486_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__27_));
OR2X2 OR2X2_3113 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9490_), .B(AES_CORE_DATAPATH__abc_16009_new_n9489_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__28_));
OR2X2 OR2X2_3114 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9493_), .B(AES_CORE_DATAPATH__abc_16009_new_n9492_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__29_));
OR2X2 OR2X2_3115 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9496_), .B(AES_CORE_DATAPATH__abc_16009_new_n9495_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__30_));
OR2X2 OR2X2_3116 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9499_), .B(AES_CORE_DATAPATH__abc_16009_new_n9498_), .Y(AES_CORE_DATAPATH__0bkp_1_2__31_0__31_));
OR2X2 OR2X2_3117 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8016_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9501_));
OR2X2 OR2X2_3118 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9502_));
OR2X2 OR2X2_3119 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9505_));
OR2X2 OR2X2_312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3062_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3063_));
OR2X2 OR2X2_3120 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9504_), .B(AES_CORE_DATAPATH__abc_16009_new_n9505_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9506_));
OR2X2 OR2X2_3121 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9507_));
OR2X2 OR2X2_3122 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8024_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9509_));
OR2X2 OR2X2_3123 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9510_));
OR2X2 OR2X2_3124 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9513_));
OR2X2 OR2X2_3125 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9512_), .B(AES_CORE_DATAPATH__abc_16009_new_n9513_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9514_));
OR2X2 OR2X2_3126 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9515_));
OR2X2 OR2X2_3127 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8032_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9517_));
OR2X2 OR2X2_3128 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9518_));
OR2X2 OR2X2_3129 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8651_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9521_));
OR2X2 OR2X2_313 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3065_));
OR2X2 OR2X2_3130 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9520_), .B(AES_CORE_DATAPATH__abc_16009_new_n9521_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9522_));
OR2X2 OR2X2_3131 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9523_));
OR2X2 OR2X2_3132 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8040_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9525_));
OR2X2 OR2X2_3133 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9526_));
OR2X2 OR2X2_3134 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8660_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9529_));
OR2X2 OR2X2_3135 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9528_), .B(AES_CORE_DATAPATH__abc_16009_new_n9529_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9530_));
OR2X2 OR2X2_3136 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9531_));
OR2X2 OR2X2_3137 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8048_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9533_));
OR2X2 OR2X2_3138 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9534_));
OR2X2 OR2X2_3139 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8669_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9537_));
OR2X2 OR2X2_314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3067_));
OR2X2 OR2X2_3140 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9536_), .B(AES_CORE_DATAPATH__abc_16009_new_n9537_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9538_));
OR2X2 OR2X2_3141 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9539_));
OR2X2 OR2X2_3142 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8056_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9541_));
OR2X2 OR2X2_3143 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9542_));
OR2X2 OR2X2_3144 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8678_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9545_));
OR2X2 OR2X2_3145 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9544_), .B(AES_CORE_DATAPATH__abc_16009_new_n9545_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9546_));
OR2X2 OR2X2_3146 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9547_));
OR2X2 OR2X2_3147 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8064_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9549_));
OR2X2 OR2X2_3148 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9550_));
OR2X2 OR2X2_3149 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9553_));
OR2X2 OR2X2_315 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3068_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3069_));
OR2X2 OR2X2_3150 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9552_), .B(AES_CORE_DATAPATH__abc_16009_new_n9553_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9554_));
OR2X2 OR2X2_3151 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9555_));
OR2X2 OR2X2_3152 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8072_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9557_));
OR2X2 OR2X2_3153 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9558_));
OR2X2 OR2X2_3154 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8696_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9561_));
OR2X2 OR2X2_3155 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9560_), .B(AES_CORE_DATAPATH__abc_16009_new_n9561_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9562_));
OR2X2 OR2X2_3156 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9563_));
OR2X2 OR2X2_3157 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8080_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9565_));
OR2X2 OR2X2_3158 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9566_));
OR2X2 OR2X2_3159 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8705_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9569_));
OR2X2 OR2X2_316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3072_), .B(AES_CORE_DATAPATH__abc_16009_new_n3073_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3074_));
OR2X2 OR2X2_3160 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9568_), .B(AES_CORE_DATAPATH__abc_16009_new_n9569_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9570_));
OR2X2 OR2X2_3161 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9571_));
OR2X2 OR2X2_3162 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8088_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9573_));
OR2X2 OR2X2_3163 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9574_));
OR2X2 OR2X2_3164 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8714_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9577_));
OR2X2 OR2X2_3165 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9576_), .B(AES_CORE_DATAPATH__abc_16009_new_n9577_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9578_));
OR2X2 OR2X2_3166 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9579_));
OR2X2 OR2X2_3167 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8096_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9581_));
OR2X2 OR2X2_3168 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9582_));
OR2X2 OR2X2_3169 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8723_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9585_));
OR2X2 OR2X2_317 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3074_), .B(AES_CORE_DATAPATH__abc_16009_new_n3071_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3075_));
OR2X2 OR2X2_3170 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9584_), .B(AES_CORE_DATAPATH__abc_16009_new_n9585_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9586_));
OR2X2 OR2X2_3171 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9587_));
OR2X2 OR2X2_3172 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8104_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9589_));
OR2X2 OR2X2_3173 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9590_));
OR2X2 OR2X2_3174 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8732_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9593_));
OR2X2 OR2X2_3175 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9592_), .B(AES_CORE_DATAPATH__abc_16009_new_n9593_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9594_));
OR2X2 OR2X2_3176 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9595_));
OR2X2 OR2X2_3177 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8112_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9597_));
OR2X2 OR2X2_3178 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9598_));
OR2X2 OR2X2_3179 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8741_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9601_));
OR2X2 OR2X2_318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3079_), .B(AES_CORE_DATAPATH__abc_16009_new_n3077_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3080_));
OR2X2 OR2X2_3180 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9600_), .B(AES_CORE_DATAPATH__abc_16009_new_n9601_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9602_));
OR2X2 OR2X2_3181 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9603_));
OR2X2 OR2X2_3182 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8120_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9605_));
OR2X2 OR2X2_3183 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9606_));
OR2X2 OR2X2_3184 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8750_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9609_));
OR2X2 OR2X2_3185 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9608_), .B(AES_CORE_DATAPATH__abc_16009_new_n9609_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9610_));
OR2X2 OR2X2_3186 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9611_));
OR2X2 OR2X2_3187 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8128_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9613_));
OR2X2 OR2X2_3188 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9614_));
OR2X2 OR2X2_3189 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9617_));
OR2X2 OR2X2_319 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3080_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3081_));
OR2X2 OR2X2_3190 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9616_), .B(AES_CORE_DATAPATH__abc_16009_new_n9617_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9618_));
OR2X2 OR2X2_3191 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9619_));
OR2X2 OR2X2_3192 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8136_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9621_));
OR2X2 OR2X2_3193 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9622_));
OR2X2 OR2X2_3194 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8768_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9625_));
OR2X2 OR2X2_3195 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9624_), .B(AES_CORE_DATAPATH__abc_16009_new_n9625_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9626_));
OR2X2 OR2X2_3196 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9627_));
OR2X2 OR2X2_3197 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8144_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9629_));
OR2X2 OR2X2_3198 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9630_));
OR2X2 OR2X2_3199 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9633_));
OR2X2 OR2X2_32 ( .A(AES_CORE_CONTROL_UNIT_state_14_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n191_));
OR2X2 OR2X2_320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3083_));
OR2X2 OR2X2_3200 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9632_), .B(AES_CORE_DATAPATH__abc_16009_new_n9633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9634_));
OR2X2 OR2X2_3201 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9635_));
OR2X2 OR2X2_3202 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8152_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9637_));
OR2X2 OR2X2_3203 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9638_));
OR2X2 OR2X2_3204 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8786_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9641_));
OR2X2 OR2X2_3205 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9640_), .B(AES_CORE_DATAPATH__abc_16009_new_n9641_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9642_));
OR2X2 OR2X2_3206 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9643_));
OR2X2 OR2X2_3207 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8160_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9645_));
OR2X2 OR2X2_3208 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9646_));
OR2X2 OR2X2_3209 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8795_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9649_));
OR2X2 OR2X2_321 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3085_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3086_));
OR2X2 OR2X2_3210 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9648_), .B(AES_CORE_DATAPATH__abc_16009_new_n9649_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9650_));
OR2X2 OR2X2_3211 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9651_));
OR2X2 OR2X2_3212 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8168_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9653_));
OR2X2 OR2X2_3213 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9654_));
OR2X2 OR2X2_3214 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8804_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9657_));
OR2X2 OR2X2_3215 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9656_), .B(AES_CORE_DATAPATH__abc_16009_new_n9657_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9658_));
OR2X2 OR2X2_3216 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9659_));
OR2X2 OR2X2_3217 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8176_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9661_));
OR2X2 OR2X2_3218 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9662_));
OR2X2 OR2X2_3219 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9665_));
OR2X2 OR2X2_322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3089_), .B(AES_CORE_DATAPATH__abc_16009_new_n3090_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3091_));
OR2X2 OR2X2_3220 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9664_), .B(AES_CORE_DATAPATH__abc_16009_new_n9665_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9666_));
OR2X2 OR2X2_3221 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9667_));
OR2X2 OR2X2_3222 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8184_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9669_));
OR2X2 OR2X2_3223 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9670_));
OR2X2 OR2X2_3224 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9673_));
OR2X2 OR2X2_3225 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9672_), .B(AES_CORE_DATAPATH__abc_16009_new_n9673_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9674_));
OR2X2 OR2X2_3226 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9675_));
OR2X2 OR2X2_3227 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8192_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9677_));
OR2X2 OR2X2_3228 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9678_));
OR2X2 OR2X2_3229 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9681_));
OR2X2 OR2X2_323 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3091_), .B(AES_CORE_DATAPATH__abc_16009_new_n3088_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3092_));
OR2X2 OR2X2_3230 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9680_), .B(AES_CORE_DATAPATH__abc_16009_new_n9681_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9682_));
OR2X2 OR2X2_3231 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9683_));
OR2X2 OR2X2_3232 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8200_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9685_));
OR2X2 OR2X2_3233 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9686_));
OR2X2 OR2X2_3234 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8840_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9689_));
OR2X2 OR2X2_3235 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9688_), .B(AES_CORE_DATAPATH__abc_16009_new_n9689_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9690_));
OR2X2 OR2X2_3236 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9691_));
OR2X2 OR2X2_3237 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8208_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9693_));
OR2X2 OR2X2_3238 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9694_));
OR2X2 OR2X2_3239 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8849_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9697_));
OR2X2 OR2X2_324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3093_));
OR2X2 OR2X2_3240 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9696_), .B(AES_CORE_DATAPATH__abc_16009_new_n9697_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9698_));
OR2X2 OR2X2_3241 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9699_));
OR2X2 OR2X2_3242 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8216_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9701_));
OR2X2 OR2X2_3243 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9702_));
OR2X2 OR2X2_3244 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8858_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9705_));
OR2X2 OR2X2_3245 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9704_), .B(AES_CORE_DATAPATH__abc_16009_new_n9705_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9706_));
OR2X2 OR2X2_3246 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9707_));
OR2X2 OR2X2_3247 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8224_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9709_));
OR2X2 OR2X2_3248 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9710_));
OR2X2 OR2X2_3249 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9713_));
OR2X2 OR2X2_325 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3097_), .B(AES_CORE_DATAPATH__abc_16009_new_n3095_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3098_));
OR2X2 OR2X2_3250 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9712_), .B(AES_CORE_DATAPATH__abc_16009_new_n9713_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9714_));
OR2X2 OR2X2_3251 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9715_));
OR2X2 OR2X2_3252 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8232_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9717_));
OR2X2 OR2X2_3253 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9718_));
OR2X2 OR2X2_3254 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8876_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9721_));
OR2X2 OR2X2_3255 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9720_), .B(AES_CORE_DATAPATH__abc_16009_new_n9721_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9722_));
OR2X2 OR2X2_3256 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9723_));
OR2X2 OR2X2_3257 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8240_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9725_));
OR2X2 OR2X2_3258 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9726_));
OR2X2 OR2X2_3259 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8885_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9729_));
OR2X2 OR2X2_326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3098_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3099_));
OR2X2 OR2X2_3260 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9728_), .B(AES_CORE_DATAPATH__abc_16009_new_n9729_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9730_));
OR2X2 OR2X2_3261 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9731_));
OR2X2 OR2X2_3262 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8248_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9733_));
OR2X2 OR2X2_3263 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9734_));
OR2X2 OR2X2_3264 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8894_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9737_));
OR2X2 OR2X2_3265 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9736_), .B(AES_CORE_DATAPATH__abc_16009_new_n9737_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9738_));
OR2X2 OR2X2_3266 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9739_));
OR2X2 OR2X2_3267 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8256_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9741_));
OR2X2 OR2X2_3268 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9742_));
OR2X2 OR2X2_3269 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8903_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9745_));
OR2X2 OR2X2_327 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3101_));
OR2X2 OR2X2_3270 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9744_), .B(AES_CORE_DATAPATH__abc_16009_new_n9745_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9746_));
OR2X2 OR2X2_3271 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9747_));
OR2X2 OR2X2_3272 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8264_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9749_));
OR2X2 OR2X2_3273 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9750_));
OR2X2 OR2X2_3274 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9404_), .B(AES_CORE_DATAPATH__abc_16009_new_n8912_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9753_));
OR2X2 OR2X2_3275 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9752_), .B(AES_CORE_DATAPATH__abc_16009_new_n9753_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9754_));
OR2X2 OR2X2_3276 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9403_), .B(AES_CORE_DATAPATH_bkp_2__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9755_));
OR2X2 OR2X2_3277 ( .A(AES_CORE_DATAPATH_iv_1__0_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9757_));
OR2X2 OR2X2_3278 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9759_));
OR2X2 OR2X2_3279 ( .A(AES_CORE_DATAPATH_iv_1__1_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9761_));
OR2X2 OR2X2_328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3103_));
OR2X2 OR2X2_3280 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9762_));
OR2X2 OR2X2_3281 ( .A(AES_CORE_DATAPATH_iv_1__2_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9764_));
OR2X2 OR2X2_3282 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9765_));
OR2X2 OR2X2_3283 ( .A(AES_CORE_DATAPATH_iv_1__3_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9767_));
OR2X2 OR2X2_3284 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9768_));
OR2X2 OR2X2_3285 ( .A(AES_CORE_DATAPATH_iv_1__4_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9770_));
OR2X2 OR2X2_3286 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9771_));
OR2X2 OR2X2_3287 ( .A(AES_CORE_DATAPATH_iv_1__5_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9773_));
OR2X2 OR2X2_3288 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9774_));
OR2X2 OR2X2_3289 ( .A(AES_CORE_DATAPATH_iv_1__6_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9776_));
OR2X2 OR2X2_329 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3104_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3105_));
OR2X2 OR2X2_3290 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9777_));
OR2X2 OR2X2_3291 ( .A(AES_CORE_DATAPATH_iv_1__7_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9779_));
OR2X2 OR2X2_3292 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9780_));
OR2X2 OR2X2_3293 ( .A(AES_CORE_DATAPATH_iv_1__8_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9782_));
OR2X2 OR2X2_3294 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9783_));
OR2X2 OR2X2_3295 ( .A(AES_CORE_DATAPATH_iv_1__9_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9785_));
OR2X2 OR2X2_3296 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9786_));
OR2X2 OR2X2_3297 ( .A(AES_CORE_DATAPATH_iv_1__10_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9788_));
OR2X2 OR2X2_3298 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9789_));
OR2X2 OR2X2_3299 ( .A(AES_CORE_DATAPATH_iv_1__11_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9791_));
OR2X2 OR2X2_33 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .B(AES_CORE_CONTROL_UNIT_state_6_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n192_));
OR2X2 OR2X2_330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3108_), .B(AES_CORE_DATAPATH__abc_16009_new_n3109_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3110_));
OR2X2 OR2X2_3300 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9792_));
OR2X2 OR2X2_3301 ( .A(AES_CORE_DATAPATH_iv_1__12_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9794_));
OR2X2 OR2X2_3302 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9795_));
OR2X2 OR2X2_3303 ( .A(AES_CORE_DATAPATH_iv_1__13_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9797_));
OR2X2 OR2X2_3304 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9798_));
OR2X2 OR2X2_3305 ( .A(AES_CORE_DATAPATH_iv_1__14_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9800_));
OR2X2 OR2X2_3306 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9801_));
OR2X2 OR2X2_3307 ( .A(AES_CORE_DATAPATH_iv_1__15_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9803_));
OR2X2 OR2X2_3308 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9804_));
OR2X2 OR2X2_3309 ( .A(AES_CORE_DATAPATH_iv_1__16_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9806_));
OR2X2 OR2X2_331 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3110_), .B(AES_CORE_DATAPATH__abc_16009_new_n3107_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3111_));
OR2X2 OR2X2_3310 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9807_));
OR2X2 OR2X2_3311 ( .A(AES_CORE_DATAPATH_iv_1__17_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9809_));
OR2X2 OR2X2_3312 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9810_));
OR2X2 OR2X2_3313 ( .A(AES_CORE_DATAPATH_iv_1__18_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9812_));
OR2X2 OR2X2_3314 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9813_));
OR2X2 OR2X2_3315 ( .A(AES_CORE_DATAPATH_iv_1__19_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9815_));
OR2X2 OR2X2_3316 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9816_));
OR2X2 OR2X2_3317 ( .A(AES_CORE_DATAPATH_iv_1__20_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9818_));
OR2X2 OR2X2_3318 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9819_));
OR2X2 OR2X2_3319 ( .A(AES_CORE_DATAPATH_iv_1__21_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9821_));
OR2X2 OR2X2_332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3115_), .B(AES_CORE_DATAPATH__abc_16009_new_n3113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3116_));
OR2X2 OR2X2_3320 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9822_));
OR2X2 OR2X2_3321 ( .A(AES_CORE_DATAPATH_iv_1__22_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9824_));
OR2X2 OR2X2_3322 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9825_));
OR2X2 OR2X2_3323 ( .A(AES_CORE_DATAPATH_iv_1__23_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9827_));
OR2X2 OR2X2_3324 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9828_));
OR2X2 OR2X2_3325 ( .A(AES_CORE_DATAPATH_iv_1__24_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9830_));
OR2X2 OR2X2_3326 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9831_));
OR2X2 OR2X2_3327 ( .A(AES_CORE_DATAPATH_iv_1__25_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9833_));
OR2X2 OR2X2_3328 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9834_));
OR2X2 OR2X2_3329 ( .A(AES_CORE_DATAPATH_iv_1__26_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9836_));
OR2X2 OR2X2_333 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3116_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3117_));
OR2X2 OR2X2_3330 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9837_));
OR2X2 OR2X2_3331 ( .A(AES_CORE_DATAPATH_iv_1__27_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9839_));
OR2X2 OR2X2_3332 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9840_));
OR2X2 OR2X2_3333 ( .A(AES_CORE_DATAPATH_iv_1__28_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9842_));
OR2X2 OR2X2_3334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9843_));
OR2X2 OR2X2_3335 ( .A(AES_CORE_DATAPATH_iv_1__29_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9845_));
OR2X2 OR2X2_3336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9846_));
OR2X2 OR2X2_3337 ( .A(AES_CORE_DATAPATH_iv_1__30_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9848_));
OR2X2 OR2X2_3338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9849_));
OR2X2 OR2X2_3339 ( .A(AES_CORE_DATAPATH_iv_1__31_), .B(\iv_en[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9851_));
OR2X2 OR2X2_334 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3121_));
OR2X2 OR2X2_3340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9758_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n9852_));
OR2X2 OR2X2_3341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9854_), .B(AES_CORE_DATAPATH__abc_16009_new_n9855_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9856_));
OR2X2 OR2X2_3342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9859_), .B(AES_CORE_DATAPATH__abc_16009_new_n9858_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__0_));
OR2X2 OR2X2_3343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9862_), .B(AES_CORE_DATAPATH__abc_16009_new_n9861_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__1_));
OR2X2 OR2X2_3344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9865_), .B(AES_CORE_DATAPATH__abc_16009_new_n9864_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__2_));
OR2X2 OR2X2_3345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9868_), .B(AES_CORE_DATAPATH__abc_16009_new_n9867_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__3_));
OR2X2 OR2X2_3346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9871_), .B(AES_CORE_DATAPATH__abc_16009_new_n9870_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__4_));
OR2X2 OR2X2_3347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9874_), .B(AES_CORE_DATAPATH__abc_16009_new_n9873_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__5_));
OR2X2 OR2X2_3348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9877_), .B(AES_CORE_DATAPATH__abc_16009_new_n9876_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__6_));
OR2X2 OR2X2_3349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9880_), .B(AES_CORE_DATAPATH__abc_16009_new_n9879_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__7_));
OR2X2 OR2X2_335 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3122_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3123_));
OR2X2 OR2X2_3350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9883_), .B(AES_CORE_DATAPATH__abc_16009_new_n9882_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__8_));
OR2X2 OR2X2_3351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9886_), .B(AES_CORE_DATAPATH__abc_16009_new_n9885_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__9_));
OR2X2 OR2X2_3352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9889_), .B(AES_CORE_DATAPATH__abc_16009_new_n9888_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__10_));
OR2X2 OR2X2_3353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9892_), .B(AES_CORE_DATAPATH__abc_16009_new_n9891_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__11_));
OR2X2 OR2X2_3354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9895_), .B(AES_CORE_DATAPATH__abc_16009_new_n9894_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__12_));
OR2X2 OR2X2_3355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9898_), .B(AES_CORE_DATAPATH__abc_16009_new_n9897_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__13_));
OR2X2 OR2X2_3356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9901_), .B(AES_CORE_DATAPATH__abc_16009_new_n9900_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__14_));
OR2X2 OR2X2_3357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9904_), .B(AES_CORE_DATAPATH__abc_16009_new_n9903_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__15_));
OR2X2 OR2X2_3358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9907_), .B(AES_CORE_DATAPATH__abc_16009_new_n9906_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__16_));
OR2X2 OR2X2_3359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9910_), .B(AES_CORE_DATAPATH__abc_16009_new_n9909_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__17_));
OR2X2 OR2X2_336 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3126_), .B(AES_CORE_DATAPATH__abc_16009_new_n3127_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3128_));
OR2X2 OR2X2_3360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9913_), .B(AES_CORE_DATAPATH__abc_16009_new_n9912_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__18_));
OR2X2 OR2X2_3361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9916_), .B(AES_CORE_DATAPATH__abc_16009_new_n9915_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__19_));
OR2X2 OR2X2_3362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9919_), .B(AES_CORE_DATAPATH__abc_16009_new_n9918_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__20_));
OR2X2 OR2X2_3363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9922_), .B(AES_CORE_DATAPATH__abc_16009_new_n9921_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__21_));
OR2X2 OR2X2_3364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9925_), .B(AES_CORE_DATAPATH__abc_16009_new_n9924_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__22_));
OR2X2 OR2X2_3365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9928_), .B(AES_CORE_DATAPATH__abc_16009_new_n9927_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__23_));
OR2X2 OR2X2_3366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9931_), .B(AES_CORE_DATAPATH__abc_16009_new_n9930_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__24_));
OR2X2 OR2X2_3367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9934_), .B(AES_CORE_DATAPATH__abc_16009_new_n9933_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__25_));
OR2X2 OR2X2_3368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9937_), .B(AES_CORE_DATAPATH__abc_16009_new_n9936_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__26_));
OR2X2 OR2X2_3369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9940_), .B(AES_CORE_DATAPATH__abc_16009_new_n9939_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__27_));
OR2X2 OR2X2_337 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3128_), .B(AES_CORE_DATAPATH__abc_16009_new_n3125_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3129_));
OR2X2 OR2X2_3370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9943_), .B(AES_CORE_DATAPATH__abc_16009_new_n9942_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__28_));
OR2X2 OR2X2_3371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9946_), .B(AES_CORE_DATAPATH__abc_16009_new_n9945_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__29_));
OR2X2 OR2X2_3372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9949_), .B(AES_CORE_DATAPATH__abc_16009_new_n9948_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__30_));
OR2X2 OR2X2_3373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9952_), .B(AES_CORE_DATAPATH__abc_16009_new_n9951_), .Y(AES_CORE_DATAPATH__0bkp_1_1__31_0__31_));
OR2X2 OR2X2_3374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8273_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9954_));
OR2X2 OR2X2_3375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9955_));
OR2X2 OR2X2_3376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9958_));
OR2X2 OR2X2_3377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9957_), .B(AES_CORE_DATAPATH__abc_16009_new_n9958_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9959_));
OR2X2 OR2X2_3378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9960_));
OR2X2 OR2X2_3379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8281_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9962_));
OR2X2 OR2X2_338 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3131_), .B(AES_CORE_DATAPATH__abc_16009_new_n3120_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3132_));
OR2X2 OR2X2_3380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9963_));
OR2X2 OR2X2_3381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9966_));
OR2X2 OR2X2_3382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9965_), .B(AES_CORE_DATAPATH__abc_16009_new_n9966_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9967_));
OR2X2 OR2X2_3383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9968_));
OR2X2 OR2X2_3384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8289_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9970_));
OR2X2 OR2X2_3385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9971_));
OR2X2 OR2X2_3386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8651_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9974_));
OR2X2 OR2X2_3387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9973_), .B(AES_CORE_DATAPATH__abc_16009_new_n9974_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9975_));
OR2X2 OR2X2_3388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9976_));
OR2X2 OR2X2_3389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8297_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9978_));
OR2X2 OR2X2_339 ( .A(\key_out[16] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3133_));
OR2X2 OR2X2_3390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9979_));
OR2X2 OR2X2_3391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8660_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9982_));
OR2X2 OR2X2_3392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9981_), .B(AES_CORE_DATAPATH__abc_16009_new_n9982_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9983_));
OR2X2 OR2X2_3393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9984_));
OR2X2 OR2X2_3394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8305_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9986_));
OR2X2 OR2X2_3395 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9987_));
OR2X2 OR2X2_3396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8669_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9990_));
OR2X2 OR2X2_3397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9989_), .B(AES_CORE_DATAPATH__abc_16009_new_n9990_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9991_));
OR2X2 OR2X2_3398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9992_));
OR2X2 OR2X2_3399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8313_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9994_));
OR2X2 OR2X2_34 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n191_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n192_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n193_));
OR2X2 OR2X2_340 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3135_), .B(AES_CORE_DATAPATH__abc_16009_new_n3119_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__16_));
OR2X2 OR2X2_3400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9995_));
OR2X2 OR2X2_3401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8678_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9998_));
OR2X2 OR2X2_3402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9997_), .B(AES_CORE_DATAPATH__abc_16009_new_n9998_), .Y(AES_CORE_DATAPATH__abc_16009_new_n9999_));
OR2X2 OR2X2_3403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10000_));
OR2X2 OR2X2_3404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8321_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10002_));
OR2X2 OR2X2_3405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10003_));
OR2X2 OR2X2_3406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10006_));
OR2X2 OR2X2_3407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10005_), .B(AES_CORE_DATAPATH__abc_16009_new_n10006_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10007_));
OR2X2 OR2X2_3408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10008_));
OR2X2 OR2X2_3409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8329_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10010_));
OR2X2 OR2X2_341 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3137_));
OR2X2 OR2X2_3410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10011_));
OR2X2 OR2X2_3411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8696_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10014_));
OR2X2 OR2X2_3412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10013_), .B(AES_CORE_DATAPATH__abc_16009_new_n10014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10015_));
OR2X2 OR2X2_3413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10016_));
OR2X2 OR2X2_3414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8337_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10018_));
OR2X2 OR2X2_3415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10019_));
OR2X2 OR2X2_3416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8705_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10022_));
OR2X2 OR2X2_3417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10021_), .B(AES_CORE_DATAPATH__abc_16009_new_n10022_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10023_));
OR2X2 OR2X2_3418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10024_));
OR2X2 OR2X2_3419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8345_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10026_));
OR2X2 OR2X2_342 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3139_));
OR2X2 OR2X2_3420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10027_));
OR2X2 OR2X2_3421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8714_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10030_));
OR2X2 OR2X2_3422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10029_), .B(AES_CORE_DATAPATH__abc_16009_new_n10030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10031_));
OR2X2 OR2X2_3423 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10032_));
OR2X2 OR2X2_3424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8353_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10034_));
OR2X2 OR2X2_3425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10035_));
OR2X2 OR2X2_3426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8723_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10038_));
OR2X2 OR2X2_3427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10037_), .B(AES_CORE_DATAPATH__abc_16009_new_n10038_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10039_));
OR2X2 OR2X2_3428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10040_));
OR2X2 OR2X2_3429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8361_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10042_));
OR2X2 OR2X2_343 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3140_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3141_));
OR2X2 OR2X2_3430 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10043_));
OR2X2 OR2X2_3431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8732_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10046_));
OR2X2 OR2X2_3432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10045_), .B(AES_CORE_DATAPATH__abc_16009_new_n10046_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10047_));
OR2X2 OR2X2_3433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10048_));
OR2X2 OR2X2_3434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8369_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10050_));
OR2X2 OR2X2_3435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10051_));
OR2X2 OR2X2_3436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8741_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10054_));
OR2X2 OR2X2_3437 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10053_), .B(AES_CORE_DATAPATH__abc_16009_new_n10054_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10055_));
OR2X2 OR2X2_3438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10056_));
OR2X2 OR2X2_3439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8377_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10058_));
OR2X2 OR2X2_344 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3144_), .B(AES_CORE_DATAPATH__abc_16009_new_n3145_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3146_));
OR2X2 OR2X2_3440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10059_));
OR2X2 OR2X2_3441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8750_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10062_));
OR2X2 OR2X2_3442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10061_), .B(AES_CORE_DATAPATH__abc_16009_new_n10062_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10063_));
OR2X2 OR2X2_3443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10064_));
OR2X2 OR2X2_3444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8385_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10066_));
OR2X2 OR2X2_3445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10067_));
OR2X2 OR2X2_3446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10070_));
OR2X2 OR2X2_3447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10069_), .B(AES_CORE_DATAPATH__abc_16009_new_n10070_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10071_));
OR2X2 OR2X2_3448 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10072_));
OR2X2 OR2X2_3449 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8393_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10074_));
OR2X2 OR2X2_345 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3146_), .B(AES_CORE_DATAPATH__abc_16009_new_n3143_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3147_));
OR2X2 OR2X2_3450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10075_));
OR2X2 OR2X2_3451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8768_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10078_));
OR2X2 OR2X2_3452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10077_), .B(AES_CORE_DATAPATH__abc_16009_new_n10078_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10079_));
OR2X2 OR2X2_3453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10080_));
OR2X2 OR2X2_3454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8401_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10082_));
OR2X2 OR2X2_3455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10083_));
OR2X2 OR2X2_3456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10086_));
OR2X2 OR2X2_3457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10085_), .B(AES_CORE_DATAPATH__abc_16009_new_n10086_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10087_));
OR2X2 OR2X2_3458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10088_));
OR2X2 OR2X2_3459 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8409_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10090_));
OR2X2 OR2X2_346 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3151_), .B(AES_CORE_DATAPATH__abc_16009_new_n3149_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3152_));
OR2X2 OR2X2_3460 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10091_));
OR2X2 OR2X2_3461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8786_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10094_));
OR2X2 OR2X2_3462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10093_), .B(AES_CORE_DATAPATH__abc_16009_new_n10094_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10095_));
OR2X2 OR2X2_3463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10096_));
OR2X2 OR2X2_3464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8417_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10098_));
OR2X2 OR2X2_3465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10099_));
OR2X2 OR2X2_3466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8795_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10102_));
OR2X2 OR2X2_3467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10101_), .B(AES_CORE_DATAPATH__abc_16009_new_n10102_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10103_));
OR2X2 OR2X2_3468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10104_));
OR2X2 OR2X2_3469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8425_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10106_));
OR2X2 OR2X2_347 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3152_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3153_));
OR2X2 OR2X2_3470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10107_));
OR2X2 OR2X2_3471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8804_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10110_));
OR2X2 OR2X2_3472 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10109_), .B(AES_CORE_DATAPATH__abc_16009_new_n10110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10111_));
OR2X2 OR2X2_3473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10112_));
OR2X2 OR2X2_3474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8433_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10114_));
OR2X2 OR2X2_3475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10115_));
OR2X2 OR2X2_3476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10118_));
OR2X2 OR2X2_3477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10117_), .B(AES_CORE_DATAPATH__abc_16009_new_n10118_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10119_));
OR2X2 OR2X2_3478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10120_));
OR2X2 OR2X2_3479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8441_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10122_));
OR2X2 OR2X2_348 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3155_));
OR2X2 OR2X2_3480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10123_));
OR2X2 OR2X2_3481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10126_));
OR2X2 OR2X2_3482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10125_), .B(AES_CORE_DATAPATH__abc_16009_new_n10126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10127_));
OR2X2 OR2X2_3483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10128_));
OR2X2 OR2X2_3484 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8449_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10130_));
OR2X2 OR2X2_3485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10131_));
OR2X2 OR2X2_3486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10134_));
OR2X2 OR2X2_3487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10133_), .B(AES_CORE_DATAPATH__abc_16009_new_n10134_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10135_));
OR2X2 OR2X2_3488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10136_));
OR2X2 OR2X2_3489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8457_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10138_));
OR2X2 OR2X2_349 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3157_));
OR2X2 OR2X2_3490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10139_));
OR2X2 OR2X2_3491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8840_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10142_));
OR2X2 OR2X2_3492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10141_), .B(AES_CORE_DATAPATH__abc_16009_new_n10142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10143_));
OR2X2 OR2X2_3493 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10144_));
OR2X2 OR2X2_3494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8465_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10146_));
OR2X2 OR2X2_3495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10147_));
OR2X2 OR2X2_3496 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8849_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10150_));
OR2X2 OR2X2_3497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10149_), .B(AES_CORE_DATAPATH__abc_16009_new_n10150_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10151_));
OR2X2 OR2X2_3498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10152_));
OR2X2 OR2X2_3499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8473_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10154_));
OR2X2 OR2X2_35 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n144_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n145_), .Y(AES_CORE_CONTROL_UNIT_col_en_0_));
OR2X2 OR2X2_350 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3158_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3159_));
OR2X2 OR2X2_3500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10155_));
OR2X2 OR2X2_3501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8858_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10158_));
OR2X2 OR2X2_3502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10157_), .B(AES_CORE_DATAPATH__abc_16009_new_n10158_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10159_));
OR2X2 OR2X2_3503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10160_));
OR2X2 OR2X2_3504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8481_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10162_));
OR2X2 OR2X2_3505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10163_));
OR2X2 OR2X2_3506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10166_));
OR2X2 OR2X2_3507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10165_), .B(AES_CORE_DATAPATH__abc_16009_new_n10166_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10167_));
OR2X2 OR2X2_3508 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10168_));
OR2X2 OR2X2_3509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8489_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10170_));
OR2X2 OR2X2_351 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3162_), .B(AES_CORE_DATAPATH__abc_16009_new_n3163_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3164_));
OR2X2 OR2X2_3510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10171_));
OR2X2 OR2X2_3511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8876_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10174_));
OR2X2 OR2X2_3512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10173_), .B(AES_CORE_DATAPATH__abc_16009_new_n10174_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10175_));
OR2X2 OR2X2_3513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10176_));
OR2X2 OR2X2_3514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8497_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10178_));
OR2X2 OR2X2_3515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10179_));
OR2X2 OR2X2_3516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8885_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10182_));
OR2X2 OR2X2_3517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10181_), .B(AES_CORE_DATAPATH__abc_16009_new_n10182_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10183_));
OR2X2 OR2X2_3518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10184_));
OR2X2 OR2X2_3519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8505_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10186_));
OR2X2 OR2X2_352 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3164_), .B(AES_CORE_DATAPATH__abc_16009_new_n3161_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3165_));
OR2X2 OR2X2_3520 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10187_));
OR2X2 OR2X2_3521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8894_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10190_));
OR2X2 OR2X2_3522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10189_), .B(AES_CORE_DATAPATH__abc_16009_new_n10190_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10191_));
OR2X2 OR2X2_3523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10192_));
OR2X2 OR2X2_3524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8513_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10194_));
OR2X2 OR2X2_3525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10195_));
OR2X2 OR2X2_3526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8903_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10198_));
OR2X2 OR2X2_3527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10197_), .B(AES_CORE_DATAPATH__abc_16009_new_n10198_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10199_));
OR2X2 OR2X2_3528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10200_));
OR2X2 OR2X2_3529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8521_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10202_));
OR2X2 OR2X2_353 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3169_), .B(AES_CORE_DATAPATH__abc_16009_new_n3167_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3170_));
OR2X2 OR2X2_3530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10203_));
OR2X2 OR2X2_3531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9857_), .B(AES_CORE_DATAPATH__abc_16009_new_n8912_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10206_));
OR2X2 OR2X2_3532 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10205_), .B(AES_CORE_DATAPATH__abc_16009_new_n10206_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10207_));
OR2X2 OR2X2_3533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n9856_), .B(AES_CORE_DATAPATH_bkp_1__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10208_));
OR2X2 OR2X2_3534 ( .A(AES_CORE_DATAPATH_iv_0__0_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10210_));
OR2X2 OR2X2_3535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10212_));
OR2X2 OR2X2_3536 ( .A(AES_CORE_DATAPATH_iv_0__1_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10214_));
OR2X2 OR2X2_3537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10215_));
OR2X2 OR2X2_3538 ( .A(AES_CORE_DATAPATH_iv_0__2_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10217_));
OR2X2 OR2X2_3539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10218_));
OR2X2 OR2X2_354 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3170_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3171_));
OR2X2 OR2X2_3540 ( .A(AES_CORE_DATAPATH_iv_0__3_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10220_));
OR2X2 OR2X2_3541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10221_));
OR2X2 OR2X2_3542 ( .A(AES_CORE_DATAPATH_iv_0__4_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10223_));
OR2X2 OR2X2_3543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[4] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10224_));
OR2X2 OR2X2_3544 ( .A(AES_CORE_DATAPATH_iv_0__5_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10226_));
OR2X2 OR2X2_3545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[5] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10227_));
OR2X2 OR2X2_3546 ( .A(AES_CORE_DATAPATH_iv_0__6_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10229_));
OR2X2 OR2X2_3547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[6] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10230_));
OR2X2 OR2X2_3548 ( .A(AES_CORE_DATAPATH_iv_0__7_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10232_));
OR2X2 OR2X2_3549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[7] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10233_));
OR2X2 OR2X2_355 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3173_));
OR2X2 OR2X2_3550 ( .A(AES_CORE_DATAPATH_iv_0__8_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10235_));
OR2X2 OR2X2_3551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[8] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10236_));
OR2X2 OR2X2_3552 ( .A(AES_CORE_DATAPATH_iv_0__9_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10238_));
OR2X2 OR2X2_3553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[9] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10239_));
OR2X2 OR2X2_3554 ( .A(AES_CORE_DATAPATH_iv_0__10_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10241_));
OR2X2 OR2X2_3555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[10] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10242_));
OR2X2 OR2X2_3556 ( .A(AES_CORE_DATAPATH_iv_0__11_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10244_));
OR2X2 OR2X2_3557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[11] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10245_));
OR2X2 OR2X2_3558 ( .A(AES_CORE_DATAPATH_iv_0__12_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10247_));
OR2X2 OR2X2_3559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[12] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10248_));
OR2X2 OR2X2_356 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3175_));
OR2X2 OR2X2_3560 ( .A(AES_CORE_DATAPATH_iv_0__13_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10250_));
OR2X2 OR2X2_3561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[13] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10251_));
OR2X2 OR2X2_3562 ( .A(AES_CORE_DATAPATH_iv_0__14_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10253_));
OR2X2 OR2X2_3563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[14] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10254_));
OR2X2 OR2X2_3564 ( .A(AES_CORE_DATAPATH_iv_0__15_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10256_));
OR2X2 OR2X2_3565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[15] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10257_));
OR2X2 OR2X2_3566 ( .A(AES_CORE_DATAPATH_iv_0__16_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10259_));
OR2X2 OR2X2_3567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[16] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10260_));
OR2X2 OR2X2_3568 ( .A(AES_CORE_DATAPATH_iv_0__17_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10262_));
OR2X2 OR2X2_3569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[17] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10263_));
OR2X2 OR2X2_357 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3176_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3177_));
OR2X2 OR2X2_3570 ( .A(AES_CORE_DATAPATH_iv_0__18_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10265_));
OR2X2 OR2X2_3571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[18] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10266_));
OR2X2 OR2X2_3572 ( .A(AES_CORE_DATAPATH_iv_0__19_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10268_));
OR2X2 OR2X2_3573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[19] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10269_));
OR2X2 OR2X2_3574 ( .A(AES_CORE_DATAPATH_iv_0__20_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10271_));
OR2X2 OR2X2_3575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[20] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10272_));
OR2X2 OR2X2_3576 ( .A(AES_CORE_DATAPATH_iv_0__21_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10274_));
OR2X2 OR2X2_3577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[21] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10275_));
OR2X2 OR2X2_3578 ( .A(AES_CORE_DATAPATH_iv_0__22_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10277_));
OR2X2 OR2X2_3579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[22] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10278_));
OR2X2 OR2X2_358 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3180_), .B(AES_CORE_DATAPATH__abc_16009_new_n3181_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3182_));
OR2X2 OR2X2_3580 ( .A(AES_CORE_DATAPATH_iv_0__23_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10280_));
OR2X2 OR2X2_3581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[23] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10281_));
OR2X2 OR2X2_3582 ( .A(AES_CORE_DATAPATH_iv_0__24_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10283_));
OR2X2 OR2X2_3583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[24] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10284_));
OR2X2 OR2X2_3584 ( .A(AES_CORE_DATAPATH_iv_0__25_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10286_));
OR2X2 OR2X2_3585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[25] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10287_));
OR2X2 OR2X2_3586 ( .A(AES_CORE_DATAPATH_iv_0__26_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10289_));
OR2X2 OR2X2_3587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[26] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10290_));
OR2X2 OR2X2_3588 ( .A(AES_CORE_DATAPATH_iv_0__27_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10292_));
OR2X2 OR2X2_3589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[27] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10293_));
OR2X2 OR2X2_359 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3182_), .B(AES_CORE_DATAPATH__abc_16009_new_n3179_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3183_));
OR2X2 OR2X2_3590 ( .A(AES_CORE_DATAPATH_iv_0__28_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10295_));
OR2X2 OR2X2_3591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[28] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10296_));
OR2X2 OR2X2_3592 ( .A(AES_CORE_DATAPATH_iv_0__29_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10298_));
OR2X2 OR2X2_3593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[29] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10299_));
OR2X2 OR2X2_3594 ( .A(AES_CORE_DATAPATH_iv_0__30_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10301_));
OR2X2 OR2X2_3595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[30] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10302_));
OR2X2 OR2X2_3596 ( .A(AES_CORE_DATAPATH_iv_0__31_), .B(\iv_en[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10304_));
OR2X2 OR2X2_3597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10211_), .B(\bus_in[31] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n10305_));
OR2X2 OR2X2_3598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10307_), .B(AES_CORE_DATAPATH__abc_16009_new_n10308_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10309_));
OR2X2 OR2X2_3599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10312_), .B(AES_CORE_DATAPATH__abc_16009_new_n10311_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__0_));
OR2X2 OR2X2_36 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n141_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n197_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n198_));
OR2X2 OR2X2_360 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3187_), .B(AES_CORE_DATAPATH__abc_16009_new_n3185_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3188_));
OR2X2 OR2X2_3600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10315_), .B(AES_CORE_DATAPATH__abc_16009_new_n10314_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__1_));
OR2X2 OR2X2_3601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10318_), .B(AES_CORE_DATAPATH__abc_16009_new_n10317_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__2_));
OR2X2 OR2X2_3602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10321_), .B(AES_CORE_DATAPATH__abc_16009_new_n10320_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__3_));
OR2X2 OR2X2_3603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10324_), .B(AES_CORE_DATAPATH__abc_16009_new_n10323_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__4_));
OR2X2 OR2X2_3604 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10327_), .B(AES_CORE_DATAPATH__abc_16009_new_n10326_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__5_));
OR2X2 OR2X2_3605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10330_), .B(AES_CORE_DATAPATH__abc_16009_new_n10329_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__6_));
OR2X2 OR2X2_3606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10333_), .B(AES_CORE_DATAPATH__abc_16009_new_n10332_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__7_));
OR2X2 OR2X2_3607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10336_), .B(AES_CORE_DATAPATH__abc_16009_new_n10335_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__8_));
OR2X2 OR2X2_3608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10339_), .B(AES_CORE_DATAPATH__abc_16009_new_n10338_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__9_));
OR2X2 OR2X2_3609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10342_), .B(AES_CORE_DATAPATH__abc_16009_new_n10341_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__10_));
OR2X2 OR2X2_361 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3188_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3189_));
OR2X2 OR2X2_3610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10345_), .B(AES_CORE_DATAPATH__abc_16009_new_n10344_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__11_));
OR2X2 OR2X2_3611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10348_), .B(AES_CORE_DATAPATH__abc_16009_new_n10347_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__12_));
OR2X2 OR2X2_3612 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10351_), .B(AES_CORE_DATAPATH__abc_16009_new_n10350_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__13_));
OR2X2 OR2X2_3613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10354_), .B(AES_CORE_DATAPATH__abc_16009_new_n10353_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__14_));
OR2X2 OR2X2_3614 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10357_), .B(AES_CORE_DATAPATH__abc_16009_new_n10356_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__15_));
OR2X2 OR2X2_3615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10360_), .B(AES_CORE_DATAPATH__abc_16009_new_n10359_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__16_));
OR2X2 OR2X2_3616 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10363_), .B(AES_CORE_DATAPATH__abc_16009_new_n10362_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__17_));
OR2X2 OR2X2_3617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10366_), .B(AES_CORE_DATAPATH__abc_16009_new_n10365_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__18_));
OR2X2 OR2X2_3618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10369_), .B(AES_CORE_DATAPATH__abc_16009_new_n10368_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__19_));
OR2X2 OR2X2_3619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10372_), .B(AES_CORE_DATAPATH__abc_16009_new_n10371_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__20_));
OR2X2 OR2X2_362 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3191_));
OR2X2 OR2X2_3620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10375_), .B(AES_CORE_DATAPATH__abc_16009_new_n10374_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__21_));
OR2X2 OR2X2_3621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10378_), .B(AES_CORE_DATAPATH__abc_16009_new_n10377_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__22_));
OR2X2 OR2X2_3622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10381_), .B(AES_CORE_DATAPATH__abc_16009_new_n10380_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__23_));
OR2X2 OR2X2_3623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10384_), .B(AES_CORE_DATAPATH__abc_16009_new_n10383_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__24_));
OR2X2 OR2X2_3624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10387_), .B(AES_CORE_DATAPATH__abc_16009_new_n10386_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__25_));
OR2X2 OR2X2_3625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10390_), .B(AES_CORE_DATAPATH__abc_16009_new_n10389_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__26_));
OR2X2 OR2X2_3626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10393_), .B(AES_CORE_DATAPATH__abc_16009_new_n10392_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__27_));
OR2X2 OR2X2_3627 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10396_), .B(AES_CORE_DATAPATH__abc_16009_new_n10395_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__28_));
OR2X2 OR2X2_3628 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10399_), .B(AES_CORE_DATAPATH__abc_16009_new_n10398_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__29_));
OR2X2 OR2X2_3629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10402_), .B(AES_CORE_DATAPATH__abc_16009_new_n10401_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__30_));
OR2X2 OR2X2_363 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3193_));
OR2X2 OR2X2_3630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10405_), .B(AES_CORE_DATAPATH__abc_16009_new_n10404_), .Y(AES_CORE_DATAPATH__0bkp_1_0__31_0__31_));
OR2X2 OR2X2_3631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7759_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10407_));
OR2X2 OR2X2_3632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10408_));
OR2X2 OR2X2_3633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10411_));
OR2X2 OR2X2_3634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10410_), .B(AES_CORE_DATAPATH__abc_16009_new_n10411_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10412_));
OR2X2 OR2X2_3635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10413_));
OR2X2 OR2X2_3636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7767_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10415_));
OR2X2 OR2X2_3637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10416_));
OR2X2 OR2X2_3638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8642_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10419_));
OR2X2 OR2X2_3639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10418_), .B(AES_CORE_DATAPATH__abc_16009_new_n10419_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10420_));
OR2X2 OR2X2_364 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3194_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3195_));
OR2X2 OR2X2_3640 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10421_));
OR2X2 OR2X2_3641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7775_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10423_));
OR2X2 OR2X2_3642 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10424_));
OR2X2 OR2X2_3643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8651_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10427_));
OR2X2 OR2X2_3644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10426_), .B(AES_CORE_DATAPATH__abc_16009_new_n10427_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10428_));
OR2X2 OR2X2_3645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10429_));
OR2X2 OR2X2_3646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7783_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10431_));
OR2X2 OR2X2_3647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10432_));
OR2X2 OR2X2_3648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8660_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10435_));
OR2X2 OR2X2_3649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10434_), .B(AES_CORE_DATAPATH__abc_16009_new_n10435_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10436_));
OR2X2 OR2X2_365 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3198_), .B(AES_CORE_DATAPATH__abc_16009_new_n3199_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3200_));
OR2X2 OR2X2_3650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10437_));
OR2X2 OR2X2_3651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7791_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10439_));
OR2X2 OR2X2_3652 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10440_));
OR2X2 OR2X2_3653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8669_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10443_));
OR2X2 OR2X2_3654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10442_), .B(AES_CORE_DATAPATH__abc_16009_new_n10443_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10444_));
OR2X2 OR2X2_3655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10445_));
OR2X2 OR2X2_3656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7799_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10447_));
OR2X2 OR2X2_3657 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10448_));
OR2X2 OR2X2_3658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8678_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10451_));
OR2X2 OR2X2_3659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10450_), .B(AES_CORE_DATAPATH__abc_16009_new_n10451_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10452_));
OR2X2 OR2X2_366 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3200_), .B(AES_CORE_DATAPATH__abc_16009_new_n3197_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3201_));
OR2X2 OR2X2_3660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10453_));
OR2X2 OR2X2_3661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7807_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10455_));
OR2X2 OR2X2_3662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10456_));
OR2X2 OR2X2_3663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8687_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10459_));
OR2X2 OR2X2_3664 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10458_), .B(AES_CORE_DATAPATH__abc_16009_new_n10459_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10460_));
OR2X2 OR2X2_3665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10461_));
OR2X2 OR2X2_3666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7815_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10463_));
OR2X2 OR2X2_3667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10464_));
OR2X2 OR2X2_3668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8696_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10467_));
OR2X2 OR2X2_3669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10466_), .B(AES_CORE_DATAPATH__abc_16009_new_n10467_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10468_));
OR2X2 OR2X2_367 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3205_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3206_));
OR2X2 OR2X2_3670 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10469_));
OR2X2 OR2X2_3671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7823_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10471_));
OR2X2 OR2X2_3672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10472_));
OR2X2 OR2X2_3673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8705_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10475_));
OR2X2 OR2X2_3674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10474_), .B(AES_CORE_DATAPATH__abc_16009_new_n10475_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10476_));
OR2X2 OR2X2_3675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__8_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10477_));
OR2X2 OR2X2_3676 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7831_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10479_));
OR2X2 OR2X2_3677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10480_));
OR2X2 OR2X2_3678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8714_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10483_));
OR2X2 OR2X2_3679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10482_), .B(AES_CORE_DATAPATH__abc_16009_new_n10483_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10484_));
OR2X2 OR2X2_368 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3206_), .B(AES_CORE_DATAPATH__abc_16009_new_n3203_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3207_));
OR2X2 OR2X2_3680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__9_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10485_));
OR2X2 OR2X2_3681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7839_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10487_));
OR2X2 OR2X2_3682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10488_));
OR2X2 OR2X2_3683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8723_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10491_));
OR2X2 OR2X2_3684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10490_), .B(AES_CORE_DATAPATH__abc_16009_new_n10491_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10492_));
OR2X2 OR2X2_3685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10493_));
OR2X2 OR2X2_3686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7847_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10495_));
OR2X2 OR2X2_3687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10496_));
OR2X2 OR2X2_3688 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8732_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10499_));
OR2X2 OR2X2_3689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10498_), .B(AES_CORE_DATAPATH__abc_16009_new_n10499_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10500_));
OR2X2 OR2X2_369 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3209_));
OR2X2 OR2X2_3690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10501_));
OR2X2 OR2X2_3691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7855_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10503_));
OR2X2 OR2X2_3692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10504_));
OR2X2 OR2X2_3693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8741_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10507_));
OR2X2 OR2X2_3694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10506_), .B(AES_CORE_DATAPATH__abc_16009_new_n10507_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10508_));
OR2X2 OR2X2_3695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10509_));
OR2X2 OR2X2_3696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7863_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10511_));
OR2X2 OR2X2_3697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10512_));
OR2X2 OR2X2_3698 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8750_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10515_));
OR2X2 OR2X2_3699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10514_), .B(AES_CORE_DATAPATH__abc_16009_new_n10515_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10516_));
OR2X2 OR2X2_37 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n198_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n200_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n201_));
OR2X2 OR2X2_370 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3211_));
OR2X2 OR2X2_3700 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10517_));
OR2X2 OR2X2_3701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7871_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10519_));
OR2X2 OR2X2_3702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10520_));
OR2X2 OR2X2_3703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8759_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10523_));
OR2X2 OR2X2_3704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10522_), .B(AES_CORE_DATAPATH__abc_16009_new_n10523_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10524_));
OR2X2 OR2X2_3705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__14_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10525_));
OR2X2 OR2X2_3706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7879_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10527_));
OR2X2 OR2X2_3707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10528_));
OR2X2 OR2X2_3708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8768_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10531_));
OR2X2 OR2X2_3709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10530_), .B(AES_CORE_DATAPATH__abc_16009_new_n10531_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10532_));
OR2X2 OR2X2_371 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3212_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3213_));
OR2X2 OR2X2_3710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__15_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10533_));
OR2X2 OR2X2_3711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7887_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10535_));
OR2X2 OR2X2_3712 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10536_));
OR2X2 OR2X2_3713 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8777_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10539_));
OR2X2 OR2X2_3714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10538_), .B(AES_CORE_DATAPATH__abc_16009_new_n10539_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10540_));
OR2X2 OR2X2_3715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10541_));
OR2X2 OR2X2_3716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7895_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10543_));
OR2X2 OR2X2_3717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10544_));
OR2X2 OR2X2_3718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8786_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10547_));
OR2X2 OR2X2_3719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10546_), .B(AES_CORE_DATAPATH__abc_16009_new_n10547_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10548_));
OR2X2 OR2X2_372 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3216_), .B(AES_CORE_DATAPATH__abc_16009_new_n3217_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3218_));
OR2X2 OR2X2_3720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10549_));
OR2X2 OR2X2_3721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7903_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10551_));
OR2X2 OR2X2_3722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10552_));
OR2X2 OR2X2_3723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8795_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10555_));
OR2X2 OR2X2_3724 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10554_), .B(AES_CORE_DATAPATH__abc_16009_new_n10555_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10556_));
OR2X2 OR2X2_3725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10557_));
OR2X2 OR2X2_3726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7911_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10559_));
OR2X2 OR2X2_3727 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10560_));
OR2X2 OR2X2_3728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8804_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10563_));
OR2X2 OR2X2_3729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10562_), .B(AES_CORE_DATAPATH__abc_16009_new_n10563_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10564_));
OR2X2 OR2X2_373 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3218_), .B(AES_CORE_DATAPATH__abc_16009_new_n3215_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3219_));
OR2X2 OR2X2_3730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__19_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10565_));
OR2X2 OR2X2_3731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7919_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10567_));
OR2X2 OR2X2_3732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10568_));
OR2X2 OR2X2_3733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8813_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10571_));
OR2X2 OR2X2_3734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10570_), .B(AES_CORE_DATAPATH__abc_16009_new_n10571_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10572_));
OR2X2 OR2X2_3735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__20_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10573_));
OR2X2 OR2X2_3736 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7927_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10575_));
OR2X2 OR2X2_3737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10576_));
OR2X2 OR2X2_3738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10579_));
OR2X2 OR2X2_3739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10578_), .B(AES_CORE_DATAPATH__abc_16009_new_n10579_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10580_));
OR2X2 OR2X2_374 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3223_), .B(AES_CORE_DATAPATH__abc_16009_new_n3221_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3224_));
OR2X2 OR2X2_3740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__21_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10581_));
OR2X2 OR2X2_3741 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7935_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10583_));
OR2X2 OR2X2_3742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10584_));
OR2X2 OR2X2_3743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8831_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10587_));
OR2X2 OR2X2_3744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10586_), .B(AES_CORE_DATAPATH__abc_16009_new_n10587_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10588_));
OR2X2 OR2X2_3745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10589_));
OR2X2 OR2X2_3746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7943_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10591_));
OR2X2 OR2X2_3747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10592_));
OR2X2 OR2X2_3748 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8840_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10595_));
OR2X2 OR2X2_3749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10594_), .B(AES_CORE_DATAPATH__abc_16009_new_n10595_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10596_));
OR2X2 OR2X2_375 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3224_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3225_));
OR2X2 OR2X2_3750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10597_));
OR2X2 OR2X2_3751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7951_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10599_));
OR2X2 OR2X2_3752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10600_));
OR2X2 OR2X2_3753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8849_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10603_));
OR2X2 OR2X2_3754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10602_), .B(AES_CORE_DATAPATH__abc_16009_new_n10603_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10604_));
OR2X2 OR2X2_3755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10605_));
OR2X2 OR2X2_3756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7959_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10607_));
OR2X2 OR2X2_3757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10608_));
OR2X2 OR2X2_3758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8858_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10611_));
OR2X2 OR2X2_3759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10610_), .B(AES_CORE_DATAPATH__abc_16009_new_n10611_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10612_));
OR2X2 OR2X2_376 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3227_));
OR2X2 OR2X2_3760 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10613_));
OR2X2 OR2X2_3761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7967_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10615_));
OR2X2 OR2X2_3762 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10616_));
OR2X2 OR2X2_3763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10619_));
OR2X2 OR2X2_3764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10618_), .B(AES_CORE_DATAPATH__abc_16009_new_n10619_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10620_));
OR2X2 OR2X2_3765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10621_));
OR2X2 OR2X2_3766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7975_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10623_));
OR2X2 OR2X2_3767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10624_));
OR2X2 OR2X2_3768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8876_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10627_));
OR2X2 OR2X2_3769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10626_), .B(AES_CORE_DATAPATH__abc_16009_new_n10627_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10628_));
OR2X2 OR2X2_377 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3229_));
OR2X2 OR2X2_3770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10629_));
OR2X2 OR2X2_3771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7983_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10631_));
OR2X2 OR2X2_3772 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10632_));
OR2X2 OR2X2_3773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8885_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10635_));
OR2X2 OR2X2_3774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10634_), .B(AES_CORE_DATAPATH__abc_16009_new_n10635_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10636_));
OR2X2 OR2X2_3775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10637_));
OR2X2 OR2X2_3776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7991_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10639_));
OR2X2 OR2X2_3777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10640_));
OR2X2 OR2X2_3778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8894_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10643_));
OR2X2 OR2X2_3779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10642_), .B(AES_CORE_DATAPATH__abc_16009_new_n10643_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10644_));
OR2X2 OR2X2_378 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3230_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3231_));
OR2X2 OR2X2_3780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10645_));
OR2X2 OR2X2_3781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n7999_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10647_));
OR2X2 OR2X2_3782 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10648_));
OR2X2 OR2X2_3783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8903_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10651_));
OR2X2 OR2X2_3784 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10650_), .B(AES_CORE_DATAPATH__abc_16009_new_n10651_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10652_));
OR2X2 OR2X2_3785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10653_));
OR2X2 OR2X2_3786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8007_), .B(AES_CORE_DATAPATH__abc_16009_new_n8628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10655_));
OR2X2 OR2X2_3787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n8527_), .B(AES_CORE_DATAPATH_bkp_1_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10656_));
OR2X2 OR2X2_3788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10310_), .B(AES_CORE_DATAPATH__abc_16009_new_n8912_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10659_));
OR2X2 OR2X2_3789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10658_), .B(AES_CORE_DATAPATH__abc_16009_new_n10659_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10660_));
OR2X2 OR2X2_379 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3234_), .B(AES_CORE_DATAPATH__abc_16009_new_n3235_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3236_));
OR2X2 OR2X2_3790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n10309_), .B(AES_CORE_DATAPATH_bkp_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10661_));
OR2X2 OR2X2_3791 ( .A(AES_CORE_CONTROL_UNIT_col_en_0_), .B(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_DATAPATH__abc_16009_new_n10663_));
OR2X2 OR2X2_3792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10664_));
OR2X2 OR2X2_3793 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10666_));
OR2X2 OR2X2_3794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10667_));
OR2X2 OR2X2_3795 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10669_));
OR2X2 OR2X2_3796 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10670_));
OR2X2 OR2X2_3797 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_CONTROL_UNIT_col_en_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10672_));
OR2X2 OR2X2_3798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10673_));
OR2X2 OR2X2_3799 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10675_));
OR2X2 OR2X2_38 ( .A(AES_CORE_CONTROL_UNIT_state_4_), .B(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_));
OR2X2 OR2X2_380 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3236_), .B(AES_CORE_DATAPATH__abc_16009_new_n3233_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3237_));
OR2X2 OR2X2_3800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10676_));
OR2X2 OR2X2_3801 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10678_));
OR2X2 OR2X2_3802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10679_));
OR2X2 OR2X2_3803 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10681_));
OR2X2 OR2X2_3804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10682_));
OR2X2 OR2X2_3805 ( .A(AES_CORE_CONTROL_UNIT_bypass_key_en), .B(AES_CORE_CONTROL_UNIT_key_en_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10684_));
OR2X2 OR2X2_3806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2807_), .B(AES_CORE_DATAPATH_key_en_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10685_));
OR2X2 OR2X2_3807 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10687_));
OR2X2 OR2X2_3808 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10688_));
OR2X2 OR2X2_3809 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10690_));
OR2X2 OR2X2_381 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3241_), .B(AES_CORE_DATAPATH__abc_16009_new_n3239_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3242_));
OR2X2 OR2X2_3810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10691_));
OR2X2 OR2X2_3811 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10693_));
OR2X2 OR2X2_3812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10694_));
OR2X2 OR2X2_3813 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp1_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10696_));
OR2X2 OR2X2_3814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2457_), .B(AES_CORE_DATAPATH_col_en_cnt_unit_pp2_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n10697_));
OR2X2 OR2X2_3815 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec));
OR2X2 OR2X2_3816 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n327_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n328_));
OR2X2 OR2X2_3817 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n329_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n330_));
OR2X2 OR2X2_3818 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n332_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n333_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n334_));
OR2X2 OR2X2_3819 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n331_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n335_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n336_));
OR2X2 OR2X2_382 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3242_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3243_));
OR2X2 OR2X2_3820 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n338_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n339_));
OR2X2 OR2X2_3821 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n340_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n341_));
OR2X2 OR2X2_3822 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n343_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n344_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n345_));
OR2X2 OR2X2_3823 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n342_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n346_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n347_));
OR2X2 OR2X2_3824 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n349_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n350_));
OR2X2 OR2X2_3825 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n351_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n352_));
OR2X2 OR2X2_3826 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n354_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n355_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n356_));
OR2X2 OR2X2_3827 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n353_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n357_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n358_));
OR2X2 OR2X2_3828 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n360_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n361_));
OR2X2 OR2X2_3829 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n362_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n363_));
OR2X2 OR2X2_383 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3245_));
OR2X2 OR2X2_3830 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n365_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n366_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n367_));
OR2X2 OR2X2_3831 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n364_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n368_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n369_));
OR2X2 OR2X2_3832 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n371_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n372_));
OR2X2 OR2X2_3833 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n373_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n374_));
OR2X2 OR2X2_3834 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n376_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n377_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n378_));
OR2X2 OR2X2_3835 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n375_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n379_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n380_));
OR2X2 OR2X2_3836 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n382_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n383_));
OR2X2 OR2X2_3837 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n384_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n385_));
OR2X2 OR2X2_3838 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n387_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n388_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n389_));
OR2X2 OR2X2_3839 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n386_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n390_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n391_));
OR2X2 OR2X2_384 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3247_));
OR2X2 OR2X2_3840 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n393_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n394_));
OR2X2 OR2X2_3841 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n395_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n396_));
OR2X2 OR2X2_3842 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n398_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n399_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n400_));
OR2X2 OR2X2_3843 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n397_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n401_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n402_));
OR2X2 OR2X2_3844 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n404_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n405_));
OR2X2 OR2X2_3845 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n406_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n407_));
OR2X2 OR2X2_3846 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n409_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n410_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n411_));
OR2X2 OR2X2_3847 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n408_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n412_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n413_));
OR2X2 OR2X2_3848 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n415_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n416_));
OR2X2 OR2X2_3849 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n417_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n418_));
OR2X2 OR2X2_385 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3248_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3249_));
OR2X2 OR2X2_3850 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n420_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n421_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n422_));
OR2X2 OR2X2_3851 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n419_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n423_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n424_));
OR2X2 OR2X2_3852 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n426_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n427_));
OR2X2 OR2X2_3853 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n428_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n429_));
OR2X2 OR2X2_3854 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n431_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n432_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n433_));
OR2X2 OR2X2_3855 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n430_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n434_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n435_));
OR2X2 OR2X2_3856 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n437_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n438_));
OR2X2 OR2X2_3857 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n439_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n440_));
OR2X2 OR2X2_3858 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n442_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n443_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n444_));
OR2X2 OR2X2_3859 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n441_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n445_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n446_));
OR2X2 OR2X2_386 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3252_), .B(AES_CORE_DATAPATH__abc_16009_new_n3253_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3254_));
OR2X2 OR2X2_3860 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n448_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n449_));
OR2X2 OR2X2_3861 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n450_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n451_));
OR2X2 OR2X2_3862 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n453_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n454_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n455_));
OR2X2 OR2X2_3863 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n452_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n456_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n457_));
OR2X2 OR2X2_3864 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n459_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n460_));
OR2X2 OR2X2_3865 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n461_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n462_));
OR2X2 OR2X2_3866 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n464_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n465_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n466_));
OR2X2 OR2X2_3867 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n463_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n467_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n468_));
OR2X2 OR2X2_3868 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n470_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n471_));
OR2X2 OR2X2_3869 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n472_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n473_));
OR2X2 OR2X2_387 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3254_), .B(AES_CORE_DATAPATH__abc_16009_new_n3251_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3255_));
OR2X2 OR2X2_3870 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n475_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n476_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n477_));
OR2X2 OR2X2_3871 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n474_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n478_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n479_));
OR2X2 OR2X2_3872 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n481_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n482_));
OR2X2 OR2X2_3873 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n483_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n484_));
OR2X2 OR2X2_3874 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n486_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n487_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n488_));
OR2X2 OR2X2_3875 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n485_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n489_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n490_));
OR2X2 OR2X2_3876 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n492_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n493_));
OR2X2 OR2X2_3877 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n494_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n495_));
OR2X2 OR2X2_3878 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n497_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n498_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n499_));
OR2X2 OR2X2_3879 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n496_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n500_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n501_));
OR2X2 OR2X2_388 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3259_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3260_));
OR2X2 OR2X2_3880 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n503_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n504_));
OR2X2 OR2X2_3881 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n505_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n506_));
OR2X2 OR2X2_3882 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n508_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n509_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n510_));
OR2X2 OR2X2_3883 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n507_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n511_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n512_));
OR2X2 OR2X2_3884 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n514_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n515_));
OR2X2 OR2X2_3885 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n516_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n517_));
OR2X2 OR2X2_3886 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n519_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n520_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n521_));
OR2X2 OR2X2_3887 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n518_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n522_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n523_));
OR2X2 OR2X2_3888 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n525_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n526_));
OR2X2 OR2X2_3889 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n527_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n528_));
OR2X2 OR2X2_389 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3260_), .B(AES_CORE_DATAPATH__abc_16009_new_n3257_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3261_));
OR2X2 OR2X2_3890 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n530_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n531_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n532_));
OR2X2 OR2X2_3891 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n529_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n533_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n534_));
OR2X2 OR2X2_3892 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n536_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n537_));
OR2X2 OR2X2_3893 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n538_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n539_));
OR2X2 OR2X2_3894 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n541_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n542_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n543_));
OR2X2 OR2X2_3895 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n540_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n544_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n545_));
OR2X2 OR2X2_3896 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n547_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n548_));
OR2X2 OR2X2_3897 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n549_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n550_));
OR2X2 OR2X2_3898 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n552_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n553_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n554_));
OR2X2 OR2X2_3899 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n551_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n555_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n556_));
OR2X2 OR2X2_39 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n203_));
OR2X2 OR2X2_390 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3265_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3266_));
OR2X2 OR2X2_3900 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n558_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n559_));
OR2X2 OR2X2_3901 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n560_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n561_));
OR2X2 OR2X2_3902 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n563_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n564_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n565_));
OR2X2 OR2X2_3903 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n562_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n566_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n567_));
OR2X2 OR2X2_3904 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n569_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n570_));
OR2X2 OR2X2_3905 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n571_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n572_));
OR2X2 OR2X2_3906 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n574_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n575_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n576_));
OR2X2 OR2X2_3907 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n573_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n577_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n578_));
OR2X2 OR2X2_3908 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n580_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n581_));
OR2X2 OR2X2_3909 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n582_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n583_));
OR2X2 OR2X2_391 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3269_), .B(AES_CORE_DATAPATH__abc_16009_new_n3270_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3271_));
OR2X2 OR2X2_3910 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n585_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n586_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n587_));
OR2X2 OR2X2_3911 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n584_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n588_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n589_));
OR2X2 OR2X2_3912 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n591_));
OR2X2 OR2X2_3913 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n599_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n601_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n602_));
OR2X2 OR2X2_3914 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n604_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n605_));
OR2X2 OR2X2_3915 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n603_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n606_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n607_));
OR2X2 OR2X2_3916 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n612_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n614_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_));
OR2X2 OR2X2_3917 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n616_));
OR2X2 OR2X2_3918 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n624_));
OR2X2 OR2X2_3919 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n626_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n627_));
OR2X2 OR2X2_392 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3271_), .B(AES_CORE_DATAPATH__abc_16009_new_n3268_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3272_));
OR2X2 OR2X2_3920 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n627_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n622_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n628_));
OR2X2 OR2X2_3921 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n632_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n633_));
OR2X2 OR2X2_3922 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n633_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n629_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n634_));
OR2X2 OR2X2_3923 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n635_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n621_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n637_));
OR2X2 OR2X2_3924 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n638_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n636_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n639_));
OR2X2 OR2X2_3925 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n644_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n645_));
OR2X2 OR2X2_3926 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n641_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n646_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_));
OR2X2 OR2X2_3927 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n648_));
OR2X2 OR2X2_3928 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n624_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n659_));
OR2X2 OR2X2_3929 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n660_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n599_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n661_));
OR2X2 OR2X2_393 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3273_));
OR2X2 OR2X2_3930 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_round_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_round_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n666_));
OR2X2 OR2X2_3931 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n666_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n655_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n667_));
OR2X2 OR2X2_3932 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n668_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n601_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n669_));
OR2X2 OR2X2_3933 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n662_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n670_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n671_));
OR2X2 OR2X2_3934 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n671_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n653_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n672_));
OR2X2 OR2X2_3935 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n673_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n657_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n674_));
OR2X2 OR2X2_3936 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n674_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n675_));
OR2X2 OR2X2_3937 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n677_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n678_));
OR2X2 OR2X2_3938 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n679_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n664_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n680_));
OR2X2 OR2X2_3939 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n681_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n682_));
OR2X2 OR2X2_394 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3275_), .B(AES_CORE_DATAPATH__abc_16009_new_n3264_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3276_));
OR2X2 OR2X2_3940 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n686_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n687_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n688_));
OR2X2 OR2X2_3941 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n688_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n689_));
OR2X2 OR2X2_3942 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n690_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n685_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_));
OR2X2 OR2X2_3943 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n692_));
OR2X2 OR2X2_3944 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n627_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n697_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n698_));
OR2X2 OR2X2_3945 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n633_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n699_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n700_));
OR2X2 OR2X2_3946 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n701_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n704_));
OR2X2 OR2X2_3947 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n708_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n702_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n709_));
OR2X2 OR2X2_3948 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n709_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n710_));
OR2X2 OR2X2_3949 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n711_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n707_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_));
OR2X2 OR2X2_395 ( .A(\key_out[24] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3277_));
OR2X2 OR2X2_3950 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n713_));
OR2X2 OR2X2_3951 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n720_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n723_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n724_));
OR2X2 OR2X2_3952 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n726_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n727_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n728_));
OR2X2 OR2X2_3953 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n731_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n733_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_));
OR2X2 OR2X2_3954 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n735_));
OR2X2 OR2X2_3955 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n741_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n742_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n743_));
OR2X2 OR2X2_3956 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n743_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n740_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n744_));
OR2X2 OR2X2_3957 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n673_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n721_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n745_));
OR2X2 OR2X2_3958 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n745_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n746_));
OR2X2 OR2X2_3959 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n679_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n718_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n747_));
OR2X2 OR2X2_396 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3279_), .B(AES_CORE_DATAPATH__abc_16009_new_n3263_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__24_));
OR2X2 OR2X2_3960 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n748_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n749_));
OR2X2 OR2X2_3961 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n753_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n754_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n755_));
OR2X2 OR2X2_3962 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n755_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n756_));
OR2X2 OR2X2_3963 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n757_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n752_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_93_));
OR2X2 OR2X2_3964 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n759_));
OR2X2 OR2X2_3965 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n699_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n764_));
OR2X2 OR2X2_3966 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n697_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n765_));
OR2X2 OR2X2_3967 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n766_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n769_));
OR2X2 OR2X2_3968 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n774_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n772_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_94_));
OR2X2 OR2X2_3969 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n776_));
OR2X2 OR2X2_397 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3281_));
OR2X2 OR2X2_3970 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n658_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n781_));
OR2X2 OR2X2_3971 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n665_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n782_));
OR2X2 OR2X2_3972 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n784_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n787_));
OR2X2 OR2X2_3973 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n791_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n785_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n792_));
OR2X2 OR2X2_3974 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n792_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n642_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n793_));
OR2X2 OR2X2_3975 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n794_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n790_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_95_));
OR2X2 OR2X2_3976 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n796_));
OR2X2 OR2X2_3977 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n800_));
OR2X2 OR2X2_3978 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n801_));
OR2X2 OR2X2_3979 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n803_));
OR2X2 OR2X2_398 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3283_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3284_));
OR2X2 OR2X2_3980 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n807_));
OR2X2 OR2X2_3981 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n808_));
OR2X2 OR2X2_3982 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n810_));
OR2X2 OR2X2_3983 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n814_));
OR2X2 OR2X2_3984 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n815_));
OR2X2 OR2X2_3985 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n817_));
OR2X2 OR2X2_3986 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n821_));
OR2X2 OR2X2_3987 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n822_));
OR2X2 OR2X2_3988 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n824_));
OR2X2 OR2X2_3989 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n828_));
OR2X2 OR2X2_399 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3287_), .B(AES_CORE_DATAPATH__abc_16009_new_n3288_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3289_));
OR2X2 OR2X2_3990 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n829_));
OR2X2 OR2X2_3991 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n831_));
OR2X2 OR2X2_3992 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n835_));
OR2X2 OR2X2_3993 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n836_));
OR2X2 OR2X2_3994 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n838_));
OR2X2 OR2X2_3995 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n842_));
OR2X2 OR2X2_3996 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n843_));
OR2X2 OR2X2_3997 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n845_));
OR2X2 OR2X2_3998 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n849_));
OR2X2 OR2X2_3999 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n850_));
OR2X2 OR2X2_4 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n108_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n106_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_));
OR2X2 OR2X2_40 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n201_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n203_), .Y(AES_CORE_CONTROL_UNIT_col_en_1_));
OR2X2 OR2X2_400 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3289_), .B(AES_CORE_DATAPATH__abc_16009_new_n3286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3290_));
OR2X2 OR2X2_4000 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n852_));
OR2X2 OR2X2_4001 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n856_));
OR2X2 OR2X2_4002 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n857_));
OR2X2 OR2X2_4003 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n859_));
OR2X2 OR2X2_4004 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n863_));
OR2X2 OR2X2_4005 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n864_));
OR2X2 OR2X2_4006 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n866_));
OR2X2 OR2X2_4007 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n870_));
OR2X2 OR2X2_4008 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n871_));
OR2X2 OR2X2_4009 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n873_));
OR2X2 OR2X2_401 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3291_));
OR2X2 OR2X2_4010 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n877_));
OR2X2 OR2X2_4011 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n878_));
OR2X2 OR2X2_4012 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n880_));
OR2X2 OR2X2_4013 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n884_));
OR2X2 OR2X2_4014 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n885_));
OR2X2 OR2X2_4015 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n887_));
OR2X2 OR2X2_4016 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n891_));
OR2X2 OR2X2_4017 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n892_));
OR2X2 OR2X2_4018 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n894_));
OR2X2 OR2X2_4019 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n898_));
OR2X2 OR2X2_402 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3295_), .B(AES_CORE_DATAPATH__abc_16009_new_n3293_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3296_));
OR2X2 OR2X2_4020 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n899_));
OR2X2 OR2X2_4021 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n901_));
OR2X2 OR2X2_4022 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n905_));
OR2X2 OR2X2_4023 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n906_));
OR2X2 OR2X2_4024 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n908_));
OR2X2 OR2X2_4025 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n912_));
OR2X2 OR2X2_4026 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n913_));
OR2X2 OR2X2_4027 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n915_));
OR2X2 OR2X2_4028 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n919_));
OR2X2 OR2X2_4029 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n920_));
OR2X2 OR2X2_403 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3296_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3297_));
OR2X2 OR2X2_4030 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n922_));
OR2X2 OR2X2_4031 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n926_));
OR2X2 OR2X2_4032 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n927_));
OR2X2 OR2X2_4033 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n929_));
OR2X2 OR2X2_4034 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n933_));
OR2X2 OR2X2_4035 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n934_));
OR2X2 OR2X2_4036 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n936_));
OR2X2 OR2X2_4037 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n940_));
OR2X2 OR2X2_4038 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n941_));
OR2X2 OR2X2_4039 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n943_));
OR2X2 OR2X2_404 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3299_));
OR2X2 OR2X2_4040 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n947_));
OR2X2 OR2X2_4041 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n948_));
OR2X2 OR2X2_4042 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n950_));
OR2X2 OR2X2_4043 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n954_));
OR2X2 OR2X2_4044 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n955_));
OR2X2 OR2X2_4045 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n957_));
OR2X2 OR2X2_4046 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n961_));
OR2X2 OR2X2_4047 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n962_));
OR2X2 OR2X2_4048 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n964_));
OR2X2 OR2X2_4049 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n968_));
OR2X2 OR2X2_405 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3301_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3302_));
OR2X2 OR2X2_4050 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n969_));
OR2X2 OR2X2_4051 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n971_));
OR2X2 OR2X2_4052 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n975_));
OR2X2 OR2X2_4053 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n976_));
OR2X2 OR2X2_4054 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n978_));
OR2X2 OR2X2_4055 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n982_));
OR2X2 OR2X2_4056 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n983_));
OR2X2 OR2X2_4057 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n985_));
OR2X2 OR2X2_4058 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n989_));
OR2X2 OR2X2_4059 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n990_));
OR2X2 OR2X2_406 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3305_), .B(AES_CORE_DATAPATH__abc_16009_new_n3306_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3307_));
OR2X2 OR2X2_4060 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n992_));
OR2X2 OR2X2_4061 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n996_));
OR2X2 OR2X2_4062 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n997_));
OR2X2 OR2X2_4063 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n999_));
OR2X2 OR2X2_4064 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1003_));
OR2X2 OR2X2_4065 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1004_));
OR2X2 OR2X2_4066 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1006_));
OR2X2 OR2X2_4067 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1010_));
OR2X2 OR2X2_4068 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1011_));
OR2X2 OR2X2_4069 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1013_));
OR2X2 OR2X2_407 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3307_), .B(AES_CORE_DATAPATH__abc_16009_new_n3304_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3308_));
OR2X2 OR2X2_4070 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1017_));
OR2X2 OR2X2_4071 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n598_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_3__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1018_));
OR2X2 OR2X2_4072 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1020_));
OR2X2 OR2X2_4073 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1024_));
OR2X2 OR2X2_4074 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1028_));
OR2X2 OR2X2_4075 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1032_));
OR2X2 OR2X2_4076 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1036_));
OR2X2 OR2X2_4077 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1040_));
OR2X2 OR2X2_4078 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1044_));
OR2X2 OR2X2_4079 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1048_));
OR2X2 OR2X2_408 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3309_));
OR2X2 OR2X2_4080 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1052_));
OR2X2 OR2X2_4081 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1056_));
OR2X2 OR2X2_4082 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1060_));
OR2X2 OR2X2_4083 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1064_));
OR2X2 OR2X2_4084 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1068_));
OR2X2 OR2X2_4085 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1072_));
OR2X2 OR2X2_4086 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1076_));
OR2X2 OR2X2_4087 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1080_));
OR2X2 OR2X2_4088 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1084_));
OR2X2 OR2X2_4089 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1088_));
OR2X2 OR2X2_409 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3313_), .B(AES_CORE_DATAPATH__abc_16009_new_n3311_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3314_));
OR2X2 OR2X2_4090 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1092_));
OR2X2 OR2X2_4091 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1096_));
OR2X2 OR2X2_4092 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1100_));
OR2X2 OR2X2_4093 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1104_));
OR2X2 OR2X2_4094 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1108_));
OR2X2 OR2X2_4095 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1112_));
OR2X2 OR2X2_4096 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1117_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1118_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_120_));
OR2X2 OR2X2_4097 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n644_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1120_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1121_));
OR2X2 OR2X2_4098 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n639_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1122_));
OR2X2 OR2X2_4099 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n688_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1124_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1125_));
OR2X2 OR2X2_41 ( .A(AES_CORE_CONTROL_UNIT_state_12_), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n205_));
OR2X2 OR2X2_410 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3314_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3315_));
OR2X2 OR2X2_4100 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n683_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1126_));
OR2X2 OR2X2_4101 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n709_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1128_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1129_));
OR2X2 OR2X2_4102 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n705_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1130_));
OR2X2 OR2X2_4103 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1135_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1133_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_124_));
OR2X2 OR2X2_4104 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n755_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1137_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1138_));
OR2X2 OR2X2_4105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n750_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1139_));
OR2X2 OR2X2_4106 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n770_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1141_));
OR2X2 OR2X2_4107 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1143_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1142_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1144_));
OR2X2 OR2X2_4108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n788_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1146_));
OR2X2 OR2X2_4109 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n792_), .B(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1147_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1148_));
OR2X2 OR2X2_411 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3317_));
OR2X2 OR2X2_4110 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__0_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1150_));
OR2X2 OR2X2_4111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__1_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__1_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1154_));
OR2X2 OR2X2_4112 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__2_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__2_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1158_));
OR2X2 OR2X2_4113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__3_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__3_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1162_));
OR2X2 OR2X2_4114 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__4_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1166_));
OR2X2 OR2X2_4115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__5_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__5_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1170_));
OR2X2 OR2X2_4116 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__6_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__6_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1174_));
OR2X2 OR2X2_4117 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__7_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1178_));
OR2X2 OR2X2_4118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__8_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__8_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1182_));
OR2X2 OR2X2_4119 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__9_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__9_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1186_));
OR2X2 OR2X2_412 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3319_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3320_));
OR2X2 OR2X2_4120 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__10_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1190_));
OR2X2 OR2X2_4121 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__11_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1194_));
OR2X2 OR2X2_4122 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__12_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1198_));
OR2X2 OR2X2_4123 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__13_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1202_));
OR2X2 OR2X2_4124 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__14_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__14_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1206_));
OR2X2 OR2X2_4125 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__15_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__15_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1210_));
OR2X2 OR2X2_4126 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__16_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1214_));
OR2X2 OR2X2_4127 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__17_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1218_));
OR2X2 OR2X2_4128 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__18_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1222_));
OR2X2 OR2X2_4129 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__19_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__19_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1226_));
OR2X2 OR2X2_413 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3323_), .B(AES_CORE_DATAPATH__abc_16009_new_n3324_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3325_));
OR2X2 OR2X2_4130 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__20_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1230_));
OR2X2 OR2X2_4131 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__21_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__21_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1234_));
OR2X2 OR2X2_4132 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__22_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1238_));
OR2X2 OR2X2_4133 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__23_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__23_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1242_));
OR2X2 OR2X2_4134 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__24_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1246_));
OR2X2 OR2X2_4135 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__25_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__25_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1250_));
OR2X2 OR2X2_4136 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__26_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1254_));
OR2X2 OR2X2_4137 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__27_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__27_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1258_));
OR2X2 OR2X2_4138 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__28_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1262_));
OR2X2 OR2X2_4139 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__29_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__29_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1266_));
OR2X2 OR2X2_414 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3325_), .B(AES_CORE_DATAPATH__abc_16009_new_n3322_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3326_));
OR2X2 OR2X2_4140 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__30_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__30_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1270_));
OR2X2 OR2X2_4141 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__31_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_2__31_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER__abc_24255_new_n1274_));
OR2X2 OR2X2_4142 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n99_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n100_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n101_));
OR2X2 OR2X2_4143 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n102_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n103_));
OR2X2 OR2X2_4144 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n104_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n105_));
OR2X2 OR2X2_4145 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n108_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n110_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n111_));
OR2X2 OR2X2_4146 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n111_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n101_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n112_));
OR2X2 OR2X2_4147 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n113_));
OR2X2 OR2X2_4148 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n116_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n115_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n117_));
OR2X2 OR2X2_4149 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n122_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n123_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_));
OR2X2 OR2X2_415 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__27_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3327_));
OR2X2 OR2X2_4150 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n125_));
OR2X2 OR2X2_4151 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n129_));
OR2X2 OR2X2_4152 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n128_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n133_));
OR2X2 OR2X2_4153 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n136_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n126_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n137_));
OR2X2 OR2X2_4154 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n140_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n130_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_));
OR2X2 OR2X2_4155 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n137_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n142_));
OR2X2 OR2X2_4156 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n144_));
OR2X2 OR2X2_4157 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n145_));
OR2X2 OR2X2_4158 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n148_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n149_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_));
OR2X2 OR2X2_4159 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n151_));
OR2X2 OR2X2_416 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3331_), .B(AES_CORE_DATAPATH__abc_16009_new_n3329_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3332_));
OR2X2 OR2X2_4160 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n119_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n153_));
OR2X2 OR2X2_4161 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n154_));
OR2X2 OR2X2_4162 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n155_));
OR2X2 OR2X2_4163 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_0_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n157_));
OR2X2 OR2X2_4164 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n98_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n159_));
OR2X2 OR2X2_4165 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n161_));
OR2X2 OR2X2_4166 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n162_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n165_));
OR2X2 OR2X2_4167 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n168_));
OR2X2 OR2X2_4168 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n176_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n169_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n177_));
OR2X2 OR2X2_4169 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n178_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n172_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n179_));
OR2X2 OR2X2_417 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3332_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3333_));
OR2X2 OR2X2_4170 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n181_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n182_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n183_));
OR2X2 OR2X2_4171 ( .A(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n185_));
OR2X2 OR2X2_4172 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n191_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n186_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_));
OR2X2 OR2X2_4173 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n189_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n193_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_));
OR2X2 OR2X2_4174 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n197_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n198_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_));
OR2X2 OR2X2_4175 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n152_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n200_));
OR2X2 OR2X2_4176 ( .A(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n201_));
OR2X2 OR2X2_4177 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n156_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n204_));
OR2X2 OR2X2_4178 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n205_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n206_));
OR2X2 OR2X2_4179 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n207_));
OR2X2 OR2X2_418 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3337_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3338_));
OR2X2 OR2X2_4180 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n208_));
OR2X2 OR2X2_4181 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n210_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n211_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n212_));
OR2X2 OR2X2_4182 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n212_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n213_));
OR2X2 OR2X2_4183 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n214_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n215_));
OR2X2 OR2X2_4184 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n212_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n216_));
OR2X2 OR2X2_4185 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n205_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n217_));
OR2X2 OR2X2_4186 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n218_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n183_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n219_));
OR2X2 OR2X2_4187 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n175_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n221_));
OR2X2 OR2X2_4188 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n222_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n223_));
OR2X2 OR2X2_4189 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n224_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n227_));
OR2X2 OR2X2_419 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3341_), .B(AES_CORE_DATAPATH__abc_16009_new_n3342_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3343_));
OR2X2 OR2X2_4190 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n231_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n233_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n234_));
OR2X2 OR2X2_4191 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n236_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n237_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_));
OR2X2 OR2X2_4192 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__0_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n239_));
OR2X2 OR2X2_4193 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n192_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n242_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n243_));
OR2X2 OR2X2_4194 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n244_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n240_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n245_));
OR2X2 OR2X2_4195 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n245_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n188_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n246_));
OR2X2 OR2X2_4196 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n249_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n250_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_));
OR2X2 OR2X2_4197 ( .A(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n253_));
OR2X2 OR2X2_4198 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n252_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n256_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n257_));
OR2X2 OR2X2_4199 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n259_));
OR2X2 OR2X2_42 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n143_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n205_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n206_));
OR2X2 OR2X2_420 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3343_), .B(AES_CORE_DATAPATH__abc_16009_new_n3340_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3344_));
OR2X2 OR2X2_4200 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n260_));
OR2X2 OR2X2_4201 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n258_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n262_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n263_));
OR2X2 OR2X2_4202 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n264_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n247_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n265_));
OR2X2 OR2X2_4203 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n266_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n267_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n268_));
OR2X2 OR2X2_4204 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n263_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n268_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n269_));
OR2X2 OR2X2_4205 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n271_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n272_));
OR2X2 OR2X2_4206 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n270_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n273_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n274_));
OR2X2 OR2X2_4207 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n230_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n276_));
OR2X2 OR2X2_4208 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n277_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n278_));
OR2X2 OR2X2_4209 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n279_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n282_));
OR2X2 OR2X2_421 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__28_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3345_));
OR2X2 OR2X2_4210 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n286_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n288_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n289_));
OR2X2 OR2X2_4211 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n293_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n290_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n294_));
OR2X2 OR2X2_4212 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n296_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n297_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n298_));
OR2X2 OR2X2_4213 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n101_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n300_));
OR2X2 OR2X2_4214 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n115_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n301_));
OR2X2 OR2X2_4215 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n247_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n303_));
OR2X2 OR2X2_4216 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n304_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n305_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n306_));
OR2X2 OR2X2_4217 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n268_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n306_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n307_));
OR2X2 OR2X2_4218 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n308_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n309_));
OR2X2 OR2X2_4219 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n310_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n311_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n312_));
OR2X2 OR2X2_422 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3347_), .B(AES_CORE_DATAPATH__abc_16009_new_n3336_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3348_));
OR2X2 OR2X2_4220 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n312_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n313_));
OR2X2 OR2X2_4221 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__1_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n315_));
OR2X2 OR2X2_4222 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n318_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n319_));
OR2X2 OR2X2_4223 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n320_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n316_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n321_));
OR2X2 OR2X2_4224 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n321_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n322_));
OR2X2 OR2X2_4225 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n314_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n323_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n324_));
OR2X2 OR2X2_4226 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n312_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n325_));
OR2X2 OR2X2_4227 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n308_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n326_));
OR2X2 OR2X2_4228 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n328_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n329_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n330_));
OR2X2 OR2X2_4229 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n330_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n331_));
OR2X2 OR2X2_423 ( .A(\key_out[28] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_4_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3349_));
OR2X2 OR2X2_4230 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n332_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n333_));
OR2X2 OR2X2_4231 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n314_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n330_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n334_));
OR2X2 OR2X2_4232 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n323_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n335_));
OR2X2 OR2X2_4233 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n336_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n298_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n337_));
OR2X2 OR2X2_4234 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n339_));
OR2X2 OR2X2_4235 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n340_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n341_));
OR2X2 OR2X2_4236 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n107_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n342_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n345_));
OR2X2 OR2X2_4237 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n348_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n349_));
OR2X2 OR2X2_4238 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n350_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n351_));
OR2X2 OR2X2_4239 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n354_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n356_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n357_));
OR2X2 OR2X2_424 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3351_), .B(AES_CORE_DATAPATH__abc_16009_new_n3335_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__28_));
OR2X2 OR2X2_4240 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n359_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n360_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n361_));
OR2X2 OR2X2_4241 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n363_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n365_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n366_));
OR2X2 OR2X2_4242 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n366_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n367_));
OR2X2 OR2X2_4243 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n368_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n369_));
OR2X2 OR2X2_4244 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n372_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n371_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n373_));
OR2X2 OR2X2_4245 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n177_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n375_));
OR2X2 OR2X2_4246 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n171_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n376_));
OR2X2 OR2X2_4247 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n378_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n374_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n379_));
OR2X2 OR2X2_4248 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n379_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n380_));
OR2X2 OR2X2_4249 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n323_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n377_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n381_));
OR2X2 OR2X2_425 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3355_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3356_));
OR2X2 OR2X2_4250 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n330_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n373_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n382_));
OR2X2 OR2X2_4251 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n383_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n384_));
OR2X2 OR2X2_4252 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n385_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n370_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n386_));
OR2X2 OR2X2_4253 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n209_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n368_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n387_));
OR2X2 OR2X2_4254 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n194_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n366_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n388_));
OR2X2 OR2X2_4255 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n383_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n390_));
OR2X2 OR2X2_4256 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n379_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n391_));
OR2X2 OR2X2_4257 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n392_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n389_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n393_));
OR2X2 OR2X2_4258 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n394_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n361_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n395_));
OR2X2 OR2X2_4259 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n392_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n370_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n396_));
OR2X2 OR2X2_426 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3359_), .B(AES_CORE_DATAPATH__abc_16009_new_n3360_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3361_));
OR2X2 OR2X2_4260 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n385_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n389_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n397_));
OR2X2 OR2X2_4261 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n398_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n399_));
OR2X2 OR2X2_4262 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n402_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n401_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n403_));
OR2X2 OR2X2_4263 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n406_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n407_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n408_));
OR2X2 OR2X2_4264 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n410_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n411_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n412_));
OR2X2 OR2X2_4265 ( .A(AES_CORE_DATAPATH_MIX_COL_col_2__3_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n414_));
OR2X2 OR2X2_4266 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n419_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n420_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n421_));
OR2X2 OR2X2_4267 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n261_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n235_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n422_));
OR2X2 OR2X2_4268 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n257_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n234_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n423_));
OR2X2 OR2X2_4269 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n389_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n424_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n425_));
OR2X2 OR2X2_427 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3361_), .B(AES_CORE_DATAPATH__abc_16009_new_n3358_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3362_));
OR2X2 OR2X2_4270 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n426_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n427_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n428_));
OR2X2 OR2X2_4271 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n428_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n370_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n429_));
OR2X2 OR2X2_4272 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n430_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n421_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n431_));
OR2X2 OR2X2_4273 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n433_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n434_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n435_));
OR2X2 OR2X2_4274 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n435_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n432_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n436_));
OR2X2 OR2X2_4275 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n437_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n438_));
OR2X2 OR2X2_4276 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n439_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n440_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n441_));
OR2X2 OR2X2_4277 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n441_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n412_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n442_));
OR2X2 OR2X2_4278 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n139_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n444_));
OR2X2 OR2X2_4279 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n134_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n445_));
OR2X2 OR2X2_428 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__29_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3363_));
OR2X2 OR2X2_4280 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n446_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n449_));
OR2X2 OR2X2_4281 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n121_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n451_));
OR2X2 OR2X2_4282 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n196_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n452_));
OR2X2 OR2X2_4283 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n450_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n453_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n454_));
OR2X2 OR2X2_4284 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n455_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n456_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n457_));
OR2X2 OR2X2_4285 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n460_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n461_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_));
OR2X2 OR2X2_4286 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n464_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n463_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n465_));
OR2X2 OR2X2_4287 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n466_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n432_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n467_));
OR2X2 OR2X2_4288 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n465_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n421_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n468_));
OR2X2 OR2X2_4289 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n469_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n462_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n470_));
OR2X2 OR2X2_429 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3365_), .B(AES_CORE_DATAPATH__abc_16009_new_n3354_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3366_));
OR2X2 OR2X2_4290 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n472_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n471_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n473_));
OR2X2 OR2X2_4291 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n476_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n477_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_6_));
OR2X2 OR2X2_4292 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n120_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n479_));
OR2X2 OR2X2_4293 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n196_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n480_));
OR2X2 OR2X2_4294 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n483_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n484_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n485_));
OR2X2 OR2X2_4295 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n485_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n251_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n486_));
OR2X2 OR2X2_4296 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n487_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n255_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n488_));
OR2X2 OR2X2_4297 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n491_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n492_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n493_));
OR2X2 OR2X2_4298 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n494_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n128_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n495_));
OR2X2 OR2X2_4299 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n493_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n137_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n496_));
OR2X2 OR2X2_43 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n201_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n206_), .Y(AES_CORE_CONTROL_UNIT_col_en_2_));
OR2X2 OR2X2_430 ( .A(\key_out[29] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_5_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3367_));
OR2X2 OR2X2_4300 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n490_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n497_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n498_));
OR2X2 OR2X2_4301 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n499_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n500_));
OR2X2 OR2X2_4302 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n104_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n502_));
OR2X2 OR2X2_4303 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n248_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n503_));
OR2X2 OR2X2_4304 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n505_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n506_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n507_));
OR2X2 OR2X2_4305 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n508_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n504_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n509_));
OR2X2 OR2X2_4306 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n507_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n510_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n511_));
OR2X2 OR2X2_4307 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n143_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n199_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n514_));
OR2X2 OR2X2_4308 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n150_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n203_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n515_));
OR2X2 OR2X2_4309 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n518_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n519_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_8_));
OR2X2 OR2X2_431 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3369_), .B(AES_CORE_DATAPATH__abc_16009_new_n3353_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__29_));
OR2X2 OR2X2_4310 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n97_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n521_));
OR2X2 OR2X2_4311 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n160_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__0_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n522_));
OR2X2 OR2X2_4312 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n525_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n526_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n527_));
OR2X2 OR2X2_4313 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n528_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n529_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n530_));
OR2X2 OR2X2_4314 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n527_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n531_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n534_));
OR2X2 OR2X2_4315 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n537_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n538_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n539_));
OR2X2 OR2X2_4316 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n542_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n540_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_9_));
OR2X2 OR2X2_4317 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n174_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n544_));
OR2X2 OR2X2_4318 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n222_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n545_));
OR2X2 OR2X2_4319 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n547_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n548_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n549_));
OR2X2 OR2X2_432 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3373_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3374_));
OR2X2 OR2X2_4320 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n550_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n546_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n551_));
OR2X2 OR2X2_4321 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n549_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n552_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n553_));
OR2X2 OR2X2_4322 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n264_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n302_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n556_));
OR2X2 OR2X2_4323 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n263_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n306_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n557_));
OR2X2 OR2X2_4324 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n558_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n555_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n559_));
OR2X2 OR2X2_4325 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n560_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_10_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n561_));
OR2X2 OR2X2_4326 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n563_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n564_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n565_));
OR2X2 OR2X2_4327 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n232_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n567_));
OR2X2 OR2X2_4328 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n277_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n568_));
OR2X2 OR2X2_4329 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n571_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n572_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n573_));
OR2X2 OR2X2_433 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3377_), .B(AES_CORE_DATAPATH__abc_16009_new_n3378_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3379_));
OR2X2 OR2X2_4330 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n575_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n576_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_11_));
OR2X2 OR2X2_4331 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n578_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n579_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n580_));
OR2X2 OR2X2_4332 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n314_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n377_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n583_));
OR2X2 OR2X2_4333 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n327_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n373_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n584_));
OR2X2 OR2X2_4334 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n581_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n586_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_11_));
OR2X2 OR2X2_4335 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n589_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n588_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n590_));
OR2X2 OR2X2_4336 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n287_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n592_));
OR2X2 OR2X2_4337 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n340_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n593_));
OR2X2 OR2X2_4338 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n596_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n597_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n598_));
OR2X2 OR2X2_4339 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n600_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n601_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_));
OR2X2 OR2X2_434 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3379_), .B(AES_CORE_DATAPATH__abc_16009_new_n3376_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3380_));
OR2X2 OR2X2_4340 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n385_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n424_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n603_));
OR2X2 OR2X2_4341 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n392_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n428_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n604_));
OR2X2 OR2X2_4342 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n605_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_12_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n606_));
OR2X2 OR2X2_4343 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n385_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n428_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n608_));
OR2X2 OR2X2_4344 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n392_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n424_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n609_));
OR2X2 OR2X2_4345 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n610_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n607_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n611_));
OR2X2 OR2X2_4346 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n348_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n613_));
OR2X2 OR2X2_4347 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n405_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__4_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n614_));
OR2X2 OR2X2_4348 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n616_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n617_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n618_));
OR2X2 OR2X2_4349 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n619_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n615_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n620_));
OR2X2 OR2X2_435 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__30_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3381_));
OR2X2 OR2X2_4350 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n618_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n621_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n622_));
OR2X2 OR2X2_4351 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n430_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n466_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n625_));
OR2X2 OR2X2_4352 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n435_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n465_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n626_));
OR2X2 OR2X2_4353 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n627_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n624_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n628_));
OR2X2 OR2X2_4354 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n435_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n466_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n629_));
OR2X2 OR2X2_4355 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n430_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n465_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n630_));
OR2X2 OR2X2_4356 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n631_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_13_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n632_));
OR2X2 OR2X2_4357 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n138_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n634_));
OR2X2 OR2X2_4358 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n134_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n635_));
OR2X2 OR2X2_4359 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n639_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n638_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n640_));
OR2X2 OR2X2_436 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3383_), .B(AES_CORE_DATAPATH__abc_16009_new_n3372_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3384_));
OR2X2 OR2X2_4360 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n642_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n643_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n644_));
OR2X2 OR2X2_4361 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n469_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n352_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n646_));
OR2X2 OR2X2_4362 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n472_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n353_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n647_));
OR2X2 OR2X2_4363 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n648_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n644_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n649_));
OR2X2 OR2X2_4364 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n650_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_14_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n651_));
OR2X2 OR2X2_4365 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n120_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n653_));
OR2X2 OR2X2_4366 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n195_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__6_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n654_));
OR2X2 OR2X2_4367 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n102_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n656_));
OR2X2 OR2X2_4368 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n190_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__7_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n657_));
OR2X2 OR2X2_4369 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n660_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n661_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n662_));
OR2X2 OR2X2_437 ( .A(\key_out[30] ), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_6_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3385_));
OR2X2 OR2X2_4370 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n663_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n655_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n664_));
OR2X2 OR2X2_4371 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n662_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n665_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n666_));
OR2X2 OR2X2_4372 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n494_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n669_));
OR2X2 OR2X2_4373 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n493_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n670_));
OR2X2 OR2X2_4374 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n671_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n667_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n672_));
OR2X2 OR2X2_4375 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n673_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_15_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n674_));
OR2X2 OR2X2_4376 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n676_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n677_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n678_));
OR2X2 OR2X2_4377 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n680_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n679_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n681_));
OR2X2 OR2X2_4378 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n683_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n685_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_16_));
OR2X2 OR2X2_4379 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n688_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n689_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_16_));
OR2X2 OR2X2_438 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3387_), .B(AES_CORE_DATAPATH__abc_16009_new_n3371_), .Y(AES_CORE_DATAPATH__0sbox_pp2_31_0__30_));
OR2X2 OR2X2_4380 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n691_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n692_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n693_));
OR2X2 OR2X2_4381 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n695_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n696_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n697_));
OR2X2 OR2X2_4382 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n699_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n700_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n701_));
OR2X2 OR2X2_4383 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n703_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n704_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n705_));
OR2X2 OR2X2_4384 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n214_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_17_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n707_));
OR2X2 OR2X2_4385 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n218_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n705_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n708_));
OR2X2 OR2X2_4386 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n710_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n711_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n712_));
OR2X2 OR2X2_4387 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n713_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n714_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n715_));
OR2X2 OR2X2_4388 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n715_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n712_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n716_));
OR2X2 OR2X2_4389 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n718_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n717_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n719_));
OR2X2 OR2X2_439 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2803_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3389_));
OR2X2 OR2X2_4390 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n270_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n721_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n722_));
OR2X2 OR2X2_4391 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n271_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_18_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n723_));
OR2X2 OR2X2_4392 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n725_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n726_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n727_));
OR2X2 OR2X2_4393 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n728_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n730_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n731_));
OR2X2 OR2X2_4394 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n594_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n285_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n732_));
OR2X2 OR2X2_4395 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n595_), .B(AES_CORE_DATAPATH_MIX_COL_col_3__3_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n733_));
OR2X2 OR2X2_4396 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n731_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n734_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n737_));
OR2X2 OR2X2_4397 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n332_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_19_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n739_));
OR2X2 OR2X2_4398 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n336_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n740_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n741_));
OR2X2 OR2X2_4399 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n743_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n744_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n745_));
OR2X2 OR2X2_44 ( .A(AES_CORE_CONTROL_UNIT_state_9_), .B(AES_CORE_CONTROL_UNIT_state_2_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_));
OR2X2 OR2X2_440 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2822_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_0__31_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3391_));
OR2X2 OR2X2_4400 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n684_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n745_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n748_));
OR2X2 OR2X2_4401 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n751_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n752_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n753_));
OR2X2 OR2X2_4402 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n755_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n756_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n757_));
OR2X2 OR2X2_4403 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n394_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n757_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n759_));
OR2X2 OR2X2_4404 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n398_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_20_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n760_));
OR2X2 OR2X2_4405 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n762_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n763_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n764_));
OR2X2 OR2X2_4406 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n764_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n767_));
OR2X2 OR2X2_4407 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n768_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n132_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n769_));
OR2X2 OR2X2_4408 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n770_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n141_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n771_));
OR2X2 OR2X2_4409 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n437_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_21_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n774_));
OR2X2 OR2X2_441 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2821_), .B(AES_CORE_DATAPATH__abc_16009_new_n3392_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3393_));
OR2X2 OR2X2_4410 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n441_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n772_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n775_));
OR2X2 OR2X2_4411 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n138_), .B(AES_CORE_DATAPATH_MIX_COL_col_2__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n777_));
OR2X2 OR2X2_4412 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n135_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__5_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n778_));
OR2X2 OR2X2_4413 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n781_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n782_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n783_));
OR2X2 OR2X2_4414 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n785_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n786_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_22_));
OR2X2 OR2X2_4415 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n789_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n790_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_22_));
OR2X2 OR2X2_4416 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n792_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n793_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n794_));
OR2X2 OR2X2_4417 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n795_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n796_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n797_));
OR2X2 OR2X2_4418 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n798_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n794_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n801_));
OR2X2 OR2X2_4419 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n802_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n497_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n804_));
OR2X2 OR2X2_442 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3396_), .B(AES_CORE_DATAPATH__abc_16009_new_n3397_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3398_));
OR2X2 OR2X2_4420 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_23_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n499_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n805_));
OR2X2 OR2X2_4421 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n807_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n808_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n809_));
OR2X2 OR2X2_4422 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n811_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n812_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_24_));
OR2X2 OR2X2_4423 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n815_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n816_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_24_));
OR2X2 OR2X2_4424 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n818_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n819_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n820_));
OR2X2 OR2X2_4425 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n820_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n823_));
OR2X2 OR2X2_4426 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n318_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n174_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n826_));
OR2X2 OR2X2_4427 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n321_), .B(AES_CORE_DATAPATH_MIX_COL_col_1__1_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n827_));
OR2X2 OR2X2_4428 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n825_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n828_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n831_));
OR2X2 OR2X2_4429 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n541_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n832_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n834_));
OR2X2 OR2X2_443 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3398_), .B(AES_CORE_DATAPATH__abc_16009_new_n3395_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3399_));
OR2X2 OR2X2_4430 ( .A(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_25_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n539_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n835_));
OR2X2 OR2X2_4431 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n837_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n838_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n839_));
OR2X2 OR2X2_4432 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n839_), .B(AES_CORE_DATAPATH_MIX_COL_col_0__2_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n841_));
OR2X2 OR2X2_4433 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n842_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n840_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n843_));
OR2X2 OR2X2_4434 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n844_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n729_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n845_));
OR2X2 OR2X2_4435 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n843_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n727_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n846_));
OR2X2 OR2X2_4436 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n849_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n850_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_26_));
OR2X2 OR2X2_4437 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n852_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n853_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n854_));
OR2X2 OR2X2_4438 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n854_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n857_));
OR2X2 OR2X2_4439 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n860_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n861_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n862_));
OR2X2 OR2X2_444 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3403_), .B(AES_CORE_DATAPATH__abc_16009_new_n3401_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3404_));
OR2X2 OR2X2_4440 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n864_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n865_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_));
OR2X2 OR2X2_4441 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n585_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_27_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n867_));
OR2X2 OR2X2_4442 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n580_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n868_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n869_));
OR2X2 OR2X2_4443 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n871_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n872_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n873_));
OR2X2 OR2X2_4444 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n875_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n876_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n877_));
OR2X2 OR2X2_4445 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n659_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n877_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n880_));
OR2X2 OR2X2_4446 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n883_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n884_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n885_));
OR2X2 OR2X2_4447 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n605_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_28_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n887_));
OR2X2 OR2X2_4448 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n610_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n885_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n888_));
OR2X2 OR2X2_4449 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n890_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n891_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n892_));
OR2X2 OR2X2_445 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3404_), .B(AES_CORE_DATAPATH__abc_16009_new_n2805_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3405_));
OR2X2 OR2X2_4450 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n894_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n895_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n896_));
OR2X2 OR2X2_4451 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n896_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n893_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n897_));
OR2X2 OR2X2_4452 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n898_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n892_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n899_));
OR2X2 OR2X2_4453 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n627_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n900_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n902_));
OR2X2 OR2X2_4454 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n631_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_29_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n903_));
OR2X2 OR2X2_4455 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n905_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n906_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n907_));
OR2X2 OR2X2_4456 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n910_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n908_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n911_));
OR2X2 OR2X2_4457 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n912_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n124_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n913_));
OR2X2 OR2X2_4458 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n911_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n147_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n914_));
OR2X2 OR2X2_4459 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n648_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n916_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n917_));
OR2X2 OR2X2_446 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3407_), .B(AES_CORE_DATAPATH__abc_16009_new_n3408_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3409_));
OR2X2 OR2X2_4460 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n650_), .B(AES_CORE_DATAPATH_MIX_COL_mix_out_enc_30_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n918_));
OR2X2 OR2X2_4461 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n921_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n920_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n922_));
OR2X2 OR2X2_4462 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n923_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n456_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n924_));
OR2X2 OR2X2_4463 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n922_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n453_), .Y(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n925_));
OR2X2 OR2X2_4464 ( .A(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n928_), .B(AES_CORE_DATAPATH_MIX_COL__abc_25207_new_n929_), .Y(AES_CORE_DATAPATH_MIX_COL_mix_out_dec_31_));
OR2X2 OR2X2_4465 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n51_));
OR2X2 OR2X2_4466 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n53_));
OR2X2 OR2X2_4467 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n55_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n56_));
OR2X2 OR2X2_4468 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n58_));
OR2X2 OR2X2_4469 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n64_));
OR2X2 OR2X2_447 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3411_), .B(AES_CORE_DATAPATH__abc_16009_new_n3412_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3413_));
OR2X2 OR2X2_4470 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n69_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n70_));
OR2X2 OR2X2_4471 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n71_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n75_));
OR2X2 OR2X2_4472 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n65_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_));
OR2X2 OR2X2_4473 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n78_));
OR2X2 OR2X2_4474 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n80_));
OR2X2 OR2X2_4475 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n86_));
OR2X2 OR2X2_4476 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n87_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n83_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n88_));
OR2X2 OR2X2_4477 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n91_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n92_));
OR2X2 OR2X2_4478 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n92_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n93_));
OR2X2 OR2X2_4479 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n94_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n96_));
OR2X2 OR2X2_448 ( .A(AES_CORE_DATAPATH_col_sel_host_0_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3417_));
OR2X2 OR2X2_4480 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n97_));
OR2X2 OR2X2_4481 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n103_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n104_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n105_));
OR2X2 OR2X2_4482 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n108_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n109_));
OR2X2 OR2X2_4483 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n111_));
OR2X2 OR2X2_4484 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n112_));
OR2X2 OR2X2_4485 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n110_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_));
OR2X2 OR2X2_4486 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n119_));
OR2X2 OR2X2_4487 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n120_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n121_));
OR2X2 OR2X2_4488 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n124_));
OR2X2 OR2X2_4489 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n125_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n126_));
OR2X2 OR2X2_449 ( .A(AES_CORE_DATAPATH_col_sel_host_1_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3420_));
OR2X2 OR2X2_4490 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n128_));
OR2X2 OR2X2_4491 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n72_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n129_));
OR2X2 OR2X2_4492 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n133_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n134_));
OR2X2 OR2X2_4493 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n134_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n135_));
OR2X2 OR2X2_4494 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n139_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n140_));
OR2X2 OR2X2_4495 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n142_));
OR2X2 OR2X2_4496 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n143_));
OR2X2 OR2X2_4497 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n144_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n145_));
OR2X2 OR2X2_4498 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n146_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n148_));
OR2X2 OR2X2_4499 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n149_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n152_));
OR2X2 OR2X2_45 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n197_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n209_));
OR2X2 OR2X2_450 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3417_), .B(AES_CORE_DATAPATH__abc_16009_new_n3419_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3426_));
OR2X2 OR2X2_4500 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n153_));
OR2X2 OR2X2_4501 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n157_));
OR2X2 OR2X2_4502 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n158_));
OR2X2 OR2X2_4503 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n162_));
OR2X2 OR2X2_4504 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n172_));
OR2X2 OR2X2_4505 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n175_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_));
OR2X2 OR2X2_4506 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n179_));
OR2X2 OR2X2_4507 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n182_));
OR2X2 OR2X2_4508 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n184_));
OR2X2 OR2X2_4509 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n188_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n189_));
OR2X2 OR2X2_451 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3426_), .B(AES_CORE_DATAPATH__abc_16009_new_n3420_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3427_));
OR2X2 OR2X2_4510 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n191_));
OR2X2 OR2X2_4511 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n202_));
OR2X2 OR2X2_4512 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n204_));
OR2X2 OR2X2_4513 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n205_));
OR2X2 OR2X2_4514 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n206_));
OR2X2 OR2X2_4515 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n212_));
OR2X2 OR2X2_4516 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n218_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n219_));
OR2X2 OR2X2_4517 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n220_));
OR2X2 OR2X2_4518 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n222_));
OR2X2 OR2X2_4519 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n224_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n225_));
OR2X2 OR2X2_452 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3425_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3428_));
OR2X2 OR2X2_4520 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n226_));
OR2X2 OR2X2_4521 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n229_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n230_));
OR2X2 OR2X2_4522 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n231_));
OR2X2 OR2X2_4523 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n235_));
OR2X2 OR2X2_4524 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n237_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n238_));
OR2X2 OR2X2_4525 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n240_));
OR2X2 OR2X2_4526 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n240_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n241_));
OR2X2 OR2X2_4527 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n243_));
OR2X2 OR2X2_4528 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n246_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n247_));
OR2X2 OR2X2_4529 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n250_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n251_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n252_));
OR2X2 OR2X2_453 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3420_), .B(AES_CORE_CONTROL_UNIT_sbox_sel_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3434_));
OR2X2 OR2X2_4530 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n252_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n253_));
OR2X2 OR2X2_4531 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n257_));
OR2X2 OR2X2_4532 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n260_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n262_));
OR2X2 OR2X2_4533 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n268_));
OR2X2 OR2X2_4534 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n273_));
OR2X2 OR2X2_4535 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n277_));
OR2X2 OR2X2_4536 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n282_));
OR2X2 OR2X2_4537 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n282_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n283_));
OR2X2 OR2X2_4538 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n287_));
OR2X2 OR2X2_4539 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n292_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n293_));
OR2X2 OR2X2_454 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3434_), .B(AES_CORE_DATAPATH__abc_16009_new_n3417_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3435_));
OR2X2 OR2X2_4540 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n295_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n297_));
OR2X2 OR2X2_4541 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n298_));
OR2X2 OR2X2_4542 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n300_));
OR2X2 OR2X2_4543 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n306_));
OR2X2 OR2X2_4544 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n312_));
OR2X2 OR2X2_4545 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n315_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n317_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n318_));
OR2X2 OR2X2_4546 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n321_));
OR2X2 OR2X2_4547 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n323_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n324_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n325_));
OR2X2 OR2X2_4548 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n325_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n326_));
OR2X2 OR2X2_4549 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n330_));
OR2X2 OR2X2_455 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3433_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3436_));
OR2X2 OR2X2_4550 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n332_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n333_));
OR2X2 OR2X2_4551 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n307_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n334_));
OR2X2 OR2X2_4552 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n340_));
OR2X2 OR2X2_4553 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n342_));
OR2X2 OR2X2_4554 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n344_));
OR2X2 OR2X2_4555 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n351_));
OR2X2 OR2X2_4556 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n352_));
OR2X2 OR2X2_4557 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n357_));
OR2X2 OR2X2_4558 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n359_));
OR2X2 OR2X2_4559 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n361_));
OR2X2 OR2X2_456 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3434_), .B(AES_CORE_DATAPATH__abc_16009_new_n3418_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3437_));
OR2X2 OR2X2_4560 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n362_));
OR2X2 OR2X2_4561 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n365_));
OR2X2 OR2X2_4562 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n367_));
OR2X2 OR2X2_4563 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n369_));
OR2X2 OR2X2_4564 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n370_));
OR2X2 OR2X2_4565 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n371_));
OR2X2 OR2X2_4566 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n373_));
OR2X2 OR2X2_4567 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n374_));
OR2X2 OR2X2_4568 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n376_));
OR2X2 OR2X2_4569 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n379_));
OR2X2 OR2X2_457 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3443_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3444_));
OR2X2 OR2X2_4570 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n380_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n381_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n382_));
OR2X2 OR2X2_4571 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n383_));
OR2X2 OR2X2_4572 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n387_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_2_));
OR2X2 OR2X2_4573 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n392_));
OR2X2 OR2X2_4574 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n395_));
OR2X2 OR2X2_4575 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n396_));
OR2X2 OR2X2_4576 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n398_));
OR2X2 OR2X2_4577 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n399_));
OR2X2 OR2X2_4578 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n400_));
OR2X2 OR2X2_4579 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n402_));
OR2X2 OR2X2_458 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3446_), .B(AES_CORE_DATAPATH__abc_16009_new_n3448_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3449_));
OR2X2 OR2X2_4580 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_7_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n404_));
OR2X2 OR2X2_4581 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n405_));
OR2X2 OR2X2_4582 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n407_));
OR2X2 OR2X2_4583 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n408_));
OR2X2 OR2X2_4584 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n411_));
OR2X2 OR2X2_4585 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n412_));
OR2X2 OR2X2_4586 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n414_));
OR2X2 OR2X2_4587 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n417_));
OR2X2 OR2X2_4588 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n385_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n418_));
OR2X2 OR2X2_4589 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n420_));
OR2X2 OR2X2_459 ( .A(\key_out[0] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3451_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3452_));
OR2X2 OR2X2_4590 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n421_));
OR2X2 OR2X2_4591 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n423_));
OR2X2 OR2X2_4592 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n424_));
OR2X2 OR2X2_4593 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_4_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n425_));
OR2X2 OR2X2_4594 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n427_));
OR2X2 OR2X2_4595 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n429_));
OR2X2 OR2X2_4596 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n430_));
OR2X2 OR2X2_4597 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n432_));
OR2X2 OR2X2_4598 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n433_));
OR2X2 OR2X2_4599 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n294_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n435_));
OR2X2 OR2X2_46 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n209_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n200_), .Y(AES_CORE_CONTROL_UNIT_col_en_3_));
OR2X2 OR2X2_460 ( .A(AES_CORE_CONTROL_UNIT_bypass_rk), .B(AES_CORE_DATAPATH_rk_out_sel_pp2), .Y(AES_CORE_DATAPATH__abc_16009_new_n3455_));
OR2X2 OR2X2_4600 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n436_));
OR2X2 OR2X2_4601 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n440_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_1_));
OR2X2 OR2X2_4602 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n442_));
OR2X2 OR2X2_4603 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n444_));
OR2X2 OR2X2_4604 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n451_));
OR2X2 OR2X2_4605 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n455_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n458_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n459_));
OR2X2 OR2X2_4606 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n462_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n463_));
OR2X2 OR2X2_4607 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n464_));
OR2X2 OR2X2_4608 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n465_));
OR2X2 OR2X2_4609 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n469_));
OR2X2 OR2X2_461 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3454_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3457_));
OR2X2 OR2X2_4610 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n470_));
OR2X2 OR2X2_4611 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n472_));
OR2X2 OR2X2_4612 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n473_));
OR2X2 OR2X2_4613 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n479_));
OR2X2 OR2X2_4614 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n483_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_0_));
OR2X2 OR2X2_4615 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n489_));
OR2X2 OR2X2_4616 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n492_));
OR2X2 OR2X2_4617 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n493_));
OR2X2 OR2X2_4618 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n468_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n496_));
OR2X2 OR2X2_4619 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n497_));
OR2X2 OR2X2_462 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3457_), .B(AES_CORE_DATAPATH__abc_16009_new_n3453_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3458_));
OR2X2 OR2X2_4620 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n500_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n501_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n502_));
OR2X2 OR2X2_4621 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n504_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n502_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n505_));
OR2X2 OR2X2_4622 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n505_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n495_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n506_));
OR2X2 OR2X2_4623 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n508_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n511_));
OR2X2 OR2X2_4624 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n511_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n491_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n512_));
OR2X2 OR2X2_4625 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n515_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n516_));
OR2X2 OR2X2_4626 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n522_));
OR2X2 OR2X2_4627 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n525_));
OR2X2 OR2X2_4628 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n527_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n519_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n528_));
OR2X2 OR2X2_4629 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n526_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n529_));
OR2X2 OR2X2_463 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3461_), .B(AES_CORE_DATAPATH__abc_16009_new_n3459_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3462_));
OR2X2 OR2X2_4630 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n533_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n531_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__out_gf_inv8_stage1_2_));
OR2X2 OR2X2_4631 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n535_));
OR2X2 OR2X2_4632 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n540_));
OR2X2 OR2X2_4633 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n542_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n536_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n543_));
OR2X2 OR2X2_4634 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n541_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n544_));
OR2X2 OR2X2_4635 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n546_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n547_));
OR2X2 OR2X2_4636 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n545_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n507_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n548_));
OR2X2 OR2X2_4637 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n552_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n550_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0__sbox_out_dec_2_));
OR2X2 OR2X2_4638 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n554_));
OR2X2 OR2X2_4639 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_0___abc_26043_new_n555_));
OR2X2 OR2X2_464 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3462_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3463_));
OR2X2 OR2X2_4640 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n51_));
OR2X2 OR2X2_4641 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n53_));
OR2X2 OR2X2_4642 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n55_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n56_));
OR2X2 OR2X2_4643 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n58_));
OR2X2 OR2X2_4644 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n64_));
OR2X2 OR2X2_4645 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n69_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n70_));
OR2X2 OR2X2_4646 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n71_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n75_));
OR2X2 OR2X2_4647 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n65_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_));
OR2X2 OR2X2_4648 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n78_));
OR2X2 OR2X2_4649 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n80_));
OR2X2 OR2X2_465 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3465_), .B(AES_CORE_DATAPATH__abc_16009_new_n3466_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_0_));
OR2X2 OR2X2_4650 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n86_));
OR2X2 OR2X2_4651 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n87_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n83_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n88_));
OR2X2 OR2X2_4652 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n91_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n92_));
OR2X2 OR2X2_4653 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n92_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n93_));
OR2X2 OR2X2_4654 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n94_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n96_));
OR2X2 OR2X2_4655 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n97_));
OR2X2 OR2X2_4656 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n103_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n104_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n105_));
OR2X2 OR2X2_4657 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n108_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n109_));
OR2X2 OR2X2_4658 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n111_));
OR2X2 OR2X2_4659 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n112_));
OR2X2 OR2X2_466 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3468_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3469_));
OR2X2 OR2X2_4660 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n110_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_));
OR2X2 OR2X2_4661 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n119_));
OR2X2 OR2X2_4662 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n120_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n121_));
OR2X2 OR2X2_4663 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n124_));
OR2X2 OR2X2_4664 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n125_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n126_));
OR2X2 OR2X2_4665 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n128_));
OR2X2 OR2X2_4666 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n72_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n129_));
OR2X2 OR2X2_4667 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n133_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n134_));
OR2X2 OR2X2_4668 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n134_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n135_));
OR2X2 OR2X2_4669 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n139_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n140_));
OR2X2 OR2X2_467 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3470_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3471_));
OR2X2 OR2X2_4670 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n142_));
OR2X2 OR2X2_4671 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n143_));
OR2X2 OR2X2_4672 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n144_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n145_));
OR2X2 OR2X2_4673 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n146_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n148_));
OR2X2 OR2X2_4674 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n149_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n152_));
OR2X2 OR2X2_4675 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n153_));
OR2X2 OR2X2_4676 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n157_));
OR2X2 OR2X2_4677 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n158_));
OR2X2 OR2X2_4678 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n162_));
OR2X2 OR2X2_4679 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n172_));
OR2X2 OR2X2_468 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3475_), .B(AES_CORE_DATAPATH__abc_16009_new_n3474_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3476_));
OR2X2 OR2X2_4680 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n175_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_));
OR2X2 OR2X2_4681 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n179_));
OR2X2 OR2X2_4682 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n182_));
OR2X2 OR2X2_4683 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n184_));
OR2X2 OR2X2_4684 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n188_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n189_));
OR2X2 OR2X2_4685 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n191_));
OR2X2 OR2X2_4686 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n202_));
OR2X2 OR2X2_4687 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n204_));
OR2X2 OR2X2_4688 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n205_));
OR2X2 OR2X2_4689 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n206_));
OR2X2 OR2X2_469 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3476_), .B(AES_CORE_DATAPATH__abc_16009_new_n3473_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3477_));
OR2X2 OR2X2_4690 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n212_));
OR2X2 OR2X2_4691 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n218_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n219_));
OR2X2 OR2X2_4692 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n220_));
OR2X2 OR2X2_4693 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n222_));
OR2X2 OR2X2_4694 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n224_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n225_));
OR2X2 OR2X2_4695 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n226_));
OR2X2 OR2X2_4696 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n229_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n230_));
OR2X2 OR2X2_4697 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n231_));
OR2X2 OR2X2_4698 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n235_));
OR2X2 OR2X2_4699 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n237_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n238_));
OR2X2 OR2X2_47 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n213_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n211_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n214_));
OR2X2 OR2X2_470 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3479_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3481_));
OR2X2 OR2X2_4700 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n240_));
OR2X2 OR2X2_4701 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n240_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n241_));
OR2X2 OR2X2_4702 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n243_));
OR2X2 OR2X2_4703 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n246_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n247_));
OR2X2 OR2X2_4704 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n250_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n251_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n252_));
OR2X2 OR2X2_4705 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n252_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n253_));
OR2X2 OR2X2_4706 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n257_));
OR2X2 OR2X2_4707 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n260_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n262_));
OR2X2 OR2X2_4708 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n268_));
OR2X2 OR2X2_4709 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n273_));
OR2X2 OR2X2_471 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3482_), .B(AES_CORE_DATAPATH__abc_16009_new_n3483_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3484_));
OR2X2 OR2X2_4710 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n277_));
OR2X2 OR2X2_4711 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n282_));
OR2X2 OR2X2_4712 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n282_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n283_));
OR2X2 OR2X2_4713 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n287_));
OR2X2 OR2X2_4714 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n292_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n293_));
OR2X2 OR2X2_4715 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n295_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n297_));
OR2X2 OR2X2_4716 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n298_));
OR2X2 OR2X2_4717 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n300_));
OR2X2 OR2X2_4718 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n306_));
OR2X2 OR2X2_4719 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n312_));
OR2X2 OR2X2_472 ( .A(\key_out[1] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3486_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3487_));
OR2X2 OR2X2_4720 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n315_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n317_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n318_));
OR2X2 OR2X2_4721 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n321_));
OR2X2 OR2X2_4722 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n323_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n324_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n325_));
OR2X2 OR2X2_4723 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n325_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n326_));
OR2X2 OR2X2_4724 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n330_));
OR2X2 OR2X2_4725 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n332_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n333_));
OR2X2 OR2X2_4726 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n307_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n334_));
OR2X2 OR2X2_4727 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n340_));
OR2X2 OR2X2_4728 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n342_));
OR2X2 OR2X2_4729 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n344_));
OR2X2 OR2X2_473 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3489_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3490_));
OR2X2 OR2X2_4730 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n351_));
OR2X2 OR2X2_4731 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n352_));
OR2X2 OR2X2_4732 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n357_));
OR2X2 OR2X2_4733 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n359_));
OR2X2 OR2X2_4734 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n361_));
OR2X2 OR2X2_4735 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n362_));
OR2X2 OR2X2_4736 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n365_));
OR2X2 OR2X2_4737 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n367_));
OR2X2 OR2X2_4738 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n369_));
OR2X2 OR2X2_4739 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n370_));
OR2X2 OR2X2_474 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3490_), .B(AES_CORE_DATAPATH__abc_16009_new_n3488_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3491_));
OR2X2 OR2X2_4740 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n371_));
OR2X2 OR2X2_4741 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n373_));
OR2X2 OR2X2_4742 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n374_));
OR2X2 OR2X2_4743 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n376_));
OR2X2 OR2X2_4744 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n379_));
OR2X2 OR2X2_4745 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n380_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n381_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n382_));
OR2X2 OR2X2_4746 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n383_));
OR2X2 OR2X2_4747 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n387_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_10_));
OR2X2 OR2X2_4748 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n392_));
OR2X2 OR2X2_4749 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n395_));
OR2X2 OR2X2_475 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3493_), .B(AES_CORE_DATAPATH__abc_16009_new_n3492_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3494_));
OR2X2 OR2X2_4750 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n396_));
OR2X2 OR2X2_4751 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n398_));
OR2X2 OR2X2_4752 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n399_));
OR2X2 OR2X2_4753 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n400_));
OR2X2 OR2X2_4754 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n402_));
OR2X2 OR2X2_4755 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_15_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n404_));
OR2X2 OR2X2_4756 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n405_));
OR2X2 OR2X2_4757 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n407_));
OR2X2 OR2X2_4758 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_14_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n408_));
OR2X2 OR2X2_4759 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n411_));
OR2X2 OR2X2_476 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3494_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3495_));
OR2X2 OR2X2_4760 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n412_));
OR2X2 OR2X2_4761 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n414_));
OR2X2 OR2X2_4762 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n417_));
OR2X2 OR2X2_4763 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_8_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n385_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n418_));
OR2X2 OR2X2_4764 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n420_));
OR2X2 OR2X2_4765 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n421_));
OR2X2 OR2X2_4766 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n423_));
OR2X2 OR2X2_4767 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n424_));
OR2X2 OR2X2_4768 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_12_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_13_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n425_));
OR2X2 OR2X2_4769 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n427_));
OR2X2 OR2X2_477 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3497_), .B(AES_CORE_DATAPATH__abc_16009_new_n3498_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_1_));
OR2X2 OR2X2_4770 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n429_));
OR2X2 OR2X2_4771 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n430_));
OR2X2 OR2X2_4772 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n432_));
OR2X2 OR2X2_4773 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n433_));
OR2X2 OR2X2_4774 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n294_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n435_));
OR2X2 OR2X2_4775 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n436_));
OR2X2 OR2X2_4776 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n440_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_9_));
OR2X2 OR2X2_4777 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n442_));
OR2X2 OR2X2_4778 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n444_));
OR2X2 OR2X2_4779 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n451_));
OR2X2 OR2X2_478 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3500_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3501_));
OR2X2 OR2X2_4780 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n455_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n458_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n459_));
OR2X2 OR2X2_4781 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n462_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n463_));
OR2X2 OR2X2_4782 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n464_));
OR2X2 OR2X2_4783 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n465_));
OR2X2 OR2X2_4784 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n469_));
OR2X2 OR2X2_4785 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n470_));
OR2X2 OR2X2_4786 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n472_));
OR2X2 OR2X2_4787 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n473_));
OR2X2 OR2X2_4788 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n479_));
OR2X2 OR2X2_4789 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n483_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_0_));
OR2X2 OR2X2_479 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3502_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3503_));
OR2X2 OR2X2_4790 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n489_));
OR2X2 OR2X2_4791 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n492_));
OR2X2 OR2X2_4792 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n493_));
OR2X2 OR2X2_4793 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n468_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n496_));
OR2X2 OR2X2_4794 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n497_));
OR2X2 OR2X2_4795 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n500_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n501_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n502_));
OR2X2 OR2X2_4796 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n504_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n502_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n505_));
OR2X2 OR2X2_4797 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n505_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n495_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n506_));
OR2X2 OR2X2_4798 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n508_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n511_));
OR2X2 OR2X2_4799 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n511_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n491_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n512_));
OR2X2 OR2X2_48 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT_last_round), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n218_));
OR2X2 OR2X2_480 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3507_), .B(AES_CORE_DATAPATH__abc_16009_new_n3506_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3508_));
OR2X2 OR2X2_4800 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n515_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n516_));
OR2X2 OR2X2_4801 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n522_));
OR2X2 OR2X2_4802 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n525_));
OR2X2 OR2X2_4803 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n527_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n519_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n528_));
OR2X2 OR2X2_4804 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n526_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n529_));
OR2X2 OR2X2_4805 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n533_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n531_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__out_gf_inv8_stage1_2_));
OR2X2 OR2X2_4806 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n535_));
OR2X2 OR2X2_4807 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n540_));
OR2X2 OR2X2_4808 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n542_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n536_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n543_));
OR2X2 OR2X2_4809 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n541_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n544_));
OR2X2 OR2X2_481 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3508_), .B(AES_CORE_DATAPATH__abc_16009_new_n3505_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3509_));
OR2X2 OR2X2_4810 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n546_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n547_));
OR2X2 OR2X2_4811 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n545_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n507_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n548_));
OR2X2 OR2X2_4812 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n552_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n550_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1__sbox_out_dec_2_));
OR2X2 OR2X2_4813 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n554_));
OR2X2 OR2X2_4814 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_1___abc_26043_new_n555_));
OR2X2 OR2X2_4815 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n51_));
OR2X2 OR2X2_4816 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n53_));
OR2X2 OR2X2_4817 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n55_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n56_));
OR2X2 OR2X2_4818 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n58_));
OR2X2 OR2X2_4819 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n64_));
OR2X2 OR2X2_482 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3511_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3513_));
OR2X2 OR2X2_4820 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n69_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n70_));
OR2X2 OR2X2_4821 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n71_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n75_));
OR2X2 OR2X2_4822 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n65_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_));
OR2X2 OR2X2_4823 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n78_));
OR2X2 OR2X2_4824 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n80_));
OR2X2 OR2X2_4825 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n86_));
OR2X2 OR2X2_4826 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n87_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n83_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n88_));
OR2X2 OR2X2_4827 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n91_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n92_));
OR2X2 OR2X2_4828 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n92_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n93_));
OR2X2 OR2X2_4829 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n94_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n96_));
OR2X2 OR2X2_483 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3514_), .B(AES_CORE_DATAPATH__abc_16009_new_n3515_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3516_));
OR2X2 OR2X2_4830 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n97_));
OR2X2 OR2X2_4831 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n103_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n104_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n105_));
OR2X2 OR2X2_4832 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n108_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n109_));
OR2X2 OR2X2_4833 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n111_));
OR2X2 OR2X2_4834 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n112_));
OR2X2 OR2X2_4835 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n110_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_));
OR2X2 OR2X2_4836 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n119_));
OR2X2 OR2X2_4837 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n120_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n121_));
OR2X2 OR2X2_4838 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n124_));
OR2X2 OR2X2_4839 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n125_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n126_));
OR2X2 OR2X2_484 ( .A(\key_out[2] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3518_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3519_));
OR2X2 OR2X2_4840 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n128_));
OR2X2 OR2X2_4841 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n72_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n129_));
OR2X2 OR2X2_4842 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n133_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n134_));
OR2X2 OR2X2_4843 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n134_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n135_));
OR2X2 OR2X2_4844 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n139_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n140_));
OR2X2 OR2X2_4845 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n142_));
OR2X2 OR2X2_4846 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n143_));
OR2X2 OR2X2_4847 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n144_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n145_));
OR2X2 OR2X2_4848 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n146_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n148_));
OR2X2 OR2X2_4849 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n149_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n152_));
OR2X2 OR2X2_485 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3521_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3522_));
OR2X2 OR2X2_4850 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n153_));
OR2X2 OR2X2_4851 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n157_));
OR2X2 OR2X2_4852 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n158_));
OR2X2 OR2X2_4853 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n162_));
OR2X2 OR2X2_4854 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n172_));
OR2X2 OR2X2_4855 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n175_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_));
OR2X2 OR2X2_4856 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n179_));
OR2X2 OR2X2_4857 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n182_));
OR2X2 OR2X2_4858 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n184_));
OR2X2 OR2X2_4859 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n188_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n189_));
OR2X2 OR2X2_486 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3522_), .B(AES_CORE_DATAPATH__abc_16009_new_n3520_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3523_));
OR2X2 OR2X2_4860 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n191_));
OR2X2 OR2X2_4861 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n202_));
OR2X2 OR2X2_4862 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n204_));
OR2X2 OR2X2_4863 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n205_));
OR2X2 OR2X2_4864 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n206_));
OR2X2 OR2X2_4865 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n212_));
OR2X2 OR2X2_4866 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n218_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n219_));
OR2X2 OR2X2_4867 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n220_));
OR2X2 OR2X2_4868 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n222_));
OR2X2 OR2X2_4869 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n224_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n225_));
OR2X2 OR2X2_487 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3525_), .B(AES_CORE_DATAPATH__abc_16009_new_n3524_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3526_));
OR2X2 OR2X2_4870 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n226_));
OR2X2 OR2X2_4871 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n229_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n230_));
OR2X2 OR2X2_4872 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n231_));
OR2X2 OR2X2_4873 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n235_));
OR2X2 OR2X2_4874 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n237_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n238_));
OR2X2 OR2X2_4875 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n240_));
OR2X2 OR2X2_4876 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n240_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n241_));
OR2X2 OR2X2_4877 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n243_));
OR2X2 OR2X2_4878 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n246_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n247_));
OR2X2 OR2X2_4879 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n250_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n251_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n252_));
OR2X2 OR2X2_488 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3526_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3527_));
OR2X2 OR2X2_4880 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n252_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n253_));
OR2X2 OR2X2_4881 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n257_));
OR2X2 OR2X2_4882 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n260_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n262_));
OR2X2 OR2X2_4883 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n268_));
OR2X2 OR2X2_4884 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n273_));
OR2X2 OR2X2_4885 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n277_));
OR2X2 OR2X2_4886 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n282_));
OR2X2 OR2X2_4887 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n282_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n283_));
OR2X2 OR2X2_4888 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n287_));
OR2X2 OR2X2_4889 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n292_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n293_));
OR2X2 OR2X2_489 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3529_), .B(AES_CORE_DATAPATH__abc_16009_new_n3530_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_2_));
OR2X2 OR2X2_4890 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n295_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n297_));
OR2X2 OR2X2_4891 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n298_));
OR2X2 OR2X2_4892 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n300_));
OR2X2 OR2X2_4893 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n306_));
OR2X2 OR2X2_4894 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n312_));
OR2X2 OR2X2_4895 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n315_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n317_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n318_));
OR2X2 OR2X2_4896 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n321_));
OR2X2 OR2X2_4897 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n323_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n324_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n325_));
OR2X2 OR2X2_4898 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n325_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n326_));
OR2X2 OR2X2_4899 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n330_));
OR2X2 OR2X2_49 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n219_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n191_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n220_));
OR2X2 OR2X2_490 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3532_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3533_));
OR2X2 OR2X2_4900 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n332_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n333_));
OR2X2 OR2X2_4901 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n307_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n334_));
OR2X2 OR2X2_4902 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n340_));
OR2X2 OR2X2_4903 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n342_));
OR2X2 OR2X2_4904 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n344_));
OR2X2 OR2X2_4905 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n351_));
OR2X2 OR2X2_4906 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n352_));
OR2X2 OR2X2_4907 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n357_));
OR2X2 OR2X2_4908 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n359_));
OR2X2 OR2X2_4909 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n361_));
OR2X2 OR2X2_491 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3534_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3535_));
OR2X2 OR2X2_4910 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n362_));
OR2X2 OR2X2_4911 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n365_));
OR2X2 OR2X2_4912 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n367_));
OR2X2 OR2X2_4913 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n369_));
OR2X2 OR2X2_4914 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n370_));
OR2X2 OR2X2_4915 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n371_));
OR2X2 OR2X2_4916 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n373_));
OR2X2 OR2X2_4917 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n374_));
OR2X2 OR2X2_4918 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n376_));
OR2X2 OR2X2_4919 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n379_));
OR2X2 OR2X2_492 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3539_), .B(AES_CORE_DATAPATH__abc_16009_new_n3538_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3540_));
OR2X2 OR2X2_4920 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n380_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n381_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n382_));
OR2X2 OR2X2_4921 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n383_));
OR2X2 OR2X2_4922 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n387_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_18_));
OR2X2 OR2X2_4923 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n392_));
OR2X2 OR2X2_4924 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n395_));
OR2X2 OR2X2_4925 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n396_));
OR2X2 OR2X2_4926 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n398_));
OR2X2 OR2X2_4927 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n399_));
OR2X2 OR2X2_4928 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n400_));
OR2X2 OR2X2_4929 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n402_));
OR2X2 OR2X2_493 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3540_), .B(AES_CORE_DATAPATH__abc_16009_new_n3537_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3541_));
OR2X2 OR2X2_4930 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_23_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n404_));
OR2X2 OR2X2_4931 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n405_));
OR2X2 OR2X2_4932 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n407_));
OR2X2 OR2X2_4933 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_22_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n408_));
OR2X2 OR2X2_4934 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n411_));
OR2X2 OR2X2_4935 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n412_));
OR2X2 OR2X2_4936 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n414_));
OR2X2 OR2X2_4937 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n417_));
OR2X2 OR2X2_4938 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_16_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n385_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n418_));
OR2X2 OR2X2_4939 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n420_));
OR2X2 OR2X2_494 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3543_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3545_));
OR2X2 OR2X2_4940 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n421_));
OR2X2 OR2X2_4941 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n423_));
OR2X2 OR2X2_4942 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n424_));
OR2X2 OR2X2_4943 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_20_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_21_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n425_));
OR2X2 OR2X2_4944 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n427_));
OR2X2 OR2X2_4945 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n429_));
OR2X2 OR2X2_4946 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n430_));
OR2X2 OR2X2_4947 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n432_));
OR2X2 OR2X2_4948 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n433_));
OR2X2 OR2X2_4949 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n294_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n435_));
OR2X2 OR2X2_495 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3546_), .B(AES_CORE_DATAPATH__abc_16009_new_n3547_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3548_));
OR2X2 OR2X2_4950 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n436_));
OR2X2 OR2X2_4951 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n440_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_func_17_));
OR2X2 OR2X2_4952 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n442_));
OR2X2 OR2X2_4953 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n444_));
OR2X2 OR2X2_4954 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n451_));
OR2X2 OR2X2_4955 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n455_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n458_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n459_));
OR2X2 OR2X2_4956 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n462_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n463_));
OR2X2 OR2X2_4957 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n464_));
OR2X2 OR2X2_4958 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n465_));
OR2X2 OR2X2_4959 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n469_));
OR2X2 OR2X2_496 ( .A(\key_out[3] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3550_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3551_));
OR2X2 OR2X2_4960 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n470_));
OR2X2 OR2X2_4961 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n472_));
OR2X2 OR2X2_4962 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n473_));
OR2X2 OR2X2_4963 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n479_));
OR2X2 OR2X2_4964 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n483_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_0_));
OR2X2 OR2X2_4965 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n489_));
OR2X2 OR2X2_4966 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n492_));
OR2X2 OR2X2_4967 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n493_));
OR2X2 OR2X2_4968 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n468_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n496_));
OR2X2 OR2X2_4969 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n497_));
OR2X2 OR2X2_497 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3553_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3554_));
OR2X2 OR2X2_4970 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n500_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n501_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n502_));
OR2X2 OR2X2_4971 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n504_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n502_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n505_));
OR2X2 OR2X2_4972 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n505_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n495_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n506_));
OR2X2 OR2X2_4973 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n508_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n511_));
OR2X2 OR2X2_4974 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n511_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n491_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n512_));
OR2X2 OR2X2_4975 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n515_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n516_));
OR2X2 OR2X2_4976 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n522_));
OR2X2 OR2X2_4977 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n525_));
OR2X2 OR2X2_4978 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n527_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n519_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n528_));
OR2X2 OR2X2_4979 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n526_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n529_));
OR2X2 OR2X2_498 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3554_), .B(AES_CORE_DATAPATH__abc_16009_new_n3552_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3555_));
OR2X2 OR2X2_4980 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n533_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n531_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__out_gf_inv8_stage1_2_));
OR2X2 OR2X2_4981 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n535_));
OR2X2 OR2X2_4982 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n540_));
OR2X2 OR2X2_4983 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n542_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n536_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n543_));
OR2X2 OR2X2_4984 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n541_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n544_));
OR2X2 OR2X2_4985 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n546_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n547_));
OR2X2 OR2X2_4986 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n545_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n507_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n548_));
OR2X2 OR2X2_4987 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n552_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n550_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2__sbox_out_dec_2_));
OR2X2 OR2X2_4988 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n554_));
OR2X2 OR2X2_4989 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_2___abc_26043_new_n555_));
OR2X2 OR2X2_499 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3557_), .B(AES_CORE_DATAPATH__abc_16009_new_n3556_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3558_));
OR2X2 OR2X2_4990 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n51_));
OR2X2 OR2X2_4991 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n53_));
OR2X2 OR2X2_4992 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n55_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n56_));
OR2X2 OR2X2_4993 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n58_));
OR2X2 OR2X2_4994 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n61_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n63_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n64_));
OR2X2 OR2X2_4995 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n68_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n69_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n70_));
OR2X2 OR2X2_4996 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n74_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n71_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n75_));
OR2X2 OR2X2_4997 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n76_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n65_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_));
OR2X2 OR2X2_4998 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n50_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n78_));
OR2X2 OR2X2_4999 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n80_));
OR2X2 OR2X2_5 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n109_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n101_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_2_));
OR2X2 OR2X2_50 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n220_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n217_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n221_));
OR2X2 OR2X2_500 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3558_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3559_));
OR2X2 OR2X2_5000 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n85_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n84_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n86_));
OR2X2 OR2X2_5001 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n87_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n83_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n88_));
OR2X2 OR2X2_5002 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n90_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n91_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n92_));
OR2X2 OR2X2_5003 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n92_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n93_));
OR2X2 OR2X2_5004 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n94_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n95_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n96_));
OR2X2 OR2X2_5005 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n96_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n97_));
OR2X2 OR2X2_5006 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n103_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n104_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n105_));
OR2X2 OR2X2_5007 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n106_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n108_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n109_));
OR2X2 OR2X2_5008 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n57_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n111_));
OR2X2 OR2X2_5009 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n112_));
OR2X2 OR2X2_501 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3561_), .B(AES_CORE_DATAPATH__abc_16009_new_n3562_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_3_));
OR2X2 OR2X2_5010 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n110_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n115_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_));
OR2X2 OR2X2_5011 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n75_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n102_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n119_));
OR2X2 OR2X2_5012 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n120_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n121_));
OR2X2 OR2X2_5013 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n86_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n79_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n124_));
OR2X2 OR2X2_5014 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n125_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n126_));
OR2X2 OR2X2_5015 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n52_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_3_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n128_));
OR2X2 OR2X2_5016 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n72_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n129_));
OR2X2 OR2X2_5017 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n133_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n134_));
OR2X2 OR2X2_5018 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n134_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n132_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n135_));
OR2X2 OR2X2_5019 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n138_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n139_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n140_));
OR2X2 OR2X2_502 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3565_));
OR2X2 OR2X2_5020 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n81_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n57_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n142_));
OR2X2 OR2X2_5021 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n82_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_in_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n143_));
OR2X2 OR2X2_5022 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n144_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_enc_dec), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n145_));
OR2X2 OR2X2_5023 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n146_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n147_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n148_));
OR2X2 OR2X2_5024 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n151_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n149_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n152_));
OR2X2 OR2X2_5025 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n152_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n66_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n153_));
OR2X2 OR2X2_5026 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_0_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n157_));
OR2X2 OR2X2_5027 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n157_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n156_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n158_));
OR2X2 OR2X2_5028 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n161_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n159_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n162_));
OR2X2 OR2X2_5029 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_pp_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n172_));
OR2X2 OR2X2_503 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3566_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3567_));
OR2X2 OR2X2_5030 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n175_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n167_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_));
OR2X2 OR2X2_5031 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n166_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n179_));
OR2X2 OR2X2_5032 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n181_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n182_));
OR2X2 OR2X2_5033 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n183_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_5_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n184_));
OR2X2 OR2X2_5034 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n188_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_6_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n189_));
OR2X2 OR2X2_5035 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n190_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_pp_4_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n191_));
OR2X2 OR2X2_5036 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n201_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n202_));
OR2X2 OR2X2_5037 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n195_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n203_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n204_));
OR2X2 OR2X2_5038 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n193_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n197_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n205_));
OR2X2 OR2X2_5039 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n205_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n202_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n206_));
OR2X2 OR2X2_504 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3571_), .B(AES_CORE_DATAPATH__abc_16009_new_n3570_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3572_));
OR2X2 OR2X2_5040 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n211_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n210_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n212_));
OR2X2 OR2X2_5041 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n218_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n177_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n219_));
OR2X2 OR2X2_5042 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n185_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n220_));
OR2X2 OR2X2_5043 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n221_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n222_));
OR2X2 OR2X2_5044 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n224_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n209_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n225_));
OR2X2 OR2X2_5045 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n176_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n205_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n226_));
OR2X2 OR2X2_5046 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n228_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n229_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n230_));
OR2X2 OR2X2_5047 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n230_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n231_));
OR2X2 OR2X2_5048 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n231_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n232_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n235_));
OR2X2 OR2X2_5049 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n237_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n238_));
OR2X2 OR2X2_505 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3572_), .B(AES_CORE_DATAPATH__abc_16009_new_n3569_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3573_));
OR2X2 OR2X2_5050 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n187_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n208_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n240_));
OR2X2 OR2X2_5051 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n240_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n213_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n241_));
OR2X2 OR2X2_5052 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n236_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n243_));
OR2X2 OR2X2_5053 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n246_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n196_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n247_));
OR2X2 OR2X2_5054 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n250_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n251_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n252_));
OR2X2 OR2X2_5055 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n252_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n253_));
OR2X2 OR2X2_5056 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n254_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n257_));
OR2X2 OR2X2_5057 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n260_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n261_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n262_));
OR2X2 OR2X2_5058 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n266_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n267_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n268_));
OR2X2 OR2X2_5059 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n264_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n270_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n273_));
OR2X2 OR2X2_506 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3575_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3577_));
OR2X2 OR2X2_5060 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n274_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n258_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n277_));
OR2X2 OR2X2_5061 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n280_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n281_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n282_));
OR2X2 OR2X2_5062 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n227_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n282_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n283_));
OR2X2 OR2X2_5063 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n284_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n287_));
OR2X2 OR2X2_5064 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n291_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n292_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n293_));
OR2X2 OR2X2_5065 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n295_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n296_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n297_));
OR2X2 OR2X2_5066 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n297_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n298_));
OR2X2 OR2X2_5067 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n299_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n300_));
OR2X2 OR2X2_5068 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n302_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n303_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n306_));
OR2X2 OR2X2_5069 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n308_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n309_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n312_));
OR2X2 OR2X2_507 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3578_), .B(AES_CORE_DATAPATH__abc_16009_new_n3579_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3580_));
OR2X2 OR2X2_5070 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n315_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n317_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n318_));
OR2X2 OR2X2_5071 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n318_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n321_));
OR2X2 OR2X2_5072 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n323_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n324_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n325_));
OR2X2 OR2X2_5073 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n247_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n325_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n326_));
OR2X2 OR2X2_5074 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n327_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n330_));
OR2X2 OR2X2_5075 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n316_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n332_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n333_));
OR2X2 OR2X2_5076 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n307_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n331_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n334_));
OR2X2 OR2X2_5077 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n326_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n337_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n340_));
OR2X2 OR2X2_5078 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n342_));
OR2X2 OR2X2_5079 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n344_));
OR2X2 OR2X2_508 ( .A(\key_out[4] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3582_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3583_));
OR2X2 OR2X2_5080 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n346_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n347_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n351_));
OR2X2 OR2X2_5081 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n351_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n350_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n352_));
OR2X2 OR2X2_5082 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n283_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n354_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n357_));
OR2X2 OR2X2_5083 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n359_));
OR2X2 OR2X2_5084 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n219_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n262_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n361_));
OR2X2 OR2X2_5085 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n212_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n269_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n362_));
OR2X2 OR2X2_5086 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n364_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n348_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n365_));
OR2X2 OR2X2_5087 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n367_));
OR2X2 OR2X2_5088 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n369_));
OR2X2 OR2X2_5089 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n242_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n343_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n370_));
OR2X2 OR2X2_509 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3585_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3586_));
OR2X2 OR2X2_5090 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n225_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n341_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n371_));
OR2X2 OR2X2_5091 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n358_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n373_));
OR2X2 OR2X2_5092 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n366_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n374_));
OR2X2 OR2X2_5093 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n376_));
OR2X2 OR2X2_5094 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n379_));
OR2X2 OR2X2_5095 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n380_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n381_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n382_));
OR2X2 OR2X2_5096 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n383_));
OR2X2 OR2X2_5097 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n386_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n387_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_26_));
OR2X2 OR2X2_5098 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n253_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n389_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n392_));
OR2X2 OR2X2_5099 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n395_));
OR2X2 OR2X2_51 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n223_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n138_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n224_));
OR2X2 OR2X2_510 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3586_), .B(AES_CORE_DATAPATH__abc_16009_new_n3584_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3587_));
OR2X2 OR2X2_5100 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n396_));
OR2X2 OR2X2_5101 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n372_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n398_));
OR2X2 OR2X2_5102 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n365_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n393_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n399_));
OR2X2 OR2X2_5103 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n353_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n394_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n400_));
OR2X2 OR2X2_5104 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n345_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n402_));
OR2X2 OR2X2_5105 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_31_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n401_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n404_));
OR2X2 OR2X2_5106 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n382_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n397_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n405_));
OR2X2 OR2X2_5107 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n299_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n407_));
OR2X2 OR2X2_5108 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_30_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n408_));
OR2X2 OR2X2_5109 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n409_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n410_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n411_));
OR2X2 OR2X2_511 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3589_), .B(AES_CORE_DATAPATH__abc_16009_new_n3588_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3590_));
OR2X2 OR2X2_5110 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n411_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n412_));
OR2X2 OR2X2_5111 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n297_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n414_));
OR2X2 OR2X2_5112 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n416_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n384_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n417_));
OR2X2 OR2X2_5113 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_24_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n385_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n418_));
OR2X2 OR2X2_5114 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n420_));
OR2X2 OR2X2_5115 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n421_));
OR2X2 OR2X2_5116 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_1_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n423_));
OR2X2 OR2X2_5117 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n406_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n378_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n424_));
OR2X2 OR2X2_5118 ( .A(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_28_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_29_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n425_));
OR2X2 OR2X2_5119 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n335_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n427_));
OR2X2 OR2X2_512 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3590_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3591_));
OR2X2 OR2X2_5120 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n422_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n429_));
OR2X2 OR2X2_5121 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n426_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n430_));
OR2X2 OR2X2_5122 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n368_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n432_));
OR2X2 OR2X2_5123 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n375_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n433_));
OR2X2 OR2X2_5124 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n294_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n435_));
OR2X2 OR2X2_5125 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n293_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n436_));
OR2X2 OR2X2_5126 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n439_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n440_), .Y(AES_CORE_DATAPATH_KEY_EXPANDER_g_out_25_));
OR2X2 OR2X2_5127 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n442_));
OR2X2 OR2X2_5128 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n444_));
OR2X2 OR2X2_5129 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_4_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n451_));
OR2X2 OR2X2_513 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3593_), .B(AES_CORE_DATAPATH__abc_16009_new_n3594_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_4_));
OR2X2 OR2X2_5130 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n455_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n458_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n459_));
OR2X2 OR2X2_5131 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n462_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n461_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n463_));
OR2X2 OR2X2_5132 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_0_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n464_));
OR2X2 OR2X2_5133 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n443_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n465_));
OR2X2 OR2X2_5134 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n468_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n88_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n469_));
OR2X2 OR2X2_5135 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_5_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n470_));
OR2X2 OR2X2_5136 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_1_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n472_));
OR2X2 OR2X2_5137 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n136_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n473_));
OR2X2 OR2X2_5138 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n467_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n476_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n479_));
OR2X2 OR2X2_5139 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n482_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n483_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_0_));
OR2X2 OR2X2_514 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3596_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3597_));
OR2X2 OR2X2_5140 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n486_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n457_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n489_));
OR2X2 OR2X2_5141 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n154_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_2_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n492_));
OR2X2 OR2X2_5142 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_3_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n140_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n493_));
OR2X2 OR2X2_5143 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_6_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n468_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n496_));
OR2X2 OR2X2_5144 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n100_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3__base_new_7_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n497_));
OR2X2 OR2X2_5145 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n500_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n501_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n502_));
OR2X2 OR2X2_5146 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n504_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n502_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n505_));
OR2X2 OR2X2_5147 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n505_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n495_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n506_));
OR2X2 OR2X2_5148 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n508_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n510_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n511_));
OR2X2 OR2X2_5149 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n511_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n491_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n512_));
OR2X2 OR2X2_515 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3598_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3599_));
OR2X2 OR2X2_5150 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n515_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n490_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n516_));
OR2X2 OR2X2_5151 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n475_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n471_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n522_));
OR2X2 OR2X2_5152 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n522_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n521_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n525_));
OR2X2 OR2X2_5153 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n527_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n519_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n528_));
OR2X2 OR2X2_5154 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n526_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n518_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n529_));
OR2X2 OR2X2_5155 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n533_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n531_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__out_gf_inv8_stage1_2_));
OR2X2 OR2X2_5156 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n466_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n463_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n535_));
OR2X2 OR2X2_5157 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n518_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n537_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n540_));
OR2X2 OR2X2_5158 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n542_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n536_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n543_));
OR2X2 OR2X2_5159 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n541_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n535_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n544_));
OR2X2 OR2X2_516 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3603_), .B(AES_CORE_DATAPATH__abc_16009_new_n3602_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3604_));
OR2X2 OR2X2_5160 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n546_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n506_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n547_));
OR2X2 OR2X2_5161 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n545_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n507_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n548_));
OR2X2 OR2X2_5162 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n552_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n550_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3__sbox_out_dec_2_));
OR2X2 OR2X2_5163 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n245_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n278_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n554_));
OR2X2 OR2X2_5164 ( .A(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n279_), .B(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n244_), .Y(AES_CORE_DATAPATH_SBOX_SBOX_3___abc_26043_new_n555_));
OR2X2 OR2X2_5165 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n69_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n73_));
OR2X2 OR2X2_5166 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n75_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n77_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n78_));
OR2X2 OR2X2_5167 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n73_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n78_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_0_));
OR2X2 OR2X2_5168 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n80_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n81_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n82_));
OR2X2 OR2X2_5169 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n83_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n84_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n85_));
OR2X2 OR2X2_517 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3604_), .B(AES_CORE_DATAPATH__abc_16009_new_n3601_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3605_));
OR2X2 OR2X2_5170 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n82_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n85_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_1_));
OR2X2 OR2X2_5171 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n87_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n88_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n89_));
OR2X2 OR2X2_5172 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n90_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n91_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n92_));
OR2X2 OR2X2_5173 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n89_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n92_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_2_));
OR2X2 OR2X2_5174 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n94_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n95_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n96_));
OR2X2 OR2X2_5175 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n97_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n98_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n99_));
OR2X2 OR2X2_5176 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n96_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n99_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_3_));
OR2X2 OR2X2_5177 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n101_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n102_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n103_));
OR2X2 OR2X2_5178 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n104_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n105_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n106_));
OR2X2 OR2X2_5179 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n103_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n106_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_4_));
OR2X2 OR2X2_518 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3607_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3609_));
OR2X2 OR2X2_5180 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n108_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n109_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n110_));
OR2X2 OR2X2_5181 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n111_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n112_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n113_));
OR2X2 OR2X2_5182 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n110_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n113_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_5_));
OR2X2 OR2X2_5183 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n115_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n116_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n117_));
OR2X2 OR2X2_5184 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n118_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n119_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n120_));
OR2X2 OR2X2_5185 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n117_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n120_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_6_));
OR2X2 OR2X2_5186 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n122_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n123_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n124_));
OR2X2 OR2X2_5187 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n125_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n126_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n127_));
OR2X2 OR2X2_5188 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n124_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n127_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_7_));
OR2X2 OR2X2_5189 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n129_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n130_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n131_));
OR2X2 OR2X2_519 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3610_), .B(AES_CORE_DATAPATH__abc_16009_new_n3611_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3612_));
OR2X2 OR2X2_5190 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n132_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n133_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n134_));
OR2X2 OR2X2_5191 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n131_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n134_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_8_));
OR2X2 OR2X2_5192 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n136_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n137_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n138_));
OR2X2 OR2X2_5193 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n139_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n140_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n141_));
OR2X2 OR2X2_5194 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n138_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n141_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_9_));
OR2X2 OR2X2_5195 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n143_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n144_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n145_));
OR2X2 OR2X2_5196 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n146_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n147_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n148_));
OR2X2 OR2X2_5197 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n145_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n148_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_10_));
OR2X2 OR2X2_5198 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n150_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n151_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n152_));
OR2X2 OR2X2_5199 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n153_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n154_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n155_));
OR2X2 OR2X2_52 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n224_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n152_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n225_));
OR2X2 OR2X2_520 ( .A(\key_out[5] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3614_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3615_));
OR2X2 OR2X2_5200 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n152_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n155_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_11_));
OR2X2 OR2X2_5201 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n157_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n158_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n159_));
OR2X2 OR2X2_5202 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n160_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n161_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n162_));
OR2X2 OR2X2_5203 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n159_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n162_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_12_));
OR2X2 OR2X2_5204 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n164_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n165_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n166_));
OR2X2 OR2X2_5205 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n167_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n168_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n169_));
OR2X2 OR2X2_5206 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n166_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n169_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_13_));
OR2X2 OR2X2_5207 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n171_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n172_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n173_));
OR2X2 OR2X2_5208 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n174_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n175_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n176_));
OR2X2 OR2X2_5209 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n173_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n176_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_14_));
OR2X2 OR2X2_521 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3617_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3618_));
OR2X2 OR2X2_5210 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n178_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n179_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n180_));
OR2X2 OR2X2_5211 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n181_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n182_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n183_));
OR2X2 OR2X2_5212 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n180_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n183_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_15_));
OR2X2 OR2X2_5213 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n185_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n186_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n187_));
OR2X2 OR2X2_5214 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n188_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n189_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n190_));
OR2X2 OR2X2_5215 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n187_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n190_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_16_));
OR2X2 OR2X2_5216 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n192_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n193_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n194_));
OR2X2 OR2X2_5217 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n195_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n196_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n197_));
OR2X2 OR2X2_5218 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n194_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n197_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_17_));
OR2X2 OR2X2_5219 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n199_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n200_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n201_));
OR2X2 OR2X2_522 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3618_), .B(AES_CORE_DATAPATH__abc_16009_new_n3616_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3619_));
OR2X2 OR2X2_5220 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n202_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n203_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n204_));
OR2X2 OR2X2_5221 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n201_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n204_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_18_));
OR2X2 OR2X2_5222 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n206_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n207_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n208_));
OR2X2 OR2X2_5223 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n209_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n210_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n211_));
OR2X2 OR2X2_5224 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n208_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n211_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_19_));
OR2X2 OR2X2_5225 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n213_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n214_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n215_));
OR2X2 OR2X2_5226 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n216_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n217_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n218_));
OR2X2 OR2X2_5227 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n215_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n218_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_20_));
OR2X2 OR2X2_5228 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n220_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n221_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n222_));
OR2X2 OR2X2_5229 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n223_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n224_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n225_));
OR2X2 OR2X2_523 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3621_), .B(AES_CORE_DATAPATH__abc_16009_new_n3620_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3622_));
OR2X2 OR2X2_5230 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n222_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n225_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_21_));
OR2X2 OR2X2_5231 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n227_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n228_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n229_));
OR2X2 OR2X2_5232 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n230_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n231_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n232_));
OR2X2 OR2X2_5233 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n229_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n232_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_22_));
OR2X2 OR2X2_5234 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n234_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n235_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n236_));
OR2X2 OR2X2_5235 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n237_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n238_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n239_));
OR2X2 OR2X2_5236 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n236_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n239_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_23_));
OR2X2 OR2X2_5237 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n241_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n242_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n243_));
OR2X2 OR2X2_5238 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n244_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n245_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n246_));
OR2X2 OR2X2_5239 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n243_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n246_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_24_));
OR2X2 OR2X2_524 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3622_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3623_));
OR2X2 OR2X2_5240 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n248_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n249_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n250_));
OR2X2 OR2X2_5241 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n251_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n252_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n253_));
OR2X2 OR2X2_5242 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n250_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n253_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_25_));
OR2X2 OR2X2_5243 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n255_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n256_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n257_));
OR2X2 OR2X2_5244 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n258_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n259_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n260_));
OR2X2 OR2X2_5245 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n257_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n260_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_26_));
OR2X2 OR2X2_5246 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n262_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n263_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n264_));
OR2X2 OR2X2_5247 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n265_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n266_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n267_));
OR2X2 OR2X2_5248 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n264_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n267_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_27_));
OR2X2 OR2X2_5249 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n269_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n270_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n271_));
OR2X2 OR2X2_525 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3625_), .B(AES_CORE_DATAPATH__abc_16009_new_n3626_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_5_));
OR2X2 OR2X2_5250 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n272_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n273_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n274_));
OR2X2 OR2X2_5251 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n271_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n274_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_28_));
OR2X2 OR2X2_5252 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n276_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n277_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n278_));
OR2X2 OR2X2_5253 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n279_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n280_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n281_));
OR2X2 OR2X2_5254 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n278_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n281_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_29_));
OR2X2 OR2X2_5255 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n283_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n284_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n285_));
OR2X2 OR2X2_5256 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n286_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n287_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n288_));
OR2X2 OR2X2_5257 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n285_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n288_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_30_));
OR2X2 OR2X2_5258 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n290_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n291_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n292_));
OR2X2 OR2X2_5259 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n293_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n294_), .Y(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n295_));
OR2X2 OR2X2_526 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3628_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3629_));
OR2X2 OR2X2_5260 ( .A(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n292_), .B(AES_CORE_DATAPATH_SWAP_IN__abc_15778_new_n295_), .Y(AES_CORE_DATAPATH_SWAP_IN_data_swap_31_));
OR2X2 OR2X2_5261 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n69_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n72_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n73_));
OR2X2 OR2X2_5262 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n75_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n77_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n78_));
OR2X2 OR2X2_5263 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n73_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n78_), .Y(\col_out[0] ));
OR2X2 OR2X2_5264 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n80_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n81_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n82_));
OR2X2 OR2X2_5265 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n83_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n84_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n85_));
OR2X2 OR2X2_5266 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n82_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n85_), .Y(\col_out[1] ));
OR2X2 OR2X2_5267 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n87_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n88_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n89_));
OR2X2 OR2X2_5268 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n90_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n91_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n92_));
OR2X2 OR2X2_5269 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n89_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n92_), .Y(\col_out[2] ));
OR2X2 OR2X2_527 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3630_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3631_));
OR2X2 OR2X2_5270 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n94_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n95_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n96_));
OR2X2 OR2X2_5271 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n97_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n98_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n99_));
OR2X2 OR2X2_5272 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n96_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n99_), .Y(\col_out[3] ));
OR2X2 OR2X2_5273 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n101_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n102_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n103_));
OR2X2 OR2X2_5274 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n104_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n105_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n106_));
OR2X2 OR2X2_5275 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n103_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n106_), .Y(\col_out[4] ));
OR2X2 OR2X2_5276 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n108_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n109_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n110_));
OR2X2 OR2X2_5277 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n111_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n112_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n113_));
OR2X2 OR2X2_5278 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n110_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n113_), .Y(\col_out[5] ));
OR2X2 OR2X2_5279 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n115_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n116_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n117_));
OR2X2 OR2X2_528 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3635_), .B(AES_CORE_DATAPATH__abc_16009_new_n3634_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3636_));
OR2X2 OR2X2_5280 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n118_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n119_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n120_));
OR2X2 OR2X2_5281 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n117_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n120_), .Y(\col_out[6] ));
OR2X2 OR2X2_5282 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n122_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n123_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n124_));
OR2X2 OR2X2_5283 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n125_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n126_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n127_));
OR2X2 OR2X2_5284 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n124_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n127_), .Y(\col_out[7] ));
OR2X2 OR2X2_5285 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n129_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n130_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n131_));
OR2X2 OR2X2_5286 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n132_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n133_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n134_));
OR2X2 OR2X2_5287 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n131_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n134_), .Y(\col_out[8] ));
OR2X2 OR2X2_5288 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n136_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n137_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n138_));
OR2X2 OR2X2_5289 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n139_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n140_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n141_));
OR2X2 OR2X2_529 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3636_), .B(AES_CORE_DATAPATH__abc_16009_new_n3633_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3637_));
OR2X2 OR2X2_5290 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n138_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n141_), .Y(\col_out[9] ));
OR2X2 OR2X2_5291 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n143_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n144_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n145_));
OR2X2 OR2X2_5292 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n146_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n147_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n148_));
OR2X2 OR2X2_5293 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n145_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n148_), .Y(\col_out[10] ));
OR2X2 OR2X2_5294 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n150_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n151_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n152_));
OR2X2 OR2X2_5295 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n153_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n154_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n155_));
OR2X2 OR2X2_5296 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n152_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n155_), .Y(\col_out[11] ));
OR2X2 OR2X2_5297 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n157_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n158_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n159_));
OR2X2 OR2X2_5298 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n160_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n161_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n162_));
OR2X2 OR2X2_5299 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n159_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n162_), .Y(\col_out[12] ));
OR2X2 OR2X2_53 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n222_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n225_), .Y(AES_CORE_CONTROL_UNIT_col_sel_0_));
OR2X2 OR2X2_530 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3639_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3641_));
OR2X2 OR2X2_5300 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n164_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n165_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n166_));
OR2X2 OR2X2_5301 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n167_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n168_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n169_));
OR2X2 OR2X2_5302 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n166_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n169_), .Y(\col_out[13] ));
OR2X2 OR2X2_5303 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n171_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n172_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n173_));
OR2X2 OR2X2_5304 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n174_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n175_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n176_));
OR2X2 OR2X2_5305 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n173_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n176_), .Y(\col_out[14] ));
OR2X2 OR2X2_5306 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n178_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n179_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n180_));
OR2X2 OR2X2_5307 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n181_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n182_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n183_));
OR2X2 OR2X2_5308 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n180_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n183_), .Y(\col_out[15] ));
OR2X2 OR2X2_5309 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n185_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n186_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n187_));
OR2X2 OR2X2_531 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3642_), .B(AES_CORE_DATAPATH__abc_16009_new_n3643_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3644_));
OR2X2 OR2X2_5310 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n188_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n189_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n190_));
OR2X2 OR2X2_5311 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n187_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n190_), .Y(\col_out[16] ));
OR2X2 OR2X2_5312 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n192_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n193_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n194_));
OR2X2 OR2X2_5313 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n195_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n196_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n197_));
OR2X2 OR2X2_5314 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n194_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n197_), .Y(\col_out[17] ));
OR2X2 OR2X2_5315 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n199_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n200_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n201_));
OR2X2 OR2X2_5316 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n202_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n203_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n204_));
OR2X2 OR2X2_5317 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n201_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n204_), .Y(\col_out[18] ));
OR2X2 OR2X2_5318 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n206_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n207_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n208_));
OR2X2 OR2X2_5319 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n209_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n210_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n211_));
OR2X2 OR2X2_532 ( .A(\key_out[6] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3646_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3647_));
OR2X2 OR2X2_5320 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n208_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n211_), .Y(\col_out[19] ));
OR2X2 OR2X2_5321 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n213_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n214_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n215_));
OR2X2 OR2X2_5322 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n216_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n217_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n218_));
OR2X2 OR2X2_5323 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n215_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n218_), .Y(\col_out[20] ));
OR2X2 OR2X2_5324 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n220_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n221_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n222_));
OR2X2 OR2X2_5325 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n223_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n224_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n225_));
OR2X2 OR2X2_5326 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n222_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n225_), .Y(\col_out[21] ));
OR2X2 OR2X2_5327 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n227_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n228_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n229_));
OR2X2 OR2X2_5328 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n230_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n231_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n232_));
OR2X2 OR2X2_5329 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n229_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n232_), .Y(\col_out[22] ));
OR2X2 OR2X2_533 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3649_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3650_));
OR2X2 OR2X2_5330 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n234_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n235_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n236_));
OR2X2 OR2X2_5331 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n237_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n238_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n239_));
OR2X2 OR2X2_5332 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n236_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n239_), .Y(\col_out[23] ));
OR2X2 OR2X2_5333 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n241_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n242_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n243_));
OR2X2 OR2X2_5334 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n244_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n245_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n246_));
OR2X2 OR2X2_5335 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n243_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n246_), .Y(\col_out[24] ));
OR2X2 OR2X2_5336 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n248_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n249_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n250_));
OR2X2 OR2X2_5337 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n251_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n252_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n253_));
OR2X2 OR2X2_5338 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n250_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n253_), .Y(\col_out[25] ));
OR2X2 OR2X2_5339 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n255_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n256_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n257_));
OR2X2 OR2X2_534 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3650_), .B(AES_CORE_DATAPATH__abc_16009_new_n3648_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3651_));
OR2X2 OR2X2_5340 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n258_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n259_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n260_));
OR2X2 OR2X2_5341 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n257_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n260_), .Y(\col_out[26] ));
OR2X2 OR2X2_5342 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n262_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n263_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n264_));
OR2X2 OR2X2_5343 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n265_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n266_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n267_));
OR2X2 OR2X2_5344 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n264_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n267_), .Y(\col_out[27] ));
OR2X2 OR2X2_5345 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n269_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n270_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n271_));
OR2X2 OR2X2_5346 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n272_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n273_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n274_));
OR2X2 OR2X2_5347 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n271_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n274_), .Y(\col_out[28] ));
OR2X2 OR2X2_5348 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n276_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n277_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n278_));
OR2X2 OR2X2_5349 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n279_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n280_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n281_));
OR2X2 OR2X2_535 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3653_), .B(AES_CORE_DATAPATH__abc_16009_new_n3652_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3654_));
OR2X2 OR2X2_5350 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n278_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n281_), .Y(\col_out[29] ));
OR2X2 OR2X2_5351 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n283_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n284_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n285_));
OR2X2 OR2X2_5352 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n286_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n287_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n288_));
OR2X2 OR2X2_5353 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n285_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n288_), .Y(\col_out[30] ));
OR2X2 OR2X2_5354 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n290_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n291_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n292_));
OR2X2 OR2X2_5355 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n293_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n294_), .Y(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n295_));
OR2X2 OR2X2_5356 ( .A(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n292_), .B(AES_CORE_DATAPATH_SWAP_OUT__abc_15778_new_n295_), .Y(\col_out[31] ));
OR2X2 OR2X2_536 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3654_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3655_));
OR2X2 OR2X2_537 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3657_), .B(AES_CORE_DATAPATH__abc_16009_new_n3658_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_6_));
OR2X2 OR2X2_538 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3660_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3661_));
OR2X2 OR2X2_539 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3662_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3663_));
OR2X2 OR2X2_54 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n227_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n234_), .Y(AES_CORE_CONTROL_UNIT_col_sel_1_));
OR2X2 OR2X2_540 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3667_), .B(AES_CORE_DATAPATH__abc_16009_new_n3666_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3668_));
OR2X2 OR2X2_541 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3668_), .B(AES_CORE_DATAPATH__abc_16009_new_n3665_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3669_));
OR2X2 OR2X2_542 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3671_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3673_));
OR2X2 OR2X2_543 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3674_), .B(AES_CORE_DATAPATH__abc_16009_new_n3675_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3676_));
OR2X2 OR2X2_544 ( .A(\key_out[7] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3678_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3679_));
OR2X2 OR2X2_545 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3681_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3682_));
OR2X2 OR2X2_546 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3682_), .B(AES_CORE_DATAPATH__abc_16009_new_n3680_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3683_));
OR2X2 OR2X2_547 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3685_), .B(AES_CORE_DATAPATH__abc_16009_new_n3684_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3686_));
OR2X2 OR2X2_548 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3686_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3687_));
OR2X2 OR2X2_549 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3689_), .B(AES_CORE_DATAPATH__abc_16009_new_n3690_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_7_));
OR2X2 OR2X2_55 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT_key_out_sel_0_));
OR2X2 OR2X2_550 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3692_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3693_));
OR2X2 OR2X2_551 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3694_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3695_));
OR2X2 OR2X2_552 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3699_), .B(AES_CORE_DATAPATH__abc_16009_new_n3698_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3700_));
OR2X2 OR2X2_553 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3700_), .B(AES_CORE_DATAPATH__abc_16009_new_n3697_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3701_));
OR2X2 OR2X2_554 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3703_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3705_));
OR2X2 OR2X2_555 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3706_), .B(AES_CORE_DATAPATH__abc_16009_new_n3707_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3708_));
OR2X2 OR2X2_556 ( .A(\key_out[8] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3710_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3711_));
OR2X2 OR2X2_557 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3713_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3714_));
OR2X2 OR2X2_558 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3714_), .B(AES_CORE_DATAPATH__abc_16009_new_n3712_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3715_));
OR2X2 OR2X2_559 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3717_), .B(AES_CORE_DATAPATH__abc_16009_new_n3716_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3718_));
OR2X2 OR2X2_56 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n205_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT_key_out_sel_1_));
OR2X2 OR2X2_560 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3718_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3719_));
OR2X2 OR2X2_561 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3721_), .B(AES_CORE_DATAPATH__abc_16009_new_n3722_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_8_));
OR2X2 OR2X2_562 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3724_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3725_));
OR2X2 OR2X2_563 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3726_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3727_));
OR2X2 OR2X2_564 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3731_), .B(AES_CORE_DATAPATH__abc_16009_new_n3730_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3732_));
OR2X2 OR2X2_565 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3732_), .B(AES_CORE_DATAPATH__abc_16009_new_n3729_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3733_));
OR2X2 OR2X2_566 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3735_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3737_));
OR2X2 OR2X2_567 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3738_), .B(AES_CORE_DATAPATH__abc_16009_new_n3739_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3740_));
OR2X2 OR2X2_568 ( .A(\key_out[9] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3742_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3743_));
OR2X2 OR2X2_569 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3745_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3746_));
OR2X2 OR2X2_57 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n150_), .B(AES_CORE_CONTROL_UNIT_key_gen), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n239_));
OR2X2 OR2X2_570 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3746_), .B(AES_CORE_DATAPATH__abc_16009_new_n3744_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3747_));
OR2X2 OR2X2_571 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3749_), .B(AES_CORE_DATAPATH__abc_16009_new_n3748_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3750_));
OR2X2 OR2X2_572 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3750_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3751_));
OR2X2 OR2X2_573 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3753_), .B(AES_CORE_DATAPATH__abc_16009_new_n3754_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_9_));
OR2X2 OR2X2_574 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3756_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3757_));
OR2X2 OR2X2_575 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3758_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3759_));
OR2X2 OR2X2_576 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3763_), .B(AES_CORE_DATAPATH__abc_16009_new_n3762_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3764_));
OR2X2 OR2X2_577 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3764_), .B(AES_CORE_DATAPATH__abc_16009_new_n3761_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3765_));
OR2X2 OR2X2_578 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3767_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3769_));
OR2X2 OR2X2_579 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3770_), .B(AES_CORE_DATAPATH__abc_16009_new_n3771_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3772_));
OR2X2 OR2X2_58 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n239_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n193_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n240_));
OR2X2 OR2X2_580 ( .A(\key_out[10] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3774_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3775_));
OR2X2 OR2X2_581 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3777_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3778_));
OR2X2 OR2X2_582 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3778_), .B(AES_CORE_DATAPATH__abc_16009_new_n3776_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3779_));
OR2X2 OR2X2_583 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3781_), .B(AES_CORE_DATAPATH__abc_16009_new_n3780_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3782_));
OR2X2 OR2X2_584 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3782_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3783_));
OR2X2 OR2X2_585 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3785_), .B(AES_CORE_DATAPATH__abc_16009_new_n3786_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_10_));
OR2X2 OR2X2_586 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3788_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3789_));
OR2X2 OR2X2_587 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3790_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3791_));
OR2X2 OR2X2_588 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3795_), .B(AES_CORE_DATAPATH__abc_16009_new_n3794_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3796_));
OR2X2 OR2X2_589 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3796_), .B(AES_CORE_DATAPATH__abc_16009_new_n3793_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3797_));
OR2X2 OR2X2_59 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n240_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n238_), .Y(AES_CORE_CONTROL_UNIT_key_sel));
OR2X2 OR2X2_590 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3799_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3801_));
OR2X2 OR2X2_591 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3802_), .B(AES_CORE_DATAPATH__abc_16009_new_n3803_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3804_));
OR2X2 OR2X2_592 ( .A(\key_out[11] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3806_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3807_));
OR2X2 OR2X2_593 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3809_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3810_));
OR2X2 OR2X2_594 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3810_), .B(AES_CORE_DATAPATH__abc_16009_new_n3808_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3811_));
OR2X2 OR2X2_595 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3813_), .B(AES_CORE_DATAPATH__abc_16009_new_n3812_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3814_));
OR2X2 OR2X2_596 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3814_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3815_));
OR2X2 OR2X2_597 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3817_), .B(AES_CORE_DATAPATH__abc_16009_new_n3818_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_11_));
OR2X2 OR2X2_598 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3820_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3821_));
OR2X2 OR2X2_599 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3822_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3823_));
OR2X2 OR2X2_6 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n112_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n115_), .Y(AES_CORE_CONTROL_UNIT__abc_10772_auto_fsm_map_cc_170_map_fsm_1782_8_));
OR2X2 OR2X2_60 ( .A(AES_CORE_CONTROL_UNIT_key_gen), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT_key_en_0_));
OR2X2 OR2X2_600 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3827_), .B(AES_CORE_DATAPATH__abc_16009_new_n3826_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3828_));
OR2X2 OR2X2_601 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3828_), .B(AES_CORE_DATAPATH__abc_16009_new_n3825_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3829_));
OR2X2 OR2X2_602 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3831_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3833_));
OR2X2 OR2X2_603 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3834_), .B(AES_CORE_DATAPATH__abc_16009_new_n3835_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3836_));
OR2X2 OR2X2_604 ( .A(\key_out[12] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3838_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3839_));
OR2X2 OR2X2_605 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3841_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3842_));
OR2X2 OR2X2_606 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3842_), .B(AES_CORE_DATAPATH__abc_16009_new_n3840_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3843_));
OR2X2 OR2X2_607 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3845_), .B(AES_CORE_DATAPATH__abc_16009_new_n3844_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3846_));
OR2X2 OR2X2_608 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3846_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3847_));
OR2X2 OR2X2_609 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3849_), .B(AES_CORE_DATAPATH__abc_16009_new_n3850_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_12_));
OR2X2 OR2X2_61 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n244_), .B(AES_CORE_CONTROL_UNIT_state_3_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n245_));
OR2X2 OR2X2_610 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3852_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3853_));
OR2X2 OR2X2_611 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3854_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3855_));
OR2X2 OR2X2_612 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3859_), .B(AES_CORE_DATAPATH__abc_16009_new_n3858_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3860_));
OR2X2 OR2X2_613 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3860_), .B(AES_CORE_DATAPATH__abc_16009_new_n3857_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3861_));
OR2X2 OR2X2_614 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3863_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3865_));
OR2X2 OR2X2_615 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3866_), .B(AES_CORE_DATAPATH__abc_16009_new_n3867_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3868_));
OR2X2 OR2X2_616 ( .A(\key_out[13] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3870_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3871_));
OR2X2 OR2X2_617 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3873_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3874_));
OR2X2 OR2X2_618 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3874_), .B(AES_CORE_DATAPATH__abc_16009_new_n3872_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3875_));
OR2X2 OR2X2_619 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3877_), .B(AES_CORE_DATAPATH__abc_16009_new_n3876_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3878_));
OR2X2 OR2X2_62 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n245_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n243_), .Y(AES_CORE_CONTROL_UNIT_key_en_1_));
OR2X2 OR2X2_620 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3878_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3879_));
OR2X2 OR2X2_621 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3881_), .B(AES_CORE_DATAPATH__abc_16009_new_n3882_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_13_));
OR2X2 OR2X2_622 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3884_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3885_));
OR2X2 OR2X2_623 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3886_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3887_));
OR2X2 OR2X2_624 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3891_), .B(AES_CORE_DATAPATH__abc_16009_new_n3890_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3892_));
OR2X2 OR2X2_625 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3892_), .B(AES_CORE_DATAPATH__abc_16009_new_n3889_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3893_));
OR2X2 OR2X2_626 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3895_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3897_));
OR2X2 OR2X2_627 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3898_), .B(AES_CORE_DATAPATH__abc_16009_new_n3899_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3900_));
OR2X2 OR2X2_628 ( .A(\key_out[14] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3902_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3903_));
OR2X2 OR2X2_629 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3905_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3906_));
OR2X2 OR2X2_63 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_1_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n247_));
OR2X2 OR2X2_630 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3906_), .B(AES_CORE_DATAPATH__abc_16009_new_n3904_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3907_));
OR2X2 OR2X2_631 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3909_), .B(AES_CORE_DATAPATH__abc_16009_new_n3908_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3910_));
OR2X2 OR2X2_632 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3910_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3911_));
OR2X2 OR2X2_633 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3913_), .B(AES_CORE_DATAPATH__abc_16009_new_n3914_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_14_));
OR2X2 OR2X2_634 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3916_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3917_));
OR2X2 OR2X2_635 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3918_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3919_));
OR2X2 OR2X2_636 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3923_), .B(AES_CORE_DATAPATH__abc_16009_new_n3922_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3924_));
OR2X2 OR2X2_637 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3924_), .B(AES_CORE_DATAPATH__abc_16009_new_n3921_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3925_));
OR2X2 OR2X2_638 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3927_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3929_));
OR2X2 OR2X2_639 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3930_), .B(AES_CORE_DATAPATH__abc_16009_new_n3931_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3932_));
OR2X2 OR2X2_64 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n153_), .B(AES_CORE_CONTROL_UNIT_state_11_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n249_));
OR2X2 OR2X2_640 ( .A(\key_out[15] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3934_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3935_));
OR2X2 OR2X2_641 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3937_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3938_));
OR2X2 OR2X2_642 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3938_), .B(AES_CORE_DATAPATH__abc_16009_new_n3936_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3939_));
OR2X2 OR2X2_643 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3941_), .B(AES_CORE_DATAPATH__abc_16009_new_n3940_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3942_));
OR2X2 OR2X2_644 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3942_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3943_));
OR2X2 OR2X2_645 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3945_), .B(AES_CORE_DATAPATH__abc_16009_new_n3946_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_15_));
OR2X2 OR2X2_646 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3948_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3949_));
OR2X2 OR2X2_647 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3950_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3951_));
OR2X2 OR2X2_648 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3955_), .B(AES_CORE_DATAPATH__abc_16009_new_n3954_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3956_));
OR2X2 OR2X2_649 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3956_), .B(AES_CORE_DATAPATH__abc_16009_new_n3953_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3957_));
OR2X2 OR2X2_65 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n248_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n249_), .Y(AES_CORE_CONTROL_UNIT_key_en_2_));
OR2X2 OR2X2_650 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3959_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3961_));
OR2X2 OR2X2_651 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3962_), .B(AES_CORE_DATAPATH__abc_16009_new_n3963_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3964_));
OR2X2 OR2X2_652 ( .A(\key_out[16] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3966_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3967_));
OR2X2 OR2X2_653 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3969_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3970_));
OR2X2 OR2X2_654 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3970_), .B(AES_CORE_DATAPATH__abc_16009_new_n3968_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3971_));
OR2X2 OR2X2_655 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3973_), .B(AES_CORE_DATAPATH__abc_16009_new_n3972_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3974_));
OR2X2 OR2X2_656 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3974_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3975_));
OR2X2 OR2X2_657 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3977_), .B(AES_CORE_DATAPATH__abc_16009_new_n3978_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_16_));
OR2X2 OR2X2_658 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n3980_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3981_));
OR2X2 OR2X2_659 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n3982_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3983_));
OR2X2 OR2X2_66 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n252_), .B(AES_CORE_CONTROL_UNIT_state_7_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n253_));
OR2X2 OR2X2_660 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3987_), .B(AES_CORE_DATAPATH__abc_16009_new_n3986_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3988_));
OR2X2 OR2X2_661 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3988_), .B(AES_CORE_DATAPATH__abc_16009_new_n3985_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3989_));
OR2X2 OR2X2_662 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3991_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3993_));
OR2X2 OR2X2_663 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3994_), .B(AES_CORE_DATAPATH__abc_16009_new_n3995_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3996_));
OR2X2 OR2X2_664 ( .A(\key_out[17] ), .B(AES_CORE_DATAPATH__abc_16009_new_n3998_), .Y(AES_CORE_DATAPATH__abc_16009_new_n3999_));
OR2X2 OR2X2_665 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4001_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4002_));
OR2X2 OR2X2_666 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4002_), .B(AES_CORE_DATAPATH__abc_16009_new_n4000_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4003_));
OR2X2 OR2X2_667 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4005_), .B(AES_CORE_DATAPATH__abc_16009_new_n4004_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4006_));
OR2X2 OR2X2_668 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4006_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4007_));
OR2X2 OR2X2_669 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4009_), .B(AES_CORE_DATAPATH__abc_16009_new_n4010_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_17_));
OR2X2 OR2X2_67 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n253_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n251_), .Y(AES_CORE_CONTROL_UNIT_key_en_3_));
OR2X2 OR2X2_670 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4012_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4013_));
OR2X2 OR2X2_671 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4014_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4015_));
OR2X2 OR2X2_672 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4019_), .B(AES_CORE_DATAPATH__abc_16009_new_n4018_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4020_));
OR2X2 OR2X2_673 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4020_), .B(AES_CORE_DATAPATH__abc_16009_new_n4017_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4021_));
OR2X2 OR2X2_674 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4023_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4025_));
OR2X2 OR2X2_675 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4026_), .B(AES_CORE_DATAPATH__abc_16009_new_n4027_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4028_));
OR2X2 OR2X2_676 ( .A(\key_out[18] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4030_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4031_));
OR2X2 OR2X2_677 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4033_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4034_));
OR2X2 OR2X2_678 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4034_), .B(AES_CORE_DATAPATH__abc_16009_new_n4032_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4035_));
OR2X2 OR2X2_679 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4037_), .B(AES_CORE_DATAPATH__abc_16009_new_n4036_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4038_));
OR2X2 OR2X2_68 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n202_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_0_));
OR2X2 OR2X2_680 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4038_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4039_));
OR2X2 OR2X2_681 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4041_), .B(AES_CORE_DATAPATH__abc_16009_new_n4042_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_18_));
OR2X2 OR2X2_682 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4044_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4045_));
OR2X2 OR2X2_683 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4046_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4047_));
OR2X2 OR2X2_684 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4051_), .B(AES_CORE_DATAPATH__abc_16009_new_n4050_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4052_));
OR2X2 OR2X2_685 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4052_), .B(AES_CORE_DATAPATH__abc_16009_new_n4049_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4053_));
OR2X2 OR2X2_686 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4055_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4057_));
OR2X2 OR2X2_687 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4058_), .B(AES_CORE_DATAPATH__abc_16009_new_n4059_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4060_));
OR2X2 OR2X2_688 ( .A(\key_out[19] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4062_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4063_));
OR2X2 OR2X2_689 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4065_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4066_));
OR2X2 OR2X2_69 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n205_), .B(AES_CORE_CONTROL_UNIT__abc_15585_new_n208_), .Y(AES_CORE_CONTROL_UNIT_sbox_sel_1_));
OR2X2 OR2X2_690 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4066_), .B(AES_CORE_DATAPATH__abc_16009_new_n4064_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4067_));
OR2X2 OR2X2_691 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4069_), .B(AES_CORE_DATAPATH__abc_16009_new_n4068_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4070_));
OR2X2 OR2X2_692 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4070_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4071_));
OR2X2 OR2X2_693 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4073_), .B(AES_CORE_DATAPATH__abc_16009_new_n4074_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_19_));
OR2X2 OR2X2_694 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4076_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4077_));
OR2X2 OR2X2_695 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4078_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4079_));
OR2X2 OR2X2_696 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4083_), .B(AES_CORE_DATAPATH__abc_16009_new_n4082_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4084_));
OR2X2 OR2X2_697 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4084_), .B(AES_CORE_DATAPATH__abc_16009_new_n4081_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4085_));
OR2X2 OR2X2_698 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4087_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4089_));
OR2X2 OR2X2_699 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4090_), .B(AES_CORE_DATAPATH__abc_16009_new_n4091_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4092_));
OR2X2 OR2X2_7 ( .A(AES_CORE_CONTROL_UNIT__abc_15585_new_n84_), .B(AES_CORE_CONTROL_UNIT_state_14_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n117_));
OR2X2 OR2X2_70 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2459_), .B(AES_CORE_DATAPATH_col_en_host_2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2460_));
OR2X2 OR2X2_700 ( .A(\key_out[20] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4094_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4095_));
OR2X2 OR2X2_701 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4097_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4098_));
OR2X2 OR2X2_702 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4098_), .B(AES_CORE_DATAPATH__abc_16009_new_n4096_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4099_));
OR2X2 OR2X2_703 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4101_), .B(AES_CORE_DATAPATH__abc_16009_new_n4100_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4102_));
OR2X2 OR2X2_704 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4102_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4103_));
OR2X2 OR2X2_705 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4105_), .B(AES_CORE_DATAPATH__abc_16009_new_n4106_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_20_));
OR2X2 OR2X2_706 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4108_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4109_));
OR2X2 OR2X2_707 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4110_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4111_));
OR2X2 OR2X2_708 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4115_), .B(AES_CORE_DATAPATH__abc_16009_new_n4114_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4116_));
OR2X2 OR2X2_709 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4116_), .B(AES_CORE_DATAPATH__abc_16009_new_n4113_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4117_));
OR2X2 OR2X2_71 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2460_), .B(AES_CORE_DATAPATH__abc_16009_new_n2458_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2461_));
OR2X2 OR2X2_710 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4119_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4121_));
OR2X2 OR2X2_711 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4122_), .B(AES_CORE_DATAPATH__abc_16009_new_n4123_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4124_));
OR2X2 OR2X2_712 ( .A(\key_out[21] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4126_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4127_));
OR2X2 OR2X2_713 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4129_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4130_));
OR2X2 OR2X2_714 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4130_), .B(AES_CORE_DATAPATH__abc_16009_new_n4128_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4131_));
OR2X2 OR2X2_715 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4133_), .B(AES_CORE_DATAPATH__abc_16009_new_n4132_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4134_));
OR2X2 OR2X2_716 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4134_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4135_));
OR2X2 OR2X2_717 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4137_), .B(AES_CORE_DATAPATH__abc_16009_new_n4138_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_21_));
OR2X2 OR2X2_718 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4140_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4141_));
OR2X2 OR2X2_719 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4142_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4143_));
OR2X2 OR2X2_72 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2461_), .B(\iv_sel_rd[2] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2462_));
OR2X2 OR2X2_720 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4147_), .B(AES_CORE_DATAPATH__abc_16009_new_n4146_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4148_));
OR2X2 OR2X2_721 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4148_), .B(AES_CORE_DATAPATH__abc_16009_new_n4145_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4149_));
OR2X2 OR2X2_722 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4151_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4153_));
OR2X2 OR2X2_723 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4154_), .B(AES_CORE_DATAPATH__abc_16009_new_n4155_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4156_));
OR2X2 OR2X2_724 ( .A(\key_out[22] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4158_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4159_));
OR2X2 OR2X2_725 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4161_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4162_));
OR2X2 OR2X2_726 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4162_), .B(AES_CORE_DATAPATH__abc_16009_new_n4160_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4163_));
OR2X2 OR2X2_727 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4165_), .B(AES_CORE_DATAPATH__abc_16009_new_n4164_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4166_));
OR2X2 OR2X2_728 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4166_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4167_));
OR2X2 OR2X2_729 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4169_), .B(AES_CORE_DATAPATH__abc_16009_new_n4170_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_22_));
OR2X2 OR2X2_73 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2464_), .B(AES_CORE_DATAPATH_col_en_host_1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2465_));
OR2X2 OR2X2_730 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4172_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4173_));
OR2X2 OR2X2_731 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4174_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4175_));
OR2X2 OR2X2_732 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4179_), .B(AES_CORE_DATAPATH__abc_16009_new_n4178_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4180_));
OR2X2 OR2X2_733 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4180_), .B(AES_CORE_DATAPATH__abc_16009_new_n4177_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4181_));
OR2X2 OR2X2_734 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4183_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4185_));
OR2X2 OR2X2_735 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4186_), .B(AES_CORE_DATAPATH__abc_16009_new_n4187_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4188_));
OR2X2 OR2X2_736 ( .A(\key_out[23] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4190_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4191_));
OR2X2 OR2X2_737 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4193_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4194_));
OR2X2 OR2X2_738 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4194_), .B(AES_CORE_DATAPATH__abc_16009_new_n4192_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4195_));
OR2X2 OR2X2_739 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4197_), .B(AES_CORE_DATAPATH__abc_16009_new_n4196_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4198_));
OR2X2 OR2X2_74 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2465_), .B(AES_CORE_DATAPATH__abc_16009_new_n2463_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2466_));
OR2X2 OR2X2_740 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4198_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4199_));
OR2X2 OR2X2_741 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4201_), .B(AES_CORE_DATAPATH__abc_16009_new_n4202_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_23_));
OR2X2 OR2X2_742 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4204_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4205_));
OR2X2 OR2X2_743 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4206_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4207_));
OR2X2 OR2X2_744 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4211_), .B(AES_CORE_DATAPATH__abc_16009_new_n4210_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4212_));
OR2X2 OR2X2_745 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4212_), .B(AES_CORE_DATAPATH__abc_16009_new_n4209_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4213_));
OR2X2 OR2X2_746 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4215_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4217_));
OR2X2 OR2X2_747 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4218_), .B(AES_CORE_DATAPATH__abc_16009_new_n4219_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4220_));
OR2X2 OR2X2_748 ( .A(\key_out[24] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4222_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4223_));
OR2X2 OR2X2_749 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4225_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4226_));
OR2X2 OR2X2_75 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2466_), .B(\iv_sel_rd[1] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2467_));
OR2X2 OR2X2_750 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4226_), .B(AES_CORE_DATAPATH__abc_16009_new_n4224_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4227_));
OR2X2 OR2X2_751 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4229_), .B(AES_CORE_DATAPATH__abc_16009_new_n4228_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4230_));
OR2X2 OR2X2_752 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4230_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4231_));
OR2X2 OR2X2_753 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4233_), .B(AES_CORE_DATAPATH__abc_16009_new_n4234_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_24_));
OR2X2 OR2X2_754 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4236_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4237_));
OR2X2 OR2X2_755 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4238_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4239_));
OR2X2 OR2X2_756 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4243_), .B(AES_CORE_DATAPATH__abc_16009_new_n4242_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4244_));
OR2X2 OR2X2_757 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4244_), .B(AES_CORE_DATAPATH__abc_16009_new_n4241_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4245_));
OR2X2 OR2X2_758 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4247_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4249_));
OR2X2 OR2X2_759 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4250_), .B(AES_CORE_DATAPATH__abc_16009_new_n4251_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4252_));
OR2X2 OR2X2_76 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2469_), .B(AES_CORE_DATAPATH_col_en_host_0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2470_));
OR2X2 OR2X2_760 ( .A(\key_out[25] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4254_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4255_));
OR2X2 OR2X2_761 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4257_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4258_));
OR2X2 OR2X2_762 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4258_), .B(AES_CORE_DATAPATH__abc_16009_new_n4256_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4259_));
OR2X2 OR2X2_763 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4261_), .B(AES_CORE_DATAPATH__abc_16009_new_n4260_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4262_));
OR2X2 OR2X2_764 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4262_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4263_));
OR2X2 OR2X2_765 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4265_), .B(AES_CORE_DATAPATH__abc_16009_new_n4266_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_25_));
OR2X2 OR2X2_766 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4268_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4269_));
OR2X2 OR2X2_767 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4270_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4271_));
OR2X2 OR2X2_768 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4275_), .B(AES_CORE_DATAPATH__abc_16009_new_n4274_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4276_));
OR2X2 OR2X2_769 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4276_), .B(AES_CORE_DATAPATH__abc_16009_new_n4273_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4277_));
OR2X2 OR2X2_77 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2470_), .B(AES_CORE_DATAPATH__abc_16009_new_n2468_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2471_));
OR2X2 OR2X2_770 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4279_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4281_));
OR2X2 OR2X2_771 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4282_), .B(AES_CORE_DATAPATH__abc_16009_new_n4283_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4284_));
OR2X2 OR2X2_772 ( .A(\key_out[26] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4286_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4287_));
OR2X2 OR2X2_773 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4289_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4290_));
OR2X2 OR2X2_774 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4290_), .B(AES_CORE_DATAPATH__abc_16009_new_n4288_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4291_));
OR2X2 OR2X2_775 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4293_), .B(AES_CORE_DATAPATH__abc_16009_new_n4292_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4294_));
OR2X2 OR2X2_776 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4294_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4295_));
OR2X2 OR2X2_777 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4297_), .B(AES_CORE_DATAPATH__abc_16009_new_n4298_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_26_));
OR2X2 OR2X2_778 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4300_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4301_));
OR2X2 OR2X2_779 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4302_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4303_));
OR2X2 OR2X2_78 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2471_), .B(\iv_sel_rd[0] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2472_));
OR2X2 OR2X2_780 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4307_), .B(AES_CORE_DATAPATH__abc_16009_new_n4306_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4308_));
OR2X2 OR2X2_781 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4308_), .B(AES_CORE_DATAPATH__abc_16009_new_n4305_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4309_));
OR2X2 OR2X2_782 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4311_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4313_));
OR2X2 OR2X2_783 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4314_), .B(AES_CORE_DATAPATH__abc_16009_new_n4315_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4316_));
OR2X2 OR2X2_784 ( .A(\key_out[27] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4318_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4319_));
OR2X2 OR2X2_785 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4321_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4322_));
OR2X2 OR2X2_786 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4322_), .B(AES_CORE_DATAPATH__abc_16009_new_n4320_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4323_));
OR2X2 OR2X2_787 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4325_), .B(AES_CORE_DATAPATH__abc_16009_new_n4324_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4326_));
OR2X2 OR2X2_788 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4326_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4327_));
OR2X2 OR2X2_789 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4329_), .B(AES_CORE_DATAPATH__abc_16009_new_n4330_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_27_));
OR2X2 OR2X2_79 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2473_), .B(AES_CORE_DATAPATH__abc_16009_new_n2467_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2474_));
OR2X2 OR2X2_790 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4332_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4333_));
OR2X2 OR2X2_791 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4334_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4335_));
OR2X2 OR2X2_792 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4339_), .B(AES_CORE_DATAPATH__abc_16009_new_n4338_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4340_));
OR2X2 OR2X2_793 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4340_), .B(AES_CORE_DATAPATH__abc_16009_new_n4337_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4341_));
OR2X2 OR2X2_794 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4343_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4345_));
OR2X2 OR2X2_795 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4346_), .B(AES_CORE_DATAPATH__abc_16009_new_n4347_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4348_));
OR2X2 OR2X2_796 ( .A(\key_out[28] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4350_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4351_));
OR2X2 OR2X2_797 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4353_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4354_));
OR2X2 OR2X2_798 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4354_), .B(AES_CORE_DATAPATH__abc_16009_new_n4352_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4355_));
OR2X2 OR2X2_799 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4357_), .B(AES_CORE_DATAPATH__abc_16009_new_n4356_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4358_));
OR2X2 OR2X2_8 ( .A(AES_CORE_CONTROL_UNIT_encrypt_decrypt), .B(AES_CORE_CONTROL_UNIT_state_9_), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n118_));
OR2X2 OR2X2_80 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2475_), .B(AES_CORE_DATAPATH_iv_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2476_));
OR2X2 OR2X2_800 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4358_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4359_));
OR2X2 OR2X2_801 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4361_), .B(AES_CORE_DATAPATH__abc_16009_new_n4362_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_28_));
OR2X2 OR2X2_802 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4364_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4365_));
OR2X2 OR2X2_803 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4366_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4367_));
OR2X2 OR2X2_804 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4371_), .B(AES_CORE_DATAPATH__abc_16009_new_n4370_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4372_));
OR2X2 OR2X2_805 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4372_), .B(AES_CORE_DATAPATH__abc_16009_new_n4369_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4373_));
OR2X2 OR2X2_806 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4375_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4377_));
OR2X2 OR2X2_807 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4378_), .B(AES_CORE_DATAPATH__abc_16009_new_n4379_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4380_));
OR2X2 OR2X2_808 ( .A(\key_out[29] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4382_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4383_));
OR2X2 OR2X2_809 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4385_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4386_));
OR2X2 OR2X2_81 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2477_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2478_));
OR2X2 OR2X2_810 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4386_), .B(AES_CORE_DATAPATH__abc_16009_new_n4384_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4387_));
OR2X2 OR2X2_811 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4389_), .B(AES_CORE_DATAPATH__abc_16009_new_n4388_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4390_));
OR2X2 OR2X2_812 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4390_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4391_));
OR2X2 OR2X2_813 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4393_), .B(AES_CORE_DATAPATH__abc_16009_new_n4394_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_29_));
OR2X2 OR2X2_814 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4396_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4397_));
OR2X2 OR2X2_815 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4398_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4399_));
OR2X2 OR2X2_816 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4403_), .B(AES_CORE_DATAPATH__abc_16009_new_n4402_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4404_));
OR2X2 OR2X2_817 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4404_), .B(AES_CORE_DATAPATH__abc_16009_new_n4401_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4405_));
OR2X2 OR2X2_818 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4407_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4409_));
OR2X2 OR2X2_819 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4410_), .B(AES_CORE_DATAPATH__abc_16009_new_n4411_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4412_));
OR2X2 OR2X2_82 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2480_), .B(AES_CORE_DATAPATH_col_en_host_3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2481_));
OR2X2 OR2X2_820 ( .A(\key_out[30] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4414_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4415_));
OR2X2 OR2X2_821 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4417_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4418_));
OR2X2 OR2X2_822 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4418_), .B(AES_CORE_DATAPATH__abc_16009_new_n4416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4419_));
OR2X2 OR2X2_823 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4421_), .B(AES_CORE_DATAPATH__abc_16009_new_n4420_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4422_));
OR2X2 OR2X2_824 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4422_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4423_));
OR2X2 OR2X2_825 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4425_), .B(AES_CORE_DATAPATH__abc_16009_new_n4426_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_30_));
OR2X2 OR2X2_826 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4428_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4429_));
OR2X2 OR2X2_827 ( .A(AES_CORE_DATAPATH__abc_16009_new_n3427_), .B(AES_CORE_DATAPATH__abc_16009_new_n4430_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4431_));
OR2X2 OR2X2_828 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4435_), .B(AES_CORE_DATAPATH__abc_16009_new_n4434_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4436_));
OR2X2 OR2X2_829 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4436_), .B(AES_CORE_DATAPATH__abc_16009_new_n4433_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4437_));
OR2X2 OR2X2_83 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2481_), .B(AES_CORE_DATAPATH__abc_16009_new_n2479_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2482_));
OR2X2 OR2X2_830 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4439_), .B(AES_CORE_DATAPATH__abc_16009_new_n3416_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4441_));
OR2X2 OR2X2_831 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4442_), .B(AES_CORE_DATAPATH__abc_16009_new_n4443_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4444_));
OR2X2 OR2X2_832 ( .A(\key_out[31] ), .B(AES_CORE_DATAPATH__abc_16009_new_n4446_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4447_));
OR2X2 OR2X2_833 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4449_), .B(AES_CORE_DATAPATH__abc_16009_new_n3456_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4450_));
OR2X2 OR2X2_834 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4450_), .B(AES_CORE_DATAPATH__abc_16009_new_n4448_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4451_));
OR2X2 OR2X2_835 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4453_), .B(AES_CORE_DATAPATH__abc_16009_new_n4452_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4454_));
OR2X2 OR2X2_836 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4454_), .B(AES_CORE_DATAPATH__abc_16009_new_n3455_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4455_));
OR2X2 OR2X2_837 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4457_), .B(AES_CORE_DATAPATH__abc_16009_new_n4458_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_31_));
OR2X2 OR2X2_838 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4461_), .B(AES_CORE_DATAPATH__abc_16009_new_n4460_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_96_));
OR2X2 OR2X2_839 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4464_), .B(AES_CORE_DATAPATH__abc_16009_new_n4463_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_97_));
OR2X2 OR2X2_84 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2482_), .B(\iv_sel_rd[3] ), .Y(AES_CORE_DATAPATH__abc_16009_new_n2483_));
OR2X2 OR2X2_840 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4467_), .B(AES_CORE_DATAPATH__abc_16009_new_n4466_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_98_));
OR2X2 OR2X2_841 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4470_), .B(AES_CORE_DATAPATH__abc_16009_new_n4469_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_99_));
OR2X2 OR2X2_842 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4473_), .B(AES_CORE_DATAPATH__abc_16009_new_n4472_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_100_));
OR2X2 OR2X2_843 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4476_), .B(AES_CORE_DATAPATH__abc_16009_new_n4475_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_101_));
OR2X2 OR2X2_844 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4479_), .B(AES_CORE_DATAPATH__abc_16009_new_n4478_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_102_));
OR2X2 OR2X2_845 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4482_), .B(AES_CORE_DATAPATH__abc_16009_new_n4481_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_103_));
OR2X2 OR2X2_846 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4485_), .B(AES_CORE_DATAPATH__abc_16009_new_n4484_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_104_));
OR2X2 OR2X2_847 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4488_), .B(AES_CORE_DATAPATH__abc_16009_new_n4487_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_105_));
OR2X2 OR2X2_848 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4491_), .B(AES_CORE_DATAPATH__abc_16009_new_n4490_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_106_));
OR2X2 OR2X2_849 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4494_), .B(AES_CORE_DATAPATH__abc_16009_new_n4493_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_107_));
OR2X2 OR2X2_85 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2486_));
OR2X2 OR2X2_850 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4497_), .B(AES_CORE_DATAPATH__abc_16009_new_n4496_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_108_));
OR2X2 OR2X2_851 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4500_), .B(AES_CORE_DATAPATH__abc_16009_new_n4499_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_109_));
OR2X2 OR2X2_852 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4503_), .B(AES_CORE_DATAPATH__abc_16009_new_n4502_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_110_));
OR2X2 OR2X2_853 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4506_), .B(AES_CORE_DATAPATH__abc_16009_new_n4505_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_111_));
OR2X2 OR2X2_854 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4509_), .B(AES_CORE_DATAPATH__abc_16009_new_n4508_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_112_));
OR2X2 OR2X2_855 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4512_), .B(AES_CORE_DATAPATH__abc_16009_new_n4511_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_113_));
OR2X2 OR2X2_856 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4515_), .B(AES_CORE_DATAPATH__abc_16009_new_n4514_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_114_));
OR2X2 OR2X2_857 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4518_), .B(AES_CORE_DATAPATH__abc_16009_new_n4517_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_115_));
OR2X2 OR2X2_858 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4521_), .B(AES_CORE_DATAPATH__abc_16009_new_n4520_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_116_));
OR2X2 OR2X2_859 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4524_), .B(AES_CORE_DATAPATH__abc_16009_new_n4523_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_117_));
OR2X2 OR2X2_86 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2488_), .B(AES_CORE_DATAPATH__abc_16009_new_n2489_), .Y(\iv_out[0] ));
OR2X2 OR2X2_860 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4527_), .B(AES_CORE_DATAPATH__abc_16009_new_n4526_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_118_));
OR2X2 OR2X2_861 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4530_), .B(AES_CORE_DATAPATH__abc_16009_new_n4529_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_119_));
OR2X2 OR2X2_862 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4533_), .B(AES_CORE_DATAPATH__abc_16009_new_n4532_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_120_));
OR2X2 OR2X2_863 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4536_), .B(AES_CORE_DATAPATH__abc_16009_new_n4535_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_121_));
OR2X2 OR2X2_864 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4539_), .B(AES_CORE_DATAPATH__abc_16009_new_n4538_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_122_));
OR2X2 OR2X2_865 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4542_), .B(AES_CORE_DATAPATH__abc_16009_new_n4541_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_123_));
OR2X2 OR2X2_866 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4545_), .B(AES_CORE_DATAPATH__abc_16009_new_n4544_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_124_));
OR2X2 OR2X2_867 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4548_), .B(AES_CORE_DATAPATH__abc_16009_new_n4547_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_125_));
OR2X2 OR2X2_868 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4551_), .B(AES_CORE_DATAPATH__abc_16009_new_n4550_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_126_));
OR2X2 OR2X2_869 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4554_), .B(AES_CORE_DATAPATH__abc_16009_new_n4553_), .Y(AES_CORE_DATAPATH_SHIFT_ROW_data_in_127_));
OR2X2 OR2X2_87 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2493_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2494_));
OR2X2 OR2X2_870 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2805_), .B(AES_CORE_CONTROL_UNIT_bypass_rk), .Y(AES_CORE_DATAPATH_rk_out_sel));
OR2X2 OR2X2_871 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4557_), .B(AES_CORE_DATAPATH__abc_16009_new_n4558_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4559_));
OR2X2 OR2X2_872 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4565_), .B(AES_CORE_DATAPATH__abc_16009_new_n4566_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4567_));
OR2X2 OR2X2_873 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4569_), .B(AES_CORE_DATAPATH__abc_16009_new_n4568_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4570_));
OR2X2 OR2X2_874 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4570_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4571_));
OR2X2 OR2X2_875 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_64_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4573_));
OR2X2 OR2X2_876 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4574_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4575_));
OR2X2 OR2X2_877 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__0_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4577_));
OR2X2 OR2X2_878 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_65_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4579_));
OR2X2 OR2X2_879 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4580_), .B(AES_CORE_DATAPATH__abc_16009_new_n4581_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4582_));
OR2X2 OR2X2_88 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2494_), .B(AES_CORE_DATAPATH__abc_16009_new_n2492_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2495_));
OR2X2 OR2X2_880 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4582_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4583_));
OR2X2 OR2X2_881 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4585_), .B(AES_CORE_DATAPATH__abc_16009_new_n4586_), .Y(AES_CORE_DATAPATH__0key_1__31_0__1_));
OR2X2 OR2X2_882 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_66_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4588_));
OR2X2 OR2X2_883 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4589_), .B(AES_CORE_DATAPATH__abc_16009_new_n4590_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4591_));
OR2X2 OR2X2_884 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4591_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4592_));
OR2X2 OR2X2_885 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4594_), .B(AES_CORE_DATAPATH__abc_16009_new_n4595_), .Y(AES_CORE_DATAPATH__0key_1__31_0__2_));
OR2X2 OR2X2_886 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_67_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4597_));
OR2X2 OR2X2_887 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4598_), .B(AES_CORE_DATAPATH__abc_16009_new_n4599_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4600_));
OR2X2 OR2X2_888 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4600_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4601_));
OR2X2 OR2X2_889 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4603_), .B(AES_CORE_DATAPATH__abc_16009_new_n4604_), .Y(AES_CORE_DATAPATH__0key_1__31_0__3_));
OR2X2 OR2X2_89 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__1_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2496_));
OR2X2 OR2X2_890 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_68_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4606_));
OR2X2 OR2X2_891 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4607_), .B(AES_CORE_DATAPATH__abc_16009_new_n4608_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4609_));
OR2X2 OR2X2_892 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4609_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4610_));
OR2X2 OR2X2_893 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4612_), .B(AES_CORE_DATAPATH__abc_16009_new_n4613_), .Y(AES_CORE_DATAPATH__0key_1__31_0__4_));
OR2X2 OR2X2_894 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_69_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4615_));
OR2X2 OR2X2_895 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4616_), .B(AES_CORE_DATAPATH__abc_16009_new_n4617_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4618_));
OR2X2 OR2X2_896 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4618_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4619_));
OR2X2 OR2X2_897 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4621_), .B(AES_CORE_DATAPATH__abc_16009_new_n4622_), .Y(AES_CORE_DATAPATH__0key_1__31_0__5_));
OR2X2 OR2X2_898 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_70_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4624_));
OR2X2 OR2X2_899 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4625_), .B(AES_CORE_DATAPATH__abc_16009_new_n4626_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4627_));
OR2X2 OR2X2_9 ( .A(disable_core), .B(end_aes), .Y(AES_CORE_CONTROL_UNIT__abc_15585_new_n123_));
OR2X2 OR2X2_90 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2498_), .B(AES_CORE_DATAPATH__abc_16009_new_n2499_), .Y(\iv_out[1] ));
OR2X2 OR2X2_900 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4627_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4628_));
OR2X2 OR2X2_901 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4630_), .B(AES_CORE_DATAPATH__abc_16009_new_n4631_), .Y(AES_CORE_DATAPATH__0key_1__31_0__6_));
OR2X2 OR2X2_902 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_71_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4633_));
OR2X2 OR2X2_903 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4634_), .B(AES_CORE_DATAPATH__abc_16009_new_n4635_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4636_));
OR2X2 OR2X2_904 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4636_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4637_));
OR2X2 OR2X2_905 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4638_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4639_));
OR2X2 OR2X2_906 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__7_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4640_));
OR2X2 OR2X2_907 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_72_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4642_));
OR2X2 OR2X2_908 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4643_), .B(AES_CORE_DATAPATH__abc_16009_new_n4644_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4645_));
OR2X2 OR2X2_909 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4645_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4646_));
OR2X2 OR2X2_91 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2503_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2504_));
OR2X2 OR2X2_910 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4648_), .B(AES_CORE_DATAPATH__abc_16009_new_n4649_), .Y(AES_CORE_DATAPATH__0key_1__31_0__8_));
OR2X2 OR2X2_911 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_73_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4651_));
OR2X2 OR2X2_912 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4652_), .B(AES_CORE_DATAPATH__abc_16009_new_n4653_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4654_));
OR2X2 OR2X2_913 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4654_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4655_));
OR2X2 OR2X2_914 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4657_), .B(AES_CORE_DATAPATH__abc_16009_new_n4658_), .Y(AES_CORE_DATAPATH__0key_1__31_0__9_));
OR2X2 OR2X2_915 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_74_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4660_));
OR2X2 OR2X2_916 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4661_), .B(AES_CORE_DATAPATH__abc_16009_new_n4662_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4663_));
OR2X2 OR2X2_917 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4663_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4664_));
OR2X2 OR2X2_918 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4665_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4666_));
OR2X2 OR2X2_919 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__10_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4667_));
OR2X2 OR2X2_92 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2504_), .B(AES_CORE_DATAPATH__abc_16009_new_n2502_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2505_));
OR2X2 OR2X2_920 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_75_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4669_));
OR2X2 OR2X2_921 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4670_), .B(AES_CORE_DATAPATH__abc_16009_new_n4671_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4672_));
OR2X2 OR2X2_922 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4672_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4673_));
OR2X2 OR2X2_923 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4674_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4675_));
OR2X2 OR2X2_924 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__11_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4676_));
OR2X2 OR2X2_925 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_76_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4678_));
OR2X2 OR2X2_926 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4679_), .B(AES_CORE_DATAPATH__abc_16009_new_n4680_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4681_));
OR2X2 OR2X2_927 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4681_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4682_));
OR2X2 OR2X2_928 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4683_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4684_));
OR2X2 OR2X2_929 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__12_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4685_));
OR2X2 OR2X2_93 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__2_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2506_));
OR2X2 OR2X2_930 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_77_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4687_));
OR2X2 OR2X2_931 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4688_), .B(AES_CORE_DATAPATH__abc_16009_new_n4689_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4690_));
OR2X2 OR2X2_932 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4690_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4691_));
OR2X2 OR2X2_933 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4692_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4693_));
OR2X2 OR2X2_934 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__13_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4694_));
OR2X2 OR2X2_935 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_78_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4696_));
OR2X2 OR2X2_936 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4697_), .B(AES_CORE_DATAPATH__abc_16009_new_n4698_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4699_));
OR2X2 OR2X2_937 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4699_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4700_));
OR2X2 OR2X2_938 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4702_), .B(AES_CORE_DATAPATH__abc_16009_new_n4703_), .Y(AES_CORE_DATAPATH__0key_1__31_0__14_));
OR2X2 OR2X2_939 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_79_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4705_));
OR2X2 OR2X2_94 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2508_), .B(AES_CORE_DATAPATH__abc_16009_new_n2509_), .Y(\iv_out[2] ));
OR2X2 OR2X2_940 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4706_), .B(AES_CORE_DATAPATH__abc_16009_new_n4707_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4708_));
OR2X2 OR2X2_941 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4708_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4709_));
OR2X2 OR2X2_942 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4711_), .B(AES_CORE_DATAPATH__abc_16009_new_n4712_), .Y(AES_CORE_DATAPATH__0key_1__31_0__15_));
OR2X2 OR2X2_943 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_80_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4714_));
OR2X2 OR2X2_944 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4715_), .B(AES_CORE_DATAPATH__abc_16009_new_n4716_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4717_));
OR2X2 OR2X2_945 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4717_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4718_));
OR2X2 OR2X2_946 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4719_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4720_));
OR2X2 OR2X2_947 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__16_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4721_));
OR2X2 OR2X2_948 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_81_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4723_));
OR2X2 OR2X2_949 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4724_), .B(AES_CORE_DATAPATH__abc_16009_new_n4725_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4726_));
OR2X2 OR2X2_95 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2513_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2514_));
OR2X2 OR2X2_950 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4726_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4727_));
OR2X2 OR2X2_951 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4728_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4729_));
OR2X2 OR2X2_952 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__17_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4730_));
OR2X2 OR2X2_953 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_82_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4732_));
OR2X2 OR2X2_954 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4733_), .B(AES_CORE_DATAPATH__abc_16009_new_n4734_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4735_));
OR2X2 OR2X2_955 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4735_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4736_));
OR2X2 OR2X2_956 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4737_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4738_));
OR2X2 OR2X2_957 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__18_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4739_));
OR2X2 OR2X2_958 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_83_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4741_));
OR2X2 OR2X2_959 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4742_), .B(AES_CORE_DATAPATH__abc_16009_new_n4743_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4744_));
OR2X2 OR2X2_96 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2514_), .B(AES_CORE_DATAPATH__abc_16009_new_n2512_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2515_));
OR2X2 OR2X2_960 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4744_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4745_));
OR2X2 OR2X2_961 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4747_), .B(AES_CORE_DATAPATH__abc_16009_new_n4748_), .Y(AES_CORE_DATAPATH__0key_1__31_0__19_));
OR2X2 OR2X2_962 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_84_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4750_));
OR2X2 OR2X2_963 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4751_), .B(AES_CORE_DATAPATH__abc_16009_new_n4752_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4753_));
OR2X2 OR2X2_964 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4753_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4754_));
OR2X2 OR2X2_965 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4756_), .B(AES_CORE_DATAPATH__abc_16009_new_n4757_), .Y(AES_CORE_DATAPATH__0key_1__31_0__20_));
OR2X2 OR2X2_966 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_85_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4759_));
OR2X2 OR2X2_967 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4760_), .B(AES_CORE_DATAPATH__abc_16009_new_n4761_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4762_));
OR2X2 OR2X2_968 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4762_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4763_));
OR2X2 OR2X2_969 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4765_), .B(AES_CORE_DATAPATH__abc_16009_new_n4766_), .Y(AES_CORE_DATAPATH__0key_1__31_0__21_));
OR2X2 OR2X2_97 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2485_), .B(AES_CORE_DATAPATH_iv_2__3_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2516_));
OR2X2 OR2X2_970 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_86_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4768_));
OR2X2 OR2X2_971 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4769_), .B(AES_CORE_DATAPATH__abc_16009_new_n4770_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4771_));
OR2X2 OR2X2_972 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4771_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4772_));
OR2X2 OR2X2_973 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4773_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4774_));
OR2X2 OR2X2_974 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__22_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4775_));
OR2X2 OR2X2_975 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_87_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4777_));
OR2X2 OR2X2_976 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4778_), .B(AES_CORE_DATAPATH__abc_16009_new_n4779_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4780_));
OR2X2 OR2X2_977 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4780_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4781_));
OR2X2 OR2X2_978 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4783_), .B(AES_CORE_DATAPATH__abc_16009_new_n4784_), .Y(AES_CORE_DATAPATH__0key_1__31_0__23_));
OR2X2 OR2X2_979 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_88_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4786_));
OR2X2 OR2X2_98 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2518_), .B(AES_CORE_DATAPATH__abc_16009_new_n2519_), .Y(\iv_out[3] ));
OR2X2 OR2X2_980 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4787_), .B(AES_CORE_DATAPATH__abc_16009_new_n4788_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4789_));
OR2X2 OR2X2_981 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4789_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4790_));
OR2X2 OR2X2_982 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4791_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4792_));
OR2X2 OR2X2_983 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__24_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4793_));
OR2X2 OR2X2_984 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_89_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4795_));
OR2X2 OR2X2_985 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4796_), .B(AES_CORE_DATAPATH__abc_16009_new_n4797_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4798_));
OR2X2 OR2X2_986 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4798_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4799_));
OR2X2 OR2X2_987 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4801_), .B(AES_CORE_DATAPATH__abc_16009_new_n4802_), .Y(AES_CORE_DATAPATH__0key_1__31_0__25_));
OR2X2 OR2X2_988 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_90_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4804_));
OR2X2 OR2X2_989 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4805_), .B(AES_CORE_DATAPATH__abc_16009_new_n4806_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4807_));
OR2X2 OR2X2_99 ( .A(AES_CORE_DATAPATH__abc_16009_new_n2523_), .B(AES_CORE_DATAPATH__abc_16009_new_n2462_), .Y(AES_CORE_DATAPATH__abc_16009_new_n2524_));
OR2X2 OR2X2_990 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4807_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4808_));
OR2X2 OR2X2_991 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4809_), .B(AES_CORE_DATAPATH__abc_16009_new_n4564_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4810_));
OR2X2 OR2X2_992 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4576_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_1__26_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4811_));
OR2X2 OR2X2_993 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_91_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4813_));
OR2X2 OR2X2_994 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4814_), .B(AES_CORE_DATAPATH__abc_16009_new_n4815_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4816_));
OR2X2 OR2X2_995 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4816_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4817_));
OR2X2 OR2X2_996 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4819_), .B(AES_CORE_DATAPATH__abc_16009_new_n4820_), .Y(AES_CORE_DATAPATH__0key_1__31_0__27_));
OR2X2 OR2X2_997 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4572_), .B(AES_CORE_DATAPATH_KEY_EXPANDER_key_out_92_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4822_));
OR2X2 OR2X2_998 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4823_), .B(AES_CORE_DATAPATH__abc_16009_new_n4824_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4825_));
OR2X2 OR2X2_999 ( .A(AES_CORE_DATAPATH__abc_16009_new_n4567_), .B(AES_CORE_DATAPATH__abc_16009_new_n4825_), .Y(AES_CORE_DATAPATH__abc_16009_new_n4826_));


endmodule